//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_200_assert(
  input        _EVAL,
  input        _EVAL_1,
  input        _EVAL_2,
  input  [3:0] _EVAL_5
);
  wire  _EVAL_4;
  wire  _EVAL_6;
  wire  _EVAL_8;
  wire  _EVAL_10;
  wire  _EVAL_13;
  wire  _EVAL_14;
  wire  _EVAL_15;
  wire  _EVAL_18;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_43;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_50;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_64;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_70;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_77;
  wire  _EVAL_80;
  wire  _EVAL_82;
  wire  _EVAL_84;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  assign _EVAL_4 = _EVAL_14 & _EVAL_80;
  assign _EVAL_73 = _EVAL_10 & _EVAL_2;
  assign _EVAL_70 = _EVAL_59 & _EVAL_24;
  assign _EVAL_10 = _EVAL_5 == 4'h6;
  assign _EVAL_96 = _EVAL_21 & _EVAL_80;
  assign _EVAL_59 = _EVAL_5 == 4'h8;
  assign _EVAL_74 = _EVAL_5 == 4'h9;
  assign _EVAL_111 = _EVAL_5 == 4'h4;
  assign _EVAL_72 = _EVAL_74 & _EVAL_2;
  assign _EVAL_62 = _EVAL_37 & _EVAL_2;
  assign _EVAL_113 = _EVAL_54 & _EVAL_80;
  assign _EVAL_28 = _EVAL_6 & _EVAL_24;
  assign _EVAL_43 = _EVAL_50 & _EVAL_80;
  assign _EVAL_106 = _EVAL_6 & _EVAL_80;
  assign _EVAL_18 = _EVAL_5 == 4'h7;
  assign _EVAL_67 = _EVAL_59 & _EVAL_80;
  assign _EVAL_13 = _EVAL_5 == 4'h2;
  assign _EVAL_45 = _EVAL_55 & _EVAL_80;
  assign _EVAL_84 = _EVAL_5 == 4'h5;
  assign _EVAL_31 = _EVAL_5 == 4'hf;
  assign _EVAL_15 = _EVAL_10 & _EVAL_80;
  assign _EVAL_46 = _EVAL_31 & _EVAL_80;
  assign _EVAL_61 = _EVAL_14 & _EVAL_2;
  assign _EVAL_54 = _EVAL_5 == 4'ha;
  assign _EVAL_109 = _EVAL_5 == 4'hb;
  assign _EVAL_58 = _EVAL_54 & _EVAL_24;
  assign _EVAL_98 = _EVAL_31 & _EVAL_24;
  assign _EVAL_23 = _EVAL_109 & _EVAL_80;
  assign _EVAL_91 = _EVAL_13 & _EVAL_24;
  assign _EVAL_21 = _EVAL_5 == 4'h3;
  assign _EVAL_89 = _EVAL_31 & _EVAL_2;
  assign _EVAL_88 = _EVAL_109 & _EVAL_24;
  assign _EVAL_50 = _EVAL_5 == 4'hc;
  assign _EVAL_47 = _EVAL_84 & _EVAL_2;
  assign _EVAL_110 = _EVAL_14 & _EVAL_24;
  assign _EVAL_53 = _EVAL_50 & _EVAL_2;
  assign _EVAL_87 = _EVAL_84 & _EVAL_80;
  assign _EVAL_37 = _EVAL_5 == 4'hd;
  assign _EVAL_56 = _EVAL_54 & _EVAL_2;
  assign _EVAL_52 = _EVAL_18 & _EVAL_80;
  assign _EVAL_82 = _EVAL_18 & _EVAL_24;
  assign _EVAL_112 = _EVAL_111 & _EVAL_80;
  assign _EVAL_80 = _EVAL_1;
  assign _EVAL_24 = ~_EVAL_2;
  assign _EVAL_64 = _EVAL_55 & _EVAL_24;
  assign _EVAL_92 = ~_EVAL_80;
  assign _EVAL_103 = _EVAL_21 & _EVAL_24;
  assign _EVAL_90 = _EVAL_74 & _EVAL_80;
  assign _EVAL_20 = _EVAL_10 & _EVAL_24;
  assign _EVAL_39 = _EVAL_84 & _EVAL_24;
  assign _EVAL_32 = _EVAL_13 & _EVAL_80;
  assign _EVAL_104 = _EVAL_37 & _EVAL_24;
  assign _EVAL_40 = _EVAL_59 & _EVAL_2;
  assign _EVAL_77 = _EVAL_21 & _EVAL_2;
  assign _EVAL_55 = _EVAL_5 == 4'h0;
  assign _EVAL_27 = _EVAL_37 & _EVAL_80;
  assign _EVAL_97 = _EVAL_111 & _EVAL_2;
  assign _EVAL_14 = _EVAL_5 == 4'h1;
  assign _EVAL_57 = _EVAL_18 & _EVAL_2;
  assign _EVAL_95 = _EVAL_50 & _EVAL_24;
  assign _EVAL_6 = _EVAL_5 == 4'he;
  assign _EVAL_66 = _EVAL_74 & _EVAL_24;
  assign _EVAL_25 = _EVAL_111 & _EVAL_24;
  assign _EVAL_36 = _EVAL_13 & _EVAL_2;
  assign _EVAL_8 = _EVAL_55 & _EVAL_2;
  assign _EVAL_94 = _EVAL_6 & _EVAL_2;
  assign _EVAL_105 = _EVAL_109 & _EVAL_2;
  always @(posedge _EVAL) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54eb487c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cec7298a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95776544)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6fec0b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bc134fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa49f817)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d494e55a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6e8c898)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af7edd20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb95267)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4063409c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(397043f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c93f6fcb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d997b4fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2f6e18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5f0a6b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b3d24d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6c7c3d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44a67fee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56d5add3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6f7736d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b1b230c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a16adac5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8282d629)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(762d94a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_70 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0a4a287)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19cccdf8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_8 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(564e0447)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9fd1fc89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbd14242)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(240b2c8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61d6fb31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a49a7b2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23209941)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e84c7f70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f1bba4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f39bb7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72ea99fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9354c8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b978e73b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d256f12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6551f21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdbf35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1889f32b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(658e600b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c456feb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8362fc97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f34e1981)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
