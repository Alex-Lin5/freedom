//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_68_assert(
  input  [3:0]  _EVAL,
  input         _EVAL_0,
  input  [11:0] _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [4:0]  _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input  [4:0]  _EVAL_8,
  input         _EVAL_9,
  input  [2:0]  _EVAL_10,
  input  [2:0]  _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input  [2:0]  _EVAL_14
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_15;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire [12:0] _EVAL_23;
  reg [2:0] _EVAL_24;
  wire [3:0] _EVAL_25;
  wire  _EVAL_26;
  wire [4:0] _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire [17:0] _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  reg [4:0] _EVAL_36;
  wire [5:0] _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_44;
  reg [3:0] _EVAL_45;
  wire [12:0] _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  reg [3:0] _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire [3:0] _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire [17:0] _EVAL_62;
  wire  _EVAL_63;
  wire [31:0] _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire [3:0] _EVAL_69;
  wire [17:0] _EVAL_70;
  wire  _EVAL_71;
  wire [4:0] _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire [31:0] _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire [11:0] _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire [5:0] _EVAL_92;
  wire [3:0] _EVAL_93;
  wire [1:0] _EVAL_94;
  wire [12:0] _EVAL_95;
  reg [2:0] _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire [12:0] _EVAL_103;
  wire [17:0] _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire [3:0] _EVAL_108;
  wire  _EVAL_109;
  reg [3:0] _EVAL_110;
  wire [2:0] _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire [17:0] _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire [5:0] _EVAL_119;
  wire [3:0] _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_124;
  wire [3:0] _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  reg [11:0] _EVAL_138;
  wire [17:0] _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire [31:0] _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire [5:0] _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire [3:0] _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  reg [4:0] _EVAL_169;
  wire [31:0] _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire [2:0] _EVAL_174;
  wire [4:0] _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  reg [31:0] _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  reg [3:0] _EVAL_193;
  reg [2:0] _EVAL_194;
  wire  _EVAL_195;
  reg [2:0] _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire [4:0] _EVAL_213;
  wire [1:0] _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire [12:0] _EVAL_230;
  reg [2:0] _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire [17:0] _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire [1:0] _EVAL_240;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire [31:0] _EVAL_246;
  wire [1:0] _EVAL_247;
  reg [17:0] _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire [11:0] _EVAL_256;
  wire  _EVAL_257;
  wire [17:0] _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire [32:0] _EVAL_271;
  wire [3:0] _EVAL_272;
  wire  _EVAL_273;
  wire [3:0] _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_173 = _EVAL_121 | _EVAL_224;
  assign _EVAL_127 = _EVAL_12 & _EVAL_176;
  assign _EVAL_269 = _EVAL_2 & _EVAL_107;
  assign _EVAL_209 = _EVAL_18 & _EVAL_57;
  assign _EVAL_79 = _EVAL_11 == 3'h7;
  assign _EVAL_200 = ~_EVAL_145;
  assign _EVAL_84 = _EVAL_8 == _EVAL_36;
  assign _EVAL_265 = _EVAL_11 == 3'h3;
  assign _EVAL_258 = _EVAL_70 & _EVAL_236;
  assign _EVAL_262 = _EVAL_30 | _EVAL_7;
  assign _EVAL_104 = _EVAL_115 >> _EVAL_4;
  assign _EVAL_254 = ~_EVAL_166;
  assign _EVAL_100 = _EVAL_3 <= 3'h3;
  assign _EVAL_19 = _EVAL_83 | _EVAL_126;
  assign _EVAL_239 = ~_EVAL_34;
  assign _EVAL_187 = _EVAL_14[0];
  assign _EVAL_116 = _EVAL_118 | _EVAL_7;
  assign _EVAL_158 = _EVAL_11[2];
  assign _EVAL_86 = {{6'd0}, _EVAL_152};
  assign _EVAL_237 = ~_EVAL_41;
  assign _EVAL_236 = ~_EVAL_32;
  assign _EVAL_256 = _EVAL_1 & _EVAL_86;
  assign _EVAL_215 = _EVAL_133 | _EVAL_7;
  assign _EVAL_69 = ~_EVAL_108;
  assign _EVAL_38 = _EVAL_219 | _EVAL_141;
  assign _EVAL_210 = _EVAL_11 == 3'h5;
  assign _EVAL_240 = _EVAL_94 | 2'h1;
  assign _EVAL_213 = _EVAL_45 - 4'h1;
  assign _EVAL_267 = ~_EVAL_191;
  assign _EVAL_17 = plusarg_reader_out == 32'h0;
  assign _EVAL_20 = _EVAL_156 == 4'h0;
  assign _EVAL_197 = _EVAL_11 == 3'h0;
  assign _EVAL_26 = _EVAL_117 & _EVAL_157;
  assign _EVAL_163 = _EVAL_3 <= 3'h2;
  assign _EVAL_128 = _EVAL_109 | _EVAL_88;
  assign _EVAL_90 = _EVAL_217 | _EVAL_7;
  assign _EVAL_148 = _EVAL_10[0];
  assign _EVAL_147 = _EVAL_124 & _EVAL_28;
  assign _EVAL_72 = _EVAL_193 - 4'h1;
  assign _EVAL_97 = _EVAL_220 | _EVAL_7;
  assign _EVAL_108 = {_EVAL_208,_EVAL_52,_EVAL_58,_EVAL_216};
  assign _EVAL_125 = _EVAL_213[3:0];
  assign _EVAL_232 = ~_EVAL_160;
  assign _EVAL_140 = ~_EVAL_276;
  assign _EVAL_70 = _EVAL_248 | _EVAL_62;
  assign _EVAL_102 = _EVAL_51 | _EVAL_223;
  assign _EVAL_33 = ~_EVAL_107;
  assign _EVAL_25 = _EVAL_175[3:0];
  assign _EVAL_118 = ~_EVAL_270;
  assign _EVAL_157 = _EVAL_45 == 4'h0;
  assign _EVAL_206 = ~_EVAL_44;
  assign _EVAL_185 = _EVAL_8 == 5'h11;
  assign _EVAL_135 = _EVAL_228 | _EVAL_7;
  assign _EVAL_273 = _EVAL_174 <= 3'h6;
  assign _EVAL_227 = 3'h6 == _EVAL_10;
  assign _EVAL_62 = _EVAL_246[17:0];
  assign _EVAL_126 = _EVAL_4 == 5'h8;
  assign _EVAL_192 = _EVAL_10 <= 3'h6;
  assign _EVAL_175 = _EVAL_110 - 4'h1;
  assign _EVAL_214 = _EVAL_8[4:3];
  assign _EVAL_167 = _EVAL_235 & _EVAL_189;
  assign _EVAL_22 = _EVAL_14 == _EVAL_196;
  assign _EVAL_238 = _EVAL_12 & _EVAL_197;
  assign _EVAL_31 = _EVAL_2 & _EVAL_243;
  assign _EVAL_137 = ~_EVAL_221;
  assign _EVAL_244 = _EVAL_10 == _EVAL_194;
  assign _EVAL_18 = _EVAL_1[1];
  assign _EVAL_80 = _EVAL_202 & _EVAL_61;
  assign _EVAL_149 = _EVAL_202 & _EVAL_129;
  assign _EVAL_46 = _EVAL_230;
  assign _EVAL_41 = _EVAL_155 | _EVAL_7;
  assign _EVAL_77 = ~_EVAL_97;
  assign _EVAL_101 = _EVAL_98 | _EVAL_165;
  assign _EVAL_21 = _EVAL_2 & _EVAL_91;
  assign _EVAL_183 = _EVAL_20 | _EVAL_7;
  assign _EVAL_276 = _EVAL_15 | _EVAL_7;
  assign _EVAL_188 = _EVAL_109 | _EVAL_73;
  assign _EVAL_178 = _EVAL_104[0];
  assign _EVAL_257 = ~_EVAL_245;
  assign _EVAL_268 = |_EVAL_248;
  assign _EVAL_247 = _EVAL_4[4:3];
  assign _EVAL_233 = _EVAL_202 & _EVAL_252;
  assign _EVAL_217 = _EVAL_192 & _EVAL_76;
  assign _EVAL_164 = _EVAL_173 | _EVAL_7;
  assign _EVAL_179 = ~_EVAL_164;
  assign _EVAL_129 = _EVAL_261 & _EVAL_266;
  assign _EVAL_203 = ~_EVAL_106;
  assign _EVAL_61 = _EVAL_18 & _EVAL_266;
  assign _EVAL_205 = _EVAL_11 == _EVAL_231;
  assign _EVAL_40 = _EVAL_244 | _EVAL_7;
  assign _EVAL_48 = _EVAL_67 | _EVAL_7;
  assign _EVAL_224 = _EVAL_8 == 5'h8;
  assign _EVAL_153 = _EVAL_199 | _EVAL_7;
  assign _EVAL_114 = _EVAL_26 & _EVAL_33;
  assign _EVAL_91 = _EVAL_14 == 3'h5;
  assign _EVAL_81 = _EVAL_3 == _EVAL_96;
  assign _EVAL_131 = _EVAL_10 <= 3'h2;
  assign _EVAL_121 = _EVAL_181 | _EVAL_59;
  assign _EVAL_162 = ~_EVAL_158;
  assign _EVAL_63 = _EVAL_3 != 3'h0;
  assign _EVAL_144 = _EVAL_205 | _EVAL_7;
  assign _EVAL_189 = _EVAL_111 <= 3'h6;
  assign _EVAL_35 = _EVAL_63 | _EVAL_7;
  assign _EVAL_107 = _EVAL_14 == 3'h6;
  assign _EVAL_195 = _EVAL_14 == 3'h0;
  assign _EVAL_263 = _EVAL_14 == 3'h1;
  assign _EVAL_223 = _EVAL_184 < plusarg_reader_out;
  assign _EVAL_261 = ~_EVAL_18;
  assign _EVAL_134 = _EVAL_117 & _EVAL_47;
  assign _EVAL_202 = _EVAL_240[0];
  assign _EVAL_50 = ~_EVAL_48;
  assign _EVAL_94 = 2'h1 << _EVAL_148;
  assign _EVAL_88 = _EVAL_260 & _EVAL_261;
  assign _EVAL_220 = _EVAL_3 == 3'h0;
  assign _EVAL_73 = _EVAL_260 & _EVAL_18;
  assign _EVAL_252 = _EVAL_261 & _EVAL_57;
  assign _EVAL_34 = _EVAL_19 | _EVAL_7;
  assign _EVAL_136 = _EVAL_49 == 4'h0;
  assign _EVAL_132 = _EVAL_185 | _EVAL_59;
  assign _EVAL_154 = _EVAL_22 | _EVAL_7;
  assign _EVAL_113 = ~_EVAL_87;
  assign _EVAL_139 = _EVAL_248 >> _EVAL_8;
  assign _EVAL_243 = _EVAL_14 == 3'h2;
  assign _EVAL_176 = _EVAL_11 == 3'h2;
  assign _EVAL_120 = _EVAL_72[3:0];
  assign _EVAL_133 = _EVAL_4 == _EVAL_169;
  assign _EVAL_52 = _EVAL_188 | _EVAL_80;
  assign _EVAL_119 = _EVAL_95[5:0];
  assign _EVAL_85 = _EVAL_2 & _EVAL_211;
  assign _EVAL_65 = ~_EVAL_7;
  assign _EVAL_216 = _EVAL_128 | _EVAL_149;
  assign _EVAL_150 = _EVAL_2 & _EVAL_263;
  assign _EVAL_270 = _EVAL_139[0];
  assign _EVAL_208 = _EVAL_188 | _EVAL_171;
  assign _EVAL_259 = ~_EVAL_161;
  assign _EVAL_201 = _EVAL_11 == 3'h4;
  assign _EVAL_181 = _EVAL_185 | _EVAL_165;
  assign _EVAL_274 = _EVAL_27[3:0];
  assign _EVAL_124 = _EVAL_0 & _EVAL_12;
  assign _EVAL_199 = _EVAL_3 <= 3'h4;
  assign _EVAL_23 = {1'b0,$signed(_EVAL_1)};
  assign _EVAL_117 = _EVAL_6 & _EVAL_2;
  assign _EVAL_83 = _EVAL_38 | _EVAL_167;
  assign _EVAL_28 = _EVAL_193 == 4'h0;
  assign _EVAL_219 = _EVAL_4 == 5'h11;
  assign _EVAL_106 = _EVAL_163 | _EVAL_7;
  assign _EVAL_172 = ~_EVAL_222;
  assign _EVAL_177 = ~_EVAL_215;
  assign _EVAL_92 = _EVAL_103[5:0];
  assign _EVAL_42 = ~_EVAL_136;
  assign _EVAL_207 = _EVAL_12 & _EVAL_151;
  assign _EVAL_146 = _EVAL_271[31:0];
  assign _EVAL_161 = _EVAL_29 | _EVAL_7;
  assign _EVAL_245 = _EVAL_178 | _EVAL_7;
  assign _EVAL_103 = 13'h3f << _EVAL_5;
  assign _EVAL_44 = _EVAL_84 | _EVAL_7;
  assign _EVAL_89 = _EVAL_12 & _EVAL_105;
  assign _EVAL_27 = _EVAL_49 - 4'h1;
  assign _EVAL_246 = _EVAL_147 ? _EVAL_64 : 32'h0;
  assign _EVAL_76 = $signed(_EVAL_46) == 13'sh0;
  assign _EVAL_109 = _EVAL_10 >= 3'h2;
  assign _EVAL_58 = _EVAL_128 | _EVAL_233;
  assign _EVAL_95 = 13'h3f << _EVAL_10;
  assign _EVAL_141 = _EVAL_4 == 5'h10;
  assign _EVAL_165 = _EVAL_8 == 5'h10;
  assign _EVAL_39 = ~_EVAL_262;
  assign _EVAL_53 = _EVAL_37[5:2];
  assign _EVAL_51 = _EVAL_43 | _EVAL_17;
  assign _EVAL_222 = _EVAL_81 | _EVAL_7;
  assign _EVAL_253 = ~_EVAL_116;
  assign _EVAL_130 = _EVAL_5 == _EVAL_24;
  assign _EVAL_250 = _EVAL_124 & _EVAL_136;
  assign _EVAL_156 = _EVAL & _EVAL_69;
  assign _EVAL_198 = _EVAL_12 & _EVAL_201;
  assign _EVAL_191 = _EVAL_100 | _EVAL_7;
  assign _EVAL_15 = _EVAL_1 == _EVAL_138;
  assign _EVAL_56 = _EVAL_249 | _EVAL_7;
  assign _EVAL_112 = _EVAL_124 | _EVAL_117;
  assign _EVAL_212 = ~_EVAL_56;
  assign _EVAL_93 = _EVAL_152[5:2];
  assign _EVAL_271 = _EVAL_184 + 32'h1;
  assign _EVAL_32 = _EVAL_82[17:0];
  assign _EVAL_87 = _EVAL_234 | _EVAL_7;
  assign _EVAL_160 = _EVAL_102 | _EVAL_7;
  assign _EVAL_111 = _EVAL_4[2:0];
  assign _EVAL_43 = ~_EVAL_268;
  assign _EVAL_82 = _EVAL_114 ? _EVAL_170 : 32'h0;
  assign _EVAL_275 = _EVAL_68 | _EVAL_7;
  assign _EVAL_170 = 32'h1 << _EVAL_4;
  assign _EVAL_142 = ~_EVAL_90;
  assign _EVAL_182 = _EVAL_12 & _EVAL_210;
  assign _EVAL_235 = _EVAL_247 == 2'h0;
  assign _EVAL_145 = _EVAL_16 | _EVAL_7;
  assign _EVAL_204 = _EVAL_2 & _EVAL_195;
  assign _EVAL_249 = _EVAL_256 == 12'h0;
  assign _EVAL_171 = _EVAL_202 & _EVAL_209;
  assign _EVAL_60 = ~_EVAL_35;
  assign _EVAL_272 = ~_EVAL;
  assign _EVAL_16 = _EVAL_101 & _EVAL_217;
  assign _EVAL_255 = ~_EVAL_135;
  assign _EVAL_71 = _EVAL_2 & _EVAL_168;
  assign _EVAL_211 = _EVAL_14 == 3'h4;
  assign _EVAL_242 = ~_EVAL_275;
  assign _EVAL_99 = _EVAL_214 == 2'h0;
  assign _EVAL_234 = _EVAL_101 | _EVAL_55;
  assign _EVAL_78 = ~_EVAL_154;
  assign _EVAL_105 = _EVAL_11 == 3'h6;
  assign _EVAL_98 = _EVAL_131 & _EVAL_132;
  assign _EVAL_221 = _EVAL_109 | _EVAL_7;
  assign _EVAL_57 = _EVAL_1[0];
  assign _EVAL_228 = _EVAL_3 <= 3'h1;
  assign _EVAL_190 = ~_EVAL_144;
  assign _EVAL_68 = _EVAL == _EVAL_108;
  assign _EVAL_229 = _EVAL_12 & _EVAL_42;
  assign _EVAL_174 = _EVAL_8[2:0];
  assign _EVAL_230 = $signed(_EVAL_23) & 13'sh1000;
  assign _EVAL_225 = _EVAL_12 & _EVAL_265;
  assign _EVAL_159 = ~_EVAL_153;
  assign _EVAL_226 = _EVAL_12 & _EVAL_79;
  assign _EVAL_30 = _EVAL_272 == 4'h0;
  assign _EVAL_67 = ~_EVAL_9;
  assign _EVAL_151 = _EVAL_11 == 3'h1;
  assign _EVAL_59 = _EVAL_99 & _EVAL_273;
  assign _EVAL_55 = _EVAL_227 & _EVAL_224;
  assign _EVAL_54 = ~_EVAL_183;
  assign _EVAL_186 = ~_EVAL_40;
  assign _EVAL_260 = _EVAL_240[1];
  assign _EVAL_166 = _EVAL_130 | _EVAL_7;
  assign _EVAL_37 = ~_EVAL_92;
  assign _EVAL_266 = ~_EVAL_57;
  assign _EVAL_168 = ~_EVAL_47;
  assign _EVAL_64 = 32'h1 << _EVAL_8;
  assign _EVAL_115 = _EVAL_62 | _EVAL_248;
  assign _EVAL_47 = _EVAL_110 == 4'h0;
  assign _EVAL_155 = _EVAL_14 <= 3'h6;
  assign _EVAL_29 = _EVAL_5 >= 3'h2;
  assign _EVAL_152 = ~_EVAL_119;
  always @(posedge _EVAL_13) begin
    if (_EVAL_134) begin
      _EVAL_24 <= _EVAL_5;
    end
    if (_EVAL_250) begin
      _EVAL_36 <= _EVAL_8;
    end
    if (_EVAL_7) begin
      _EVAL_45 <= 4'h0;
    end else if (_EVAL_117) begin
      if (_EVAL_157) begin
        if (_EVAL_187) begin
          _EVAL_45 <= _EVAL_53;
        end else begin
          _EVAL_45 <= 4'h0;
        end
      end else begin
        _EVAL_45 <= _EVAL_125;
      end
    end
    if (_EVAL_7) begin
      _EVAL_49 <= 4'h0;
    end else if (_EVAL_124) begin
      if (_EVAL_136) begin
        if (_EVAL_162) begin
          _EVAL_49 <= _EVAL_93;
        end else begin
          _EVAL_49 <= 4'h0;
        end
      end else begin
        _EVAL_49 <= _EVAL_274;
      end
    end
    if (_EVAL_250) begin
      _EVAL_96 <= _EVAL_3;
    end
    if (_EVAL_7) begin
      _EVAL_110 <= 4'h0;
    end else if (_EVAL_117) begin
      if (_EVAL_47) begin
        if (_EVAL_187) begin
          _EVAL_110 <= _EVAL_53;
        end else begin
          _EVAL_110 <= 4'h0;
        end
      end else begin
        _EVAL_110 <= _EVAL_25;
      end
    end
    if (_EVAL_250) begin
      _EVAL_138 <= _EVAL_1;
    end
    if (_EVAL_134) begin
      _EVAL_169 <= _EVAL_4;
    end
    if (_EVAL_7) begin
      _EVAL_184 <= 32'h0;
    end else if (_EVAL_112) begin
      _EVAL_184 <= 32'h0;
    end else begin
      _EVAL_184 <= _EVAL_146;
    end
    if (_EVAL_7) begin
      _EVAL_193 <= 4'h0;
    end else if (_EVAL_124) begin
      if (_EVAL_28) begin
        if (_EVAL_162) begin
          _EVAL_193 <= _EVAL_93;
        end else begin
          _EVAL_193 <= 4'h0;
        end
      end else begin
        _EVAL_193 <= _EVAL_120;
      end
    end
    if (_EVAL_250) begin
      _EVAL_194 <= _EVAL_10;
    end
    if (_EVAL_134) begin
      _EVAL_196 <= _EVAL_14;
    end
    if (_EVAL_250) begin
      _EVAL_231 <= _EVAL_11;
    end
    if (_EVAL_7) begin
      _EVAL_248 <= 18'h0;
    end else begin
      _EVAL_248 <= _EVAL_258;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da42291e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26697185)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28bc5df7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3fdfc95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_253) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(920959eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8e514b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ee3bf80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5514d4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed60f264)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7639758)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c3e0eea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bcce211d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ac5a913)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fa7cc01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2db0cd8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3da3a92f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_2 & _EVAL_237) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_255) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6466af0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f96703eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e512437a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c96e8f73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8af2f797)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(491cbc42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a9f035e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53240ec3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bbf44f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad6a3611)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96a5fbbc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c96e8f73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d834082)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ef53847)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54a72cbc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db5c61a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d76848ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc514a3c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(303d585d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bcfabb06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6239728)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33fc1c70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b238c9ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_255) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a076097)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_257) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0517337)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f131d60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bb0c7d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97bd8286)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c54cdb65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb87e12f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aed5fe4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16730d6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_257) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b4c73d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(903e60a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4fc4b89b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7fc275c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4c0816f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38d8f5bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ae00a9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4384e04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(586b7843)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d72467e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b80c3a30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b23a01af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_204 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd42350)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12d9914b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f98f66a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(451fb18c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99af38eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a3d71bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37fd066a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85e7c361)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc031c9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be6cd8f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(355ddd28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b776e3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_253) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d8c6c47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2 & _EVAL_237) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5041fa4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90e61bff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_24 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_36 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_45 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_49 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_96 = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_110 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_138 = _RAND_6[11:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_169 = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_184 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_193 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_194 = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_196 = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_231 = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_248 = _RAND_13[17:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
