//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_30_assert(
  input         _EVAL,
  input  [1:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input  [3:0]  _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [2:0]  _EVAL_9,
  input         _EVAL_10,
  input  [3:0]  _EVAL_11,
  input         _EVAL_12,
  input  [31:0] _EVAL_13
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_14;
  wire [32:0] _EVAL_15;
  wire [31:0] _EVAL_16;
  wire [32:0] _EVAL_17;
  wire [32:0] _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  reg  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire [32:0] _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire [7:0] _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire [7:0] _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire [32:0] _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  reg [7:0] _EVAL_47;
  reg [31:0] _EVAL_48;
  wire  _EVAL_49;
  wire [31:0] _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire [32:0] _EVAL_53;
  wire [8:0] _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire [1:0] _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire [32:0] _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_66;
  wire  _EVAL_67;
  reg  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire [7:0] _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_76;
  reg [3:0] _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire [31:0] _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire [31:0] _EVAL_97;
  reg [7:0] _EVAL_98;
  wire [32:0] _EVAL_99;
  wire [32:0] _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire [32:0] _EVAL_112;
  wire [8:0] _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  reg [2:0] _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire [7:0] _EVAL_128;
  wire  _EVAL_129;
  reg  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire [7:0] _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire [32:0] _EVAL_139;
  wire  _EVAL_140;
  wire [32:0] _EVAL_141;
  wire  _EVAL_142;
  wire [31:0] _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire [32:0] _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  reg [7:0] _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire [7:0] _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  reg [2:0] _EVAL_164;
  wire  _EVAL_165;
  wire [32:0] _EVAL_166;
  wire [32:0] _EVAL_167;
  reg [3:0] _EVAL_168;
  wire  _EVAL_169;
  wire [31:0] _EVAL_170;
  wire  _EVAL_171;
  wire [31:0] _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire [31:0] _EVAL_185;
  wire  _EVAL_186;
  reg [7:0] _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire [32:0] _EVAL_190;
  wire [32:0] _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire [31:0] _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire [8:0] _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  reg [1:0] _EVAL_201;
  wire [32:0] _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_205;
  wire [32:0] _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire [32:0] _EVAL_212;
  wire [7:0] _EVAL_213;
  wire  _EVAL_214;
  wire [8:0] _EVAL_215;
  wire [7:0] _EVAL_216;
  wire [31:0] _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire [1:0] _EVAL_221;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire [32:0] _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire [22:0] _EVAL_233;
  wire  _EVAL_235;
  wire [22:0] _EVAL_236;
  reg [31:0] _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire [32:0] _EVAL_240;
  wire [32:0] _EVAL_241;
  wire  _EVAL_242;
  wire [32:0] _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire [32:0] _EVAL_248;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_27 = _EVAL_125 | _EVAL;
  assign _EVAL_148 = ~_EVAL_107;
  assign _EVAL_84 = ~_EVAL_1;
  assign _EVAL_49 = ~_EVAL_109;
  assign _EVAL_78 = _EVAL_46 | _EVAL_132;
  assign _EVAL_15 = _EVAL_100;
  assign _EVAL_14 = _EVAL_163 & _EVAL_220;
  assign _EVAL_241 = $signed(_EVAL_243) & -33'sh2000;
  assign _EVAL_194 = _EVAL_13 ^ 32'hc000000;
  assign _EVAL_141 = $signed(_EVAL_202) & -33'sh5000;
  assign _EVAL_147 = _EVAL_125 | _EVAL_1;
  assign _EVAL_93 = ~_EVAL_70;
  assign _EVAL_103 = ~_EVAL_186;
  assign _EVAL_132 = plusarg_reader_out == 32'h0;
  assign _EVAL_245 = ~_EVAL_101;
  assign _EVAL_100 = $signed(_EVAL_191) & -33'sh400000;
  assign _EVAL_34 = _EVAL_81 | _EVAL_1;
  assign _EVAL_175 = _EVAL_8 & _EVAL_188;
  assign _EVAL_196 = $signed(_EVAL_53) == 33'sh0;
  assign _EVAL_43 = _EVAL_6 & _EVAL_121;
  assign _EVAL_235 = ~_EVAL_37;
  assign _EVAL_118 = _EVAL_31 | _EVAL_1;
  assign _EVAL_231 = _EVAL_173 | _EVAL_96;
  assign _EVAL_127 = _EVAL_110 | _EVAL_203;
  assign _EVAL_32 = _EVAL_54[7:0];
  assign _EVAL_243 = {1'b0,$signed(_EVAL_16)};
  assign _EVAL_125 = ~_EVAL_10;
  assign _EVAL_227 = $signed(_EVAL_15) == 33'sh0;
  assign _EVAL_85 = _EVAL_9 == 3'h2;
  assign _EVAL_95 = _EVAL_5 <= 3'h6;
  assign _EVAL_137 = _EVAL_40 | _EVAL_1;
  assign _EVAL_92 = |_EVAL_20;
  assign _EVAL_143 = _EVAL_13 & _EVAL_185;
  assign _EVAL_53 = _EVAL_241;
  assign _EVAL_21 = _EVAL_221[0];
  assign _EVAL_63 = _EVAL_112;
  assign _EVAL_22 = ~_EVAL_184;
  assign _EVAL_229 = ~_EVAL_76;
  assign _EVAL_244 = $signed(_EVAL_206) == 33'sh0;
  assign _EVAL_197 = ~_EVAL_71;
  assign _EVAL_202 = {1'b0,$signed(_EVAL_13)};
  assign _EVAL_150 = $signed(_EVAL_99) & -33'sh4000;
  assign _EVAL_55 = _EVAL_8 & _EVAL_171;
  assign _EVAL_121 = _EVAL_5 == 3'h5;
  assign _EVAL_61 = _EVAL_224 | _EVAL_176;
  assign _EVAL_126 = _EVAL_6 & _EVAL_24;
  assign _EVAL_142 = _EVAL_0 != 2'h2;
  assign _EVAL_156 = ~_EVAL_137;
  assign _EVAL_64 = ~_EVAL_200;
  assign _EVAL_89 = _EVAL_5 == 3'h0;
  assign _EVAL_96 = ~_EVAL_92;
  assign _EVAL_169 = ~_EVAL;
  assign _EVAL_186 = _EVAL_25 | _EVAL_1;
  assign _EVAL_177 = ~_EVAL_118;
  assign _EVAL_70 = _EVAL_117 | _EVAL_1;
  assign _EVAL_172 = _EVAL_13 ^ 32'h20000000;
  assign _EVAL_230 = _EVAL_9 == 3'h0;
  assign _EVAL_152 = _EVAL_8 & _EVAL_230;
  assign _EVAL_41 = _EVAL_226;
  assign _EVAL_120 = ~_EVAL_124;
  assign _EVAL_33 = $signed(_EVAL_212) == 33'sh0;
  assign _EVAL_44 = $signed(_EVAL_41) == 33'sh0;
  assign _EVAL_62 = _EVAL_104 & _EVAL_91;
  assign _EVAL_54 = _EVAL_47 - 8'h1;
  assign _EVAL_179 = _EVAL_9 == 3'h7;
  assign _EVAL_57 = _EVAL_14 ? 2'h1 : 2'h0;
  assign _EVAL_25 = _EVAL_4 <= 4'h2;
  assign _EVAL_224 = _EVAL_45 | _EVAL_227;
  assign _EVAL_76 = _EVAL_82 | _EVAL_1;
  assign _EVAL_17 = {1'b0,$signed(_EVAL_172)};
  assign _EVAL_66 = _EVAL_20 | _EVAL_23;
  assign _EVAL_171 = ~_EVAL_67;
  assign _EVAL_214 = _EVAL_48 < plusarg_reader_out;
  assign _EVAL_31 = _EVAL_0 == _EVAL_201;
  assign _EVAL_189 = _EVAL_9 == 3'h5;
  assign _EVAL_80 = ~_EVAL_21;
  assign _EVAL_212 = _EVAL_190;
  assign _EVAL_117 = ~_EVAL_23;
  assign _EVAL_30 = $signed(_EVAL_63) == 33'sh0;
  assign _EVAL_86 = _EVAL_13 ^ 32'h2000000;
  assign _EVAL_238 = $signed(_EVAL_166) == 33'sh0;
  assign _EVAL_88 = _EVAL_5 == _EVAL_164;
  assign _EVAL_50 = _EVAL_13 ^ 32'h3000;
  assign _EVAL_45 = _EVAL_181 | _EVAL_30;
  assign _EVAL_205 = _EVAL_138 | _EVAL_1;
  assign _EVAL_144 = _EVAL_10 == _EVAL_68;
  assign _EVAL_104 = _EVAL_7 & _EVAL_6;
  assign _EVAL_38 = _EVAL_198[7:0];
  assign _EVAL_131 = _EVAL_142 | _EVAL_1;
  assign _EVAL_225 = _EVAL_6 & _EVAL_19;
  assign _EVAL_203 = _EVAL_174 & _EVAL_209;
  assign _EVAL_81 = _EVAL_78 | _EVAL_214;
  assign _EVAL_114 = _EVAL_154 - 8'h1;
  assign _EVAL_167 = {1'b0,$signed(_EVAL_97)};
  assign _EVAL_185 = {{24'd0}, _EVAL_128};
  assign _EVAL_160 = _EVAL_163 | _EVAL_104;
  assign _EVAL_192 = _EVAL_6 & _EVAL_89;
  assign _EVAL_200 = _EVAL_193 | _EVAL_1;
  assign _EVAL_174 = _EVAL_4 <= 4'h6;
  assign _EVAL_217 = _EVAL_29[31:0];
  assign _EVAL_79 = _EVAL_174 & _EVAL_195;
  assign _EVAL_165 = _EVAL_144 | _EVAL_1;
  assign _EVAL_82 = _EVAL_4 == _EVAL_168;
  assign _EVAL_232 = _EVAL_5 == 3'h1;
  assign _EVAL_162 = _EVAL_8 & _EVAL_146;
  assign _EVAL_138 = _EVAL_143 == 32'h0;
  assign _EVAL_20 = _EVAL_57[0];
  assign _EVAL_163 = _EVAL_3 & _EVAL_8;
  assign _EVAL_136 = _EVAL_0 == 2'h0;
  assign _EVAL_102 = ~_EVAL_147;
  assign _EVAL_91 = _EVAL_47 == 8'h0;
  assign _EVAL_40 = _EVAL_110 | _EVAL_79;
  assign _EVAL_74 = ~_EVAL_205;
  assign _EVAL_210 = ~_EVAL_218;
  assign _EVAL_107 = _EVAL_94 | _EVAL_1;
  assign _EVAL_206 = _EVAL_150;
  assign _EVAL_240 = _EVAL_248;
  assign _EVAL_112 = $signed(_EVAL_18) & -33'sh10000;
  assign _EVAL_18 = {1'b0,$signed(_EVAL_86)};
  assign _EVAL_246 = _EVAL_136 | _EVAL_1;
  assign _EVAL_52 = ~_EVAL_131;
  assign _EVAL_182 = _EVAL_6 & _EVAL_232;
  assign _EVAL_140 = _EVAL_169 | _EVAL_1;
  assign _EVAL_191 = {1'b0,$signed(_EVAL_194)};
  assign _EVAL_199 = _EVAL_231 | _EVAL_1;
  assign _EVAL_133 = ~_EVAL_159;
  assign _EVAL_94 = _EVAL_11 == _EVAL_77;
  assign _EVAL_135 = _EVAL_9 == 3'h4;
  assign _EVAL_123 = _EVAL_27 | _EVAL_1;
  assign _EVAL_219 = _EVAL_9 == 3'h3;
  assign _EVAL_170 = _EVAL_13 ^ 32'h80000000;
  assign _EVAL_24 = _EVAL_5 == 3'h6;
  assign _EVAL_58 = _EVAL_66 | _EVAL_1;
  assign _EVAL_111 = _EVAL_23 | _EVAL_20;
  assign _EVAL_180 = _EVAL_8 & _EVAL_179;
  assign _EVAL_173 = _EVAL_20 != _EVAL_21;
  assign _EVAL_124 = _EVAL_95 | _EVAL_1;
  assign _EVAL_248 = $signed(_EVAL_17) & -33'sh2000;
  assign _EVAL_108 = _EVAL_0 <= 2'h2;
  assign _EVAL_90 = _EVAL_183 & _EVAL_36;
  assign _EVAL_101 = _EVAL_88 | _EVAL_1;
  assign _EVAL_42 = ~_EVAL_123;
  assign _EVAL_145 = ~_EVAL_58;
  assign _EVAL_99 = {1'b0,$signed(_EVAL_170)};
  assign _EVAL_190 = $signed(_EVAL_139) & -33'sh1000;
  assign _EVAL_56 = _EVAL_5[0];
  assign _EVAL_73 = _EVAL_233[7:0];
  assign _EVAL_134 = ~_EVAL_165;
  assign _EVAL_105 = _EVAL_116 | _EVAL_1;
  assign _EVAL_146 = _EVAL_9 == 3'h1;
  assign _EVAL_128 = ~_EVAL_73;
  assign _EVAL_106 = _EVAL_8 & _EVAL_85;
  assign _EVAL_184 = _EVAL_9[2];
  assign _EVAL_181 = _EVAL_238 | _EVAL_44;
  assign _EVAL_36 = ~_EVAL_24;
  assign _EVAL_159 = _EVAL_236[7:0];
  assign _EVAL_119 = ~_EVAL_228;
  assign _EVAL_198 = _EVAL_98 - 8'h1;
  assign _EVAL_208 = ~_EVAL_246;
  assign _EVAL_220 = _EVAL_154 == 8'h0;
  assign _EVAL_209 = _EVAL_176 | _EVAL_196;
  assign _EVAL_166 = _EVAL_141;
  assign _EVAL_26 = ~_EVAL_91;
  assign _EVAL_216 = _EVAL_114[7:0];
  assign _EVAL_176 = $signed(_EVAL_240) == 33'sh0;
  assign _EVAL_60 = _EVAL_8 & _EVAL_219;
  assign _EVAL_183 = _EVAL_104 & _EVAL_35;
  assign _EVAL_178 = ~_EVAL_105;
  assign _EVAL_16 = _EVAL_13 ^ 32'h40000000;
  assign _EVAL_247 = _EVAL_61 | _EVAL_196;
  assign _EVAL_233 = 23'hff << _EVAL_4;
  assign _EVAL_151 = ~_EVAL_140;
  assign _EVAL_19 = _EVAL_5 == 3'h4;
  assign _EVAL_228 = _EVAL_127 | _EVAL_1;
  assign _EVAL_129 = _EVAL_4 <= 4'h8;
  assign _EVAL_213 = _EVAL_215[7:0];
  assign _EVAL_157 = _EVAL_8 & _EVAL_189;
  assign _EVAL_155 = _EVAL_6 & _EVAL_26;
  assign _EVAL_37 = _EVAL_207 | _EVAL_1;
  assign _EVAL_115 = |_EVAL_23;
  assign _EVAL_195 = _EVAL_224 | _EVAL_244;
  assign _EVAL_46 = ~_EVAL_115;
  assign _EVAL_226 = $signed(_EVAL_167) & -33'sh4000;
  assign _EVAL_83 = _EVAL_111 & _EVAL_80;
  assign _EVAL_218 = _EVAL_108 | _EVAL_1;
  assign _EVAL_97 = _EVAL_13 ^ 32'h1800000;
  assign _EVAL_69 = _EVAL_247 | _EVAL_244;
  assign _EVAL_35 = _EVAL_98 == 8'h0;
  assign _EVAL_139 = {1'b0,$signed(_EVAL_50)};
  assign _EVAL_71 = _EVAL_72 | _EVAL_1;
  assign _EVAL_109 = _EVAL_59 | _EVAL_1;
  assign _EVAL_211 = _EVAL_8 & _EVAL_135;
  assign _EVAL_51 = _EVAL_174 & _EVAL_69;
  assign _EVAL_116 = _EVAL_12 == _EVAL_130;
  assign _EVAL_215 = _EVAL_187 - 8'h1;
  assign _EVAL_242 = ~_EVAL_34;
  assign _EVAL_239 = ~_EVAL_199;
  assign _EVAL_236 = 23'hff << _EVAL_11;
  assign _EVAL_110 = _EVAL_129 & _EVAL_33;
  assign _EVAL_161 = _EVAL_5 == 3'h2;
  assign _EVAL_87 = _EVAL_163 & _EVAL_67;
  assign _EVAL_207 = _EVAL_25 & _EVAL_59;
  assign _EVAL_188 = _EVAL_9 == 3'h6;
  assign _EVAL_29 = _EVAL_48 + 32'h1;
  assign _EVAL_221 = _EVAL_90 ? 2'h1 : 2'h0;
  assign _EVAL_67 = _EVAL_187 == 8'h0;
  assign _EVAL_193 = _EVAL_13 == _EVAL_237;
  assign _EVAL_72 = _EVAL_9 == _EVAL_122;
  assign _EVAL_39 = _EVAL_6 & _EVAL_161;
  assign _EVAL_59 = _EVAL_110 | _EVAL_51;
  always @(posedge _EVAL_2) begin
    if (_EVAL_1) begin
      _EVAL_23 <= 1'h0;
    end else begin
      _EVAL_23 <= _EVAL_83;
    end
    if (_EVAL_1) begin
      _EVAL_47 <= 8'h0;
    end else if (_EVAL_104) begin
      if (_EVAL_91) begin
        if (_EVAL_56) begin
          _EVAL_47 <= _EVAL_133;
        end else begin
          _EVAL_47 <= 8'h0;
        end
      end else begin
        _EVAL_47 <= _EVAL_32;
      end
    end
    if (_EVAL_1) begin
      _EVAL_48 <= 32'h0;
    end else if (_EVAL_160) begin
      _EVAL_48 <= 32'h0;
    end else begin
      _EVAL_48 <= _EVAL_217;
    end
    if (_EVAL_62) begin
      _EVAL_68 <= _EVAL_10;
    end
    if (_EVAL_62) begin
      _EVAL_77 <= _EVAL_11;
    end
    if (_EVAL_1) begin
      _EVAL_98 <= 8'h0;
    end else if (_EVAL_104) begin
      if (_EVAL_35) begin
        if (_EVAL_56) begin
          _EVAL_98 <= _EVAL_133;
        end else begin
          _EVAL_98 <= 8'h0;
        end
      end else begin
        _EVAL_98 <= _EVAL_38;
      end
    end
    if (_EVAL_87) begin
      _EVAL_122 <= _EVAL_9;
    end
    if (_EVAL_62) begin
      _EVAL_130 <= _EVAL_12;
    end
    if (_EVAL_1) begin
      _EVAL_154 <= 8'h0;
    end else if (_EVAL_163) begin
      if (_EVAL_220) begin
        if (_EVAL_22) begin
          _EVAL_154 <= _EVAL_128;
        end else begin
          _EVAL_154 <= 8'h0;
        end
      end else begin
        _EVAL_154 <= _EVAL_216;
      end
    end
    if (_EVAL_62) begin
      _EVAL_164 <= _EVAL_5;
    end
    if (_EVAL_87) begin
      _EVAL_168 <= _EVAL_4;
    end
    if (_EVAL_1) begin
      _EVAL_187 <= 8'h0;
    end else if (_EVAL_163) begin
      if (_EVAL_67) begin
        if (_EVAL_22) begin
          _EVAL_187 <= _EVAL_128;
        end else begin
          _EVAL_187 <= 8'h0;
        end
      end else begin
        _EVAL_187 <= _EVAL_213;
      end
    end
    if (_EVAL_62) begin
      _EVAL_201 <= _EVAL_0;
    end
    if (_EVAL_87) begin
      _EVAL_237 <= _EVAL_13;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2231e4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1eb984bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d020a1b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4772d1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34e02f82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d355e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a9a0d71)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78c69d88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91b40da1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a6739d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94b16906)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10a28220)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce54e693)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84679890)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a866a24e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84303985)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_145) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d42b0ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa844a35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(104af1fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(584bc9a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c33d84fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_208) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f01adf64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(967a339b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6f9a055)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_208) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a356462b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(858e0eee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46373c55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9de88409)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb09a648)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_208) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(592a86e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f206eaf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f2e1599)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad417e92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b556e56a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e0ce2e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d321d3f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_208) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_208) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3523e111)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4fb71a7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_208) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65f2828d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94b16906)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54af0018)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d57a52ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60760135)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6efe613d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb224472)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(961a162)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ec886d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_208) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4ca392f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d57937ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d37f3e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63426212)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_208) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc5d6cb2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_23 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_47 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_48 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_68 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_77 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_98 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_122 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_130 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_154 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_164 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_168 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_187 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_201 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_237 = _RAND_13[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
