//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_85_assert(
  input  [4:0]  _EVAL,
  input  [2:0]  _EVAL_0,
  input         _EVAL_1,
  input  [1:0]  _EVAL_2,
  input  [4:0]  _EVAL_3,
  input  [2:0]  _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  input         _EVAL_8,
  input  [2:0]  _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input  [29:0] _EVAL_16,
  input         _EVAL_17,
  input  [3:0]  _EVAL_18
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  reg [2:0] _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire [32:0] _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  reg [3:0] _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire [17:0] _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  reg [1:0] _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire [30:0] _EVAL_61;
  reg  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  reg [3:0] _EVAL_69;
  wire  _EVAL_70;
  wire [3:0] _EVAL_71;
  wire [5:0] _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  reg [2:0] _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire [3:0] _EVAL_89;
  wire  _EVAL_90;
  wire [3:0] _EVAL_91;
  wire [31:0] _EVAL_92;
  wire  _EVAL_93;
  wire [29:0] _EVAL_94;
  wire [12:0] _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire [4:0] _EVAL_115;
  reg  _EVAL_116;
  wire [30:0] _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  reg [2:0] _EVAL_120;
  wire  _EVAL_121;
  wire [17:0] _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire [31:0] _EVAL_125;
  wire  _EVAL_126;
  wire [2:0] _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire [4:0] _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire [3:0] _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire [3:0] _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire [1:0] _EVAL_154;
  wire  _EVAL_155;
  wire [31:0] _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire [3:0] _EVAL_159;
  wire [1:0] _EVAL_160;
  wire  _EVAL_161;
  wire [31:0] plusarg_reader_out;
  wire [17:0] _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  reg [2:0] _EVAL_165;
  wire  _EVAL_166;
  reg [17:0] _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire [3:0] _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire [31:0] _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  reg [3:0] _EVAL_182;
  wire [3:0] _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire [17:0] _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire [5:0] _EVAL_201;
  wire [3:0] _EVAL_202;
  wire [29:0] _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  reg [31:0] _EVAL_207;
  wire [17:0] _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire [1:0] _EVAL_222;
  wire  _EVAL_223;
  wire [4:0] _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire [17:0] _EVAL_236;
  wire  _EVAL_238;
  wire  _EVAL_239;
  reg [4:0] _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire [31:0] _EVAL_244;
  wire [2:0] _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire [17:0] _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire [1:0] _EVAL_257;
  wire [5:0] _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  reg [3:0] _EVAL_273;
  wire  _EVAL_274;
  wire [30:0] _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire  _EVAL_280;
  wire [12:0] _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire [4:0] _EVAL_286;
  reg [29:0] _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire [5:0] _EVAL_293;
  wire [17:0] _EVAL_294;
  wire  _EVAL_295;
  wire  _EVAL_296;
  wire [29:0] _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire [3:0] _EVAL_301;
  wire  _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_308;
  wire  _EVAL_309;
  wire  _EVAL_310;
  wire  _EVAL_311;
  wire  _EVAL_312;
  reg [4:0] _EVAL_313;
  wire  _EVAL_314;
  reg [2:0] _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_317;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_274 = _EVAL_257 == 2'h0;
  assign _EVAL_89 = _EVAL_286[3:0];
  assign _EVAL_36 = ~_EVAL_270;
  assign _EVAL_142 = _EVAL_3 == 5'h8;
  assign _EVAL_193 = _EVAL_9 == 3'h5;
  assign _EVAL_244 = _EVAL_253 ? _EVAL_125 : 32'h0;
  assign _EVAL_60 = ~_EVAL_97;
  assign _EVAL_21 = _EVAL_194 | _EVAL_12;
  assign _EVAL_264 = ~_EVAL_13;
  assign _EVAL_204 = _EVAL_197 | _EVAL_271;
  assign _EVAL_115 = _EVAL_69 - 4'h1;
  assign _EVAL_43 = _EVAL_148 | _EVAL_12;
  assign _EVAL_46 = ~_EVAL_73;
  assign _EVAL_33 = _EVAL_294 != _EVAL_162;
  assign _EVAL_177 = ~_EVAL_241;
  assign _EVAL_215 = ~_EVAL_126;
  assign _EVAL_157 = _EVAL_106 | _EVAL_12;
  assign _EVAL_239 = _EVAL_0[0];
  assign _EVAL_171 = _EVAL_37 | _EVAL_12;
  assign _EVAL_191 = _EVAL_167 >> _EVAL_3;
  assign _EVAL_312 = _EVAL_172 | _EVAL_12;
  assign _EVAL_102 = $signed(_EVAL_117) == 31'sh0;
  assign _EVAL_168 = _EVAL_6 & _EVAL_1;
  assign _EVAL_155 = ~_EVAL_196;
  assign _EVAL_146 = _EVAL_63 | _EVAL_295;
  assign _EVAL_32 = _EVAL_41 == 4'h0;
  assign _EVAL_109 = _EVAL_2 == _EVAL_57;
  assign _EVAL_252 = _EVAL_101 & _EVAL_263;
  assign _EVAL_230 = _EVAL_50 | _EVAL_133;
  assign _EVAL_199 = _EVAL_5 <= 3'h2;
  assign _EVAL_134 = _EVAL_8 & _EVAL_17;
  assign _EVAL_251 = _EVAL_294 | _EVAL_167;
  assign _EVAL_192 = _EVAL_0 >= 3'h2;
  assign _EVAL_133 = _EVAL_3 == 5'h10;
  assign _EVAL_263 = _EVAL_272 & _EVAL_139;
  assign _EVAL_106 = ~_EVAL_14;
  assign _EVAL_85 = _EVAL_7 == _EVAL_120;
  assign _EVAL_254 = ~_EVAL_206;
  assign _EVAL_301 = _EVAL_224[3:0];
  assign _EVAL_61 = $signed(_EVAL_275) & -31'sh2000;
  assign _EVAL_38 = _EVAL_230 | _EVAL_289;
  assign _EVAL_190 = _EVAL_199 | _EVAL_12;
  assign _EVAL_74 = |_EVAL_294;
  assign _EVAL_310 = _EVAL_17 & _EVAL_166;
  assign _EVAL_245 = _EVAL[2:0];
  assign _EVAL_216 = _EVAL_5 == _EVAL_78;
  assign _EVAL_92 = _EVAL_198 ? _EVAL_156 : 32'h0;
  assign _EVAL_242 = _EVAL_17 & _EVAL_29;
  assign _EVAL_280 = _EVAL_17 & _EVAL_247;
  assign _EVAL_292 = _EVAL_75 | _EVAL_12;
  assign _EVAL_121 = _EVAL_33 | _EVAL_26;
  assign _EVAL_151 = ~_EVAL_65;
  assign _EVAL_73 = _EVAL_226 | _EVAL_12;
  assign _EVAL_317 = _EVAL_168 & _EVAL_220;
  assign _EVAL_118 = _EVAL_189 | _EVAL_12;
  assign _EVAL_261 = _EVAL == _EVAL_240;
  assign _EVAL_197 = _EVAL_192 | _EVAL_179;
  assign _EVAL_163 = _EVAL_127 <= 3'h6;
  assign _EVAL_298 = _EVAL_106 | _EVAL_13;
  assign _EVAL_232 = _EVAL_3 == _EVAL_313;
  assign _EVAL_210 = _EVAL_146 | _EVAL_12;
  assign _EVAL_52 = ~_EVAL_76;
  assign _EVAL_198 = _EVAL_317 & _EVAL_39;
  assign _EVAL_218 = _EVAL_272 & _EVAL_143;
  assign _EVAL_260 = _EVAL_134 & _EVAL_49;
  assign _EVAL_200 = ~_EVAL_267;
  assign _EVAL_70 = ~_EVAL_98;
  assign _EVAL_150 = {_EVAL_149,_EVAL_204,_EVAL_153,_EVAL_77};
  assign _EVAL_66 = _EVAL_85 | _EVAL_12;
  assign _EVAL_47 = _EVAL_207 < plusarg_reader_out;
  assign _EVAL_101 = _EVAL_222[0];
  assign _EVAL_138 = _EVAL_9 == 3'h6;
  assign _EVAL_217 = ~_EVAL_212;
  assign _EVAL_136 = ~_EVAL_157;
  assign _EVAL_145 = _EVAL_264 | _EVAL_12;
  assign _EVAL_156 = 32'h1 << _EVAL;
  assign _EVAL_309 = _EVAL_1 & _EVAL_243;
  assign _EVAL_279 = ~_EVAL_265;
  assign _EVAL_169 = _EVAL_5 <= 3'h1;
  assign _EVAL_44 = ~_EVAL_228;
  assign _EVAL_188 = ~_EVAL_238;
  assign _EVAL_214 = ~_EVAL_312;
  assign _EVAL_42 = _EVAL_1 & _EVAL_195;
  assign _EVAL_94 = _EVAL_16 ^ 30'h20000000;
  assign _EVAL_306 = ~_EVAL_19;
  assign _EVAL_294 = _EVAL_244[17:0];
  assign _EVAL_122 = _EVAL_251 >> _EVAL;
  assign _EVAL_241 = _EVAL_216 | _EVAL_12;
  assign _EVAL_270 = _EVAL_7[2];
  assign _EVAL_205 = _EVAL_1 & _EVAL_305;
  assign _EVAL_119 = _EVAL_14 == _EVAL_62;
  assign _EVAL_255 = _EVAL_7 == 3'h1;
  assign _EVAL_114 = _EVAL_18 == _EVAL_150;
  assign _EVAL_76 = _EVAL_58 | _EVAL_12;
  assign _EVAL_113 = _EVAL_266 | _EVAL_124;
  assign _EVAL_84 = _EVAL_5 == 3'h0;
  assign _EVAL_286 = _EVAL_182 - 4'h1;
  assign _EVAL_233 = ~_EVAL_288;
  assign _EVAL_126 = _EVAL_284 | _EVAL_12;
  assign _EVAL_51 = _EVAL_1 & _EVAL_110;
  assign _EVAL_297 = {{24'd0}, _EVAL_293};
  assign _EVAL_299 = ~_EVAL_66;
  assign _EVAL_135 = _EVAL_87 & _EVAL_143;
  assign _EVAL_24 = ~_EVAL_107;
  assign _EVAL_111 = ~_EVAL_99;
  assign _EVAL_128 = _EVAL_16 == _EVAL_287;
  assign _EVAL_224 = _EVAL_41 - 4'h1;
  assign _EVAL_249 = _EVAL_5 <= 3'h3;
  assign _EVAL_222 = _EVAL_154 | 2'h1;
  assign _EVAL_55 = _EVAL_160 == 2'h0;
  assign _EVAL_267 = |_EVAL_167;
  assign _EVAL_148 = _EVAL_11 == _EVAL_116;
  assign _EVAL_160 = _EVAL_3[4:3];
  assign _EVAL_28 = _EVAL_17 & _EVAL_67;
  assign _EVAL_49 = _EVAL_182 == 4'h0;
  assign _EVAL_144 = _EVAL_248 | _EVAL_12;
  assign _EVAL_203 = _EVAL_16 & _EVAL_297;
  assign _EVAL_276 = _EVAL_101 & _EVAL_135;
  assign _EVAL_149 = _EVAL_197 | _EVAL_252;
  assign _EVAL_107 = _EVAL_83 | _EVAL_12;
  assign _EVAL_68 = ~_EVAL_190;
  assign _EVAL_37 = _EVAL_122[0];
  assign _EVAL_19 = _EVAL_64 | _EVAL_12;
  assign _EVAL_225 = plusarg_reader_out == 32'h0;
  assign _EVAL_202 = _EVAL_18 & _EVAL_71;
  assign _EVAL_265 = _EVAL_249 | _EVAL_12;
  assign _EVAL_262 = ~_EVAL_314;
  assign _EVAL_93 = ~_EVAL_316;
  assign _EVAL_175 = _EVAL_123 | _EVAL_12;
  assign _EVAL_27 = _EVAL_222[1];
  assign _EVAL_277 = _EVAL_269 & _EVAL_235;
  assign _EVAL_246 = _EVAL_53 | _EVAL_47;
  assign _EVAL_54 = _EVAL_7 == 3'h5;
  assign _EVAL_91 = _EVAL_132[3:0];
  assign _EVAL_212 = _EVAL_109 | _EVAL_12;
  assign _EVAL_79 = _EVAL_17 & _EVAL_80;
  assign _EVAL_247 = _EVAL_7 == 3'h7;
  assign _EVAL_289 = _EVAL_55 & _EVAL_163;
  assign _EVAL_266 = _EVAL_234 | _EVAL_285;
  assign _EVAL_293 = ~_EVAL_258;
  assign _EVAL_316 = _EVAL_161 | _EVAL_12;
  assign _EVAL_31 = _EVAL_256 & _EVAL_102;
  assign _EVAL_303 = _EVAL_141 | _EVAL_12;
  assign _EVAL_159 = _EVAL_115[3:0];
  assign _EVAL_29 = _EVAL_7 == 3'h2;
  assign _EVAL_40 = ~_EVAL_12;
  assign _EVAL_234 = _EVAL == 5'h11;
  assign _EVAL_208 = ~_EVAL_162;
  assign _EVAL_123 = _EVAL_4 >= 3'h2;
  assign _EVAL_161 = _EVAL_9 == _EVAL_165;
  assign _EVAL_117 = _EVAL_61;
  assign _EVAL_75 = _EVAL_2 <= 2'h2;
  assign _EVAL_213 = ~_EVAL_43;
  assign _EVAL_127 = _EVAL_3[2:0];
  assign _EVAL_181 = _EVAL_202 == 4'h0;
  assign _EVAL_86 = _EVAL_168 & _EVAL_296;
  assign _EVAL_26 = ~_EVAL_74;
  assign _EVAL_184 = ~_EVAL_18;
  assign _EVAL_132 = _EVAL_273 - 4'h1;
  assign _EVAL_223 = ~_EVAL_118;
  assign _EVAL_147 = _EVAL_245 <= 3'h6;
  assign _EVAL_295 = _EVAL_104 & _EVAL_142;
  assign _EVAL_228 = _EVAL_232 | _EVAL_12;
  assign _EVAL_96 = ~_EVAL_131;
  assign _EVAL_288 = _EVAL_31 | _EVAL_12;
  assign _EVAL_99 = _EVAL_84 | _EVAL_12;
  assign _EVAL_256 = _EVAL_0 <= 3'h6;
  assign _EVAL_35 = ~_EVAL_129;
  assign _EVAL_174 = _EVAL_293[5:2];
  assign _EVAL_296 = _EVAL_273 == 4'h0;
  assign _EVAL_112 = _EVAL_9[0];
  assign _EVAL_201 = ~_EVAL_72;
  assign _EVAL_271 = _EVAL_101 & _EVAL_218;
  assign _EVAL_125 = 32'h1 << _EVAL_3;
  assign _EVAL_164 = _EVAL == 5'h8;
  assign _EVAL_278 = ~_EVAL_185;
  assign _EVAL_83 = ~_EVAL_82;
  assign _EVAL_281 = 13'h3f << _EVAL_0;
  assign _EVAL_67 = ~_EVAL_49;
  assign _EVAL_275 = {1'b0,$signed(_EVAL_94)};
  assign _EVAL_141 = _EVAL_5 != 3'h0;
  assign _EVAL_185 = _EVAL_298 | _EVAL_12;
  assign _EVAL_87 = ~_EVAL_272;
  assign _EVAL_97 = _EVAL_180 | _EVAL_12;
  assign _EVAL_285 = _EVAL == 5'h10;
  assign _EVAL_243 = ~_EVAL_296;
  assign _EVAL_302 = _EVAL_1 & _EVAL_193;
  assign _EVAL_259 = ~_EVAL_210;
  assign _EVAL_250 = ~_EVAL_175;
  assign _EVAL_291 = _EVAL_169 | _EVAL_12;
  assign _EVAL_45 = _EVAL_167 | _EVAL_294;
  assign _EVAL_82 = _EVAL_191[0];
  assign _EVAL_194 = _EVAL_184 == 4'h0;
  assign _EVAL_248 = _EVAL_5 <= 3'h4;
  assign _EVAL_104 = 3'h6 == _EVAL_0;
  assign _EVAL_282 = ~_EVAL_25;
  assign _EVAL_152 = _EVAL_2 == 2'h0;
  assign _EVAL_153 = _EVAL_130 | _EVAL_186;
  assign _EVAL_56 = _EVAL_87 & _EVAL_139;
  assign _EVAL_80 = _EVAL_7 == 3'h6;
  assign _EVAL_65 = _EVAL_152 | _EVAL_12;
  assign _EVAL_231 = ~_EVAL_303;
  assign _EVAL_206 = _EVAL_128 | _EVAL_12;
  assign _EVAL_235 = _EVAL_50 | _EVAL_289;
  assign _EVAL_258 = _EVAL_281[5:0];
  assign _EVAL_305 = _EVAL_9 == 3'h1;
  assign _EVAL_22 = _EVAL_7 == 3'h0;
  assign _EVAL_129 = _EVAL_119 | _EVAL_12;
  assign _EVAL_257 = _EVAL[4:3];
  assign _EVAL_64 = _EVAL_203 == 30'h0;
  assign _EVAL_180 = _EVAL_0 == _EVAL_23;
  assign _EVAL_34 = _EVAL_207 + 32'h1;
  assign _EVAL_300 = ~_EVAL_145;
  assign _EVAL_25 = _EVAL_261 | _EVAL_12;
  assign _EVAL_311 = _EVAL_1 & _EVAL_138;
  assign _EVAL_130 = _EVAL_192 | _EVAL_304;
  assign _EVAL_100 = _EVAL_113 | _EVAL_164;
  assign _EVAL_71 = ~_EVAL_150;
  assign _EVAL_283 = ~_EVAL_144;
  assign _EVAL_195 = _EVAL_9 == 3'h4;
  assign _EVAL_143 = ~_EVAL_139;
  assign _EVAL_229 = _EVAL_17 & _EVAL_255;
  assign _EVAL_90 = _EVAL_17 & _EVAL_105;
  assign _EVAL_98 = _EVAL_181 | _EVAL_12;
  assign _EVAL_162 = _EVAL_92[17:0];
  assign _EVAL_272 = _EVAL_16[1];
  assign _EVAL_140 = _EVAL_201[5:2];
  assign _EVAL_105 = _EVAL_7 == 3'h4;
  assign _EVAL_20 = ~_EVAL_292;
  assign _EVAL_77 = _EVAL_130 | _EVAL_276;
  assign _EVAL_179 = _EVAL_27 & _EVAL_272;
  assign _EVAL_173 = ~_EVAL_176;
  assign _EVAL_131 = _EVAL_48 | _EVAL_12;
  assign _EVAL_63 = _EVAL_277 | _EVAL_133;
  assign _EVAL_219 = ~_EVAL_291;
  assign _EVAL_189 = _EVAL_38 | _EVAL_142;
  assign _EVAL_59 = _EVAL_246 | _EVAL_12;
  assign _EVAL_50 = _EVAL_3 == 5'h11;
  assign _EVAL_236 = _EVAL_45 & _EVAL_208;
  assign _EVAL_110 = _EVAL_9 == 3'h2;
  assign _EVAL_284 = _EVAL_9 <= 3'h6;
  assign _EVAL_304 = _EVAL_27 & _EVAL_87;
  assign _EVAL_308 = _EVAL_17 & _EVAL_54;
  assign _EVAL_176 = _EVAL_100 | _EVAL_12;
  assign _EVAL_39 = ~_EVAL_138;
  assign _EVAL_58 = _EVAL_63 & _EVAL_31;
  assign _EVAL_268 = _EVAL_9 == 3'h0;
  assign _EVAL_72 = _EVAL_95[5:0];
  assign _EVAL_95 = 13'h3f << _EVAL_4;
  assign _EVAL_238 = _EVAL_192 | _EVAL_12;
  assign _EVAL_154 = 2'h1 << _EVAL_239;
  assign _EVAL_186 = _EVAL_101 & _EVAL_56;
  assign _EVAL_172 = _EVAL_2 != 2'h2;
  assign _EVAL_314 = _EVAL_121 | _EVAL_12;
  assign _EVAL_124 = _EVAL_274 & _EVAL_147;
  assign _EVAL_103 = _EVAL_17 & _EVAL_22;
  assign _EVAL_227 = ~_EVAL_171;
  assign _EVAL_196 = _EVAL_114 | _EVAL_12;
  assign _EVAL_269 = _EVAL_0 <= 3'h2;
  assign _EVAL_178 = _EVAL_34[31:0];
  assign _EVAL_253 = _EVAL_134 & _EVAL_32;
  assign _EVAL_139 = _EVAL_16[0];
  assign _EVAL_158 = _EVAL_134 | _EVAL_168;
  assign _EVAL_221 = ~_EVAL_59;
  assign _EVAL_220 = _EVAL_69 == 4'h0;
  assign _EVAL_226 = ~_EVAL_10;
  assign _EVAL_137 = _EVAL_1 & _EVAL_268;
  assign _EVAL_209 = ~_EVAL_21;
  assign _EVAL_48 = _EVAL_4 == _EVAL_315;
  assign _EVAL_166 = _EVAL_7 == 3'h3;
  assign _EVAL_53 = _EVAL_200 | _EVAL_225;
  always @(posedge _EVAL_15) begin
    if (_EVAL_260) begin
      _EVAL_23 <= _EVAL_0;
    end
    if (_EVAL_12) begin
      _EVAL_41 <= 4'h0;
    end else if (_EVAL_134) begin
      if (_EVAL_32) begin
        if (_EVAL_36) begin
          _EVAL_41 <= _EVAL_174;
        end else begin
          _EVAL_41 <= 4'h0;
        end
      end else begin
        _EVAL_41 <= _EVAL_301;
      end
    end
    if (_EVAL_86) begin
      _EVAL_57 <= _EVAL_2;
    end
    if (_EVAL_86) begin
      _EVAL_62 <= _EVAL_14;
    end
    if (_EVAL_12) begin
      _EVAL_69 <= 4'h0;
    end else if (_EVAL_168) begin
      if (_EVAL_220) begin
        if (_EVAL_112) begin
          _EVAL_69 <= _EVAL_140;
        end else begin
          _EVAL_69 <= 4'h0;
        end
      end else begin
        _EVAL_69 <= _EVAL_159;
      end
    end
    if (_EVAL_260) begin
      _EVAL_78 <= _EVAL_5;
    end
    if (_EVAL_86) begin
      _EVAL_116 <= _EVAL_11;
    end
    if (_EVAL_260) begin
      _EVAL_120 <= _EVAL_7;
    end
    if (_EVAL_86) begin
      _EVAL_165 <= _EVAL_9;
    end
    if (_EVAL_12) begin
      _EVAL_167 <= 18'h0;
    end else begin
      _EVAL_167 <= _EVAL_236;
    end
    if (_EVAL_12) begin
      _EVAL_182 <= 4'h0;
    end else if (_EVAL_134) begin
      if (_EVAL_49) begin
        if (_EVAL_36) begin
          _EVAL_182 <= _EVAL_174;
        end else begin
          _EVAL_182 <= 4'h0;
        end
      end else begin
        _EVAL_182 <= _EVAL_89;
      end
    end
    if (_EVAL_12) begin
      _EVAL_207 <= 32'h0;
    end else if (_EVAL_158) begin
      _EVAL_207 <= 32'h0;
    end else begin
      _EVAL_207 <= _EVAL_178;
    end
    if (_EVAL_86) begin
      _EVAL_240 <= _EVAL;
    end
    if (_EVAL_12) begin
      _EVAL_273 <= 4'h0;
    end else if (_EVAL_168) begin
      if (_EVAL_296) begin
        if (_EVAL_112) begin
          _EVAL_273 <= _EVAL_140;
        end else begin
          _EVAL_273 <= 4'h0;
        end
      end else begin
        _EVAL_273 <= _EVAL_91;
      end
    end
    if (_EVAL_260) begin
      _EVAL_287 <= _EVAL_16;
    end
    if (_EVAL_260) begin
      _EVAL_313 <= _EVAL_3;
    end
    if (_EVAL_86) begin
      _EVAL_315 <= _EVAL_4;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b96985ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(932e0574)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b918715)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76761e3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87943758)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_306) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2ebcf9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a3196c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(339a0b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf47f60d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8876fe4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_306) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(387e39fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33b1587c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a0fabe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a4b1252)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(283d4a21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c95ba5e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_306) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8db48486)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae5c180b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_300) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acc597a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a32219b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_306) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae7c013f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da392600)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_306) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(608f2c55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_306) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_306) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c4959c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(492119b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_306) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9ab57b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f091d851)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d542fb9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dae1136f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_300) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a29d4ce1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec65e88e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69bcbe7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_283) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2702538)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f61f5aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_300) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_300) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51928819)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc7677f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3aba11ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9be0c70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bcdd5fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c053818b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6bf0ceb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_306) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_306) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3a239b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e52752b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_306) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c56c2872)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_306) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f2010fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f173add4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59716615)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4abe0253)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bece0222)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(746026c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e6f3ff2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10fce9fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f27e1504)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_300) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad16e840)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2f6d158)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a4edd31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_300) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf511015)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bdf0204)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_300) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c20a5f21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bcab4512)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_306) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51db4b80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_283) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7b259fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7175abf1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a5e9938)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43d61f5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e2e396d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f32d61f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_306) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95ad4e95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_306) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_306) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2b3710d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_137 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46483f3c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c0db303)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfca4f1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a9359e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7566a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc85310e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_300) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1db6bb16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82be8983)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bcdd5fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e92f7a81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1135de04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(426cd13f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a67e3655)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5110ad38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc9cd39a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_308 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33b3e95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd68ba4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9cf59b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5802543)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49dc2fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d7f5992)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e90fcd0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f13c114b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9dd4f98a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18ee29eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_299) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5502c6ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_299) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3527e74d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_23 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_41 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_57 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_62 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_69 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_78 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_116 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_120 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_165 = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_167 = _RAND_9[17:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_182 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_207 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_240 = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_273 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_287 = _RAND_14[29:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_313 = _RAND_15[4:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_315 = _RAND_16[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
