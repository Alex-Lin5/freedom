//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL(
  output  _EVAL,
  input   _EVAL_0,
  output  _EVAL_1,
  input   _EVAL_2,
  output  _EVAL_3,
  output  _EVAL_4,
  output  _EVAL_5,
  output  _EVAL_6,
  input   _EVAL_7,
  input   _EVAL_8,
  output  _EVAL_9,
  output  _EVAL_10,
  input   _EVAL_11,
  input   _EVAL_12,
  output  _EVAL_13,
  input   _EVAL_14,
  input   _EVAL_15,
  input   _EVAL_16,
  output  _EVAL_17,
  input   _EVAL_18,
  input   _EVAL_19,
  input   _EVAL_20,
  input   _EVAL_21,
  input   _EVAL_22,
  input   _EVAL_23,
  output  _EVAL_24,
  output  _EVAL_25,
  input   _EVAL_26,
  output  _EVAL_27,
  input   _EVAL_28,
  output  _EVAL_29,
  input   _EVAL_30,
  output  _EVAL_31,
  input   _EVAL_32,
  input   _EVAL_33,
  input   _EVAL_34,
  output  _EVAL_35,
  output  _EVAL_36,
  input   _EVAL_37,
  input   _EVAL_38,
  input   _EVAL_39,
  input   _EVAL_40,
  input   _EVAL_41,
  input   _EVAL_42,
  output  _EVAL_43,
  output  _EVAL_44,
  input   _EVAL_45,
  output  _EVAL_46,
  output  _EVAL_47,
  output  _EVAL_48,
  output  _EVAL_49,
  input   _EVAL_50,
  input   _EVAL_51,
  output  _EVAL_52,
  output  _EVAL_53,
  input   _EVAL_54,
  output  _EVAL_55,
  input   _EVAL_56,
  output  _EVAL_57,
  input   _EVAL_58,
  input   _EVAL_59,
  output  _EVAL_60,
  input   _EVAL_61,
  output  _EVAL_62,
  input   _EVAL_63,
  input   _EVAL_64,
  output  _EVAL_65,
  input   _EVAL_66,
  input   _EVAL_67,
  output  _EVAL_68,
  input   _EVAL_69,
  output  _EVAL_70,
  output  _EVAL_71,
  input   _EVAL_72,
  output  _EVAL_73,
  output  _EVAL_74,
  input   _EVAL_75,
  output  _EVAL_76,
  input   _EVAL_77,
  output  _EVAL_78,
  input   _EVAL_79,
  output  _EVAL_80,
  input   _EVAL_81,
  output  _EVAL_82,
  output  _EVAL_83,
  output  _EVAL_84,
  output  _EVAL_85,
  input   _EVAL_86,
  input   _EVAL_87,
  input   _EVAL_88,
  input   _EVAL_89,
  input   _EVAL_90,
  output  _EVAL_91,
  input   _EVAL_92,
  input   _EVAL_93,
  input   _EVAL_94,
  input   _EVAL_95,
  output  _EVAL_96,
  output  _EVAL_97,
  input   _EVAL_98,
  input   _EVAL_99,
  input   _EVAL_100,
  output  _EVAL_101,
  input   _EVAL_102,
  input   _EVAL_103,
  input   _EVAL_104,
  output  _EVAL_105,
  input   _EVAL_106,
  input   _EVAL_107,
  output  _EVAL_108,
  output  _EVAL_109,
  output  _EVAL_110,
  input   _EVAL_111,
  output  _EVAL_112,
  input   _EVAL_113,
  input   _EVAL_114,
  output  _EVAL_115,
  input   _EVAL_116,
  output  _EVAL_117,
  input   _EVAL_118,
  input   _EVAL_119,
  input   _EVAL_120,
  input   _EVAL_121,
  output  _EVAL_122,
  input   _EVAL_123,
  output  _EVAL_124,
  output  _EVAL_125,
  input   _EVAL_126,
  input   _EVAL_127,
  output  _EVAL_128,
  input   _EVAL_129,
  input   _EVAL_130,
  input   _EVAL_131,
  output  _EVAL_132,
  output  _EVAL_133,
  output  _EVAL_134,
  output  _EVAL_135,
  output  _EVAL_136,
  input   _EVAL_137,
  output  _EVAL_138,
  output  _EVAL_139,
  input   _EVAL_140,
  output  _EVAL_141,
  input   _EVAL_142,
  output  _EVAL_143,
  input   _EVAL_144,
  output  _EVAL_145,
  input   _EVAL_146,
  output  _EVAL_147,
  output  _EVAL_148,
  input   _EVAL_149,
  output  _EVAL_150,
  output  _EVAL_151,
  input   _EVAL_152,
  input   _EVAL_153,
  input   _EVAL_154,
  input   _EVAL_155,
  output  _EVAL_156,
  input   _EVAL_157,
  input   _EVAL_158,
  output  _EVAL_159,
  input   _EVAL_160,
  input   _EVAL_161,
  output  _EVAL_162,
  input   _EVAL_163,
  input   _EVAL_164,
  output  _EVAL_165,
  output  _EVAL_166,
  output  _EVAL_167,
  output  _EVAL_168,
  output  _EVAL_169,
  input   _EVAL_170,
  output  _EVAL_171,
  output  _EVAL_172,
  output  _EVAL_173,
  input   _EVAL_174,
  input   _EVAL_175,
  output  _EVAL_176,
  output  _EVAL_177,
  output  _EVAL_178,
  output  _EVAL_179,
  input   _EVAL_180,
  output  _EVAL_181,
  input   _EVAL_182,
  output  _EVAL_183,
  output  _EVAL_184,
  input   _EVAL_185,
  input   _EVAL_186,
  input   _EVAL_187,
  output  _EVAL_188,
  output  _EVAL_189,
  input   _EVAL_190,
  input   _EVAL_191,
  output  _EVAL_192,
  output  _EVAL_193,
  output  _EVAL_194,
  output  _EVAL_195,
  input   _EVAL_196,
  input   _EVAL_197,
  input   _EVAL_198,
  input   _EVAL_199,
  input   _EVAL_200,
  input   _EVAL_201,
  input   _EVAL_202,
  output  _EVAL_203,
  output  _EVAL_204,
  output  _EVAL_205,
  output  _EVAL_206,
  output  _EVAL_207,
  output  _EVAL_208,
  input   _EVAL_209,
  input   _EVAL_210,
  input   _EVAL_211,
  output  _EVAL_212,
  input   _EVAL_213,
  output  _EVAL_214,
  output  _EVAL_215,
  output  _EVAL_216,
  output  _EVAL_217,
  output  _EVAL_218,
  output  _EVAL_219,
  output  _EVAL_220,
  output  _EVAL_221,
  input   _EVAL_222,
  input   _EVAL_223,
  output  _EVAL_224,
  input   _EVAL_225,
  output  _EVAL_226,
  input   _EVAL_227,
  output  _EVAL_228,
  output  _EVAL_229,
  input   _EVAL_230,
  input   _EVAL_231,
  input   _EVAL_232,
  input   _EVAL_233,
  input   _EVAL_234,
  output  _EVAL_235,
  output  _EVAL_236,
  output  _EVAL_237,
  input   _EVAL_238,
  output  _EVAL_239,
  output  _EVAL_240,
  input   _EVAL_241,
  output  _EVAL_242,
  output  _EVAL_243,
  output  _EVAL_244,
  output  _EVAL_245,
  output  _EVAL_246,
  input   _EVAL_247,
  output  _EVAL_248,
  input   _EVAL_249,
  input   _EVAL_250,
  output  _EVAL_251,
  output  _EVAL_252
);
  assign _EVAL_78 = _EVAL_99;
  assign _EVAL_229 = _EVAL_92;
  assign _EVAL_193 = _EVAL_241;
  assign _EVAL_35 = _EVAL_164;
  assign _EVAL_6 = _EVAL_186;
  assign _EVAL_228 = _EVAL_93;
  assign _EVAL_145 = _EVAL_187;
  assign _EVAL_134 = _EVAL_81;
  assign _EVAL_83 = _EVAL_22;
  assign _EVAL_147 = _EVAL_11;
  assign _EVAL_46 = _EVAL_90;
  assign _EVAL_181 = _EVAL_249;
  assign _EVAL_226 = _EVAL_26;
  assign _EVAL = _EVAL_21;
  assign _EVAL_125 = _EVAL_232;
  assign _EVAL_60 = _EVAL_58;
  assign _EVAL_151 = _EVAL_16;
  assign _EVAL_189 = _EVAL_12;
  assign _EVAL_165 = _EVAL_170;
  assign _EVAL_244 = _EVAL_116;
  assign _EVAL_239 = _EVAL_67;
  assign _EVAL_110 = _EVAL_40;
  assign _EVAL_52 = _EVAL_211;
  assign _EVAL_206 = _EVAL_102;
  assign _EVAL_9 = _EVAL_180;
  assign _EVAL_48 = _EVAL_87;
  assign _EVAL_235 = _EVAL_185;
  assign _EVAL_242 = _EVAL_30;
  assign _EVAL_70 = _EVAL_213;
  assign _EVAL_141 = _EVAL_41;
  assign _EVAL_136 = _EVAL_155;
  assign _EVAL_49 = _EVAL_157;
  assign _EVAL_246 = _EVAL_196;
  assign _EVAL_240 = _EVAL_39;
  assign _EVAL_214 = _EVAL_15;
  assign _EVAL_251 = _EVAL_174;
  assign _EVAL_143 = _EVAL_161;
  assign _EVAL_245 = _EVAL_182;
  assign _EVAL_177 = _EVAL_202;
  assign _EVAL_171 = _EVAL_51;
  assign _EVAL_101 = _EVAL_121;
  assign _EVAL_117 = _EVAL_7;
  assign _EVAL_80 = _EVAL_32;
  assign _EVAL_148 = _EVAL_19;
  assign _EVAL_195 = _EVAL_66;
  assign _EVAL_248 = _EVAL_198;
  assign _EVAL_24 = _EVAL_88;
  assign _EVAL_82 = _EVAL_230;
  assign _EVAL_184 = _EVAL_146;
  assign _EVAL_85 = _EVAL_222;
  assign _EVAL_236 = _EVAL_111;
  assign _EVAL_139 = _EVAL_140;
  assign _EVAL_133 = _EVAL_104;
  assign _EVAL_188 = _EVAL_200;
  assign _EVAL_179 = _EVAL_158;
  assign _EVAL_1 = _EVAL_69;
  assign _EVAL_57 = _EVAL_144;
  assign _EVAL_183 = _EVAL_233;
  assign _EVAL_252 = _EVAL_154;
  assign _EVAL_224 = _EVAL_152;
  assign _EVAL_17 = _EVAL_103;
  assign _EVAL_47 = _EVAL_119;
  assign _EVAL_65 = _EVAL_95;
  assign _EVAL_221 = _EVAL_98;
  assign _EVAL_216 = _EVAL_37;
  assign _EVAL_162 = _EVAL_64;
  assign _EVAL_44 = _EVAL_130;
  assign _EVAL_91 = _EVAL_126;
  assign _EVAL_115 = _EVAL_38;
  assign _EVAL_169 = _EVAL_153;
  assign _EVAL_53 = _EVAL_8;
  assign _EVAL_220 = _EVAL_137;
  assign _EVAL_159 = _EVAL_100;
  assign _EVAL_218 = _EVAL_54;
  assign _EVAL_62 = _EVAL_238;
  assign _EVAL_76 = _EVAL_209;
  assign _EVAL_124 = _EVAL_160;
  assign _EVAL_178 = _EVAL_107;
  assign _EVAL_29 = _EVAL_34;
  assign _EVAL_43 = _EVAL_163;
  assign _EVAL_10 = _EVAL_61;
  assign _EVAL_132 = _EVAL_142;
  assign _EVAL_27 = _EVAL_231;
  assign _EVAL_173 = _EVAL_18;
  assign _EVAL_68 = _EVAL_247;
  assign _EVAL_55 = _EVAL_113;
  assign _EVAL_109 = _EVAL_50;
  assign _EVAL_150 = _EVAL_28;
  assign _EVAL_13 = _EVAL_72;
  assign _EVAL_217 = _EVAL_190;
  assign _EVAL_219 = _EVAL_197;
  assign _EVAL_36 = _EVAL_201;
  assign _EVAL_176 = _EVAL_23;
  assign _EVAL_73 = _EVAL_123;
  assign _EVAL_156 = _EVAL_118;
  assign _EVAL_167 = _EVAL_234;
  assign _EVAL_172 = _EVAL_20;
  assign _EVAL_84 = _EVAL_191;
  assign _EVAL_4 = _EVAL_59;
  assign _EVAL_207 = _EVAL_120;
  assign _EVAL_212 = _EVAL_94;
  assign _EVAL_128 = _EVAL_225;
  assign _EVAL_31 = _EVAL_0;
  assign _EVAL_96 = _EVAL_63;
  assign _EVAL_105 = _EVAL_106;
  assign _EVAL_166 = _EVAL_56;
  assign _EVAL_194 = _EVAL_131;
  assign _EVAL_138 = _EVAL_42;
  assign _EVAL_208 = _EVAL_129;
  assign _EVAL_74 = _EVAL_45;
  assign _EVAL_203 = _EVAL_86;
  assign _EVAL_205 = _EVAL_114;
  assign _EVAL_5 = _EVAL_127;
  assign _EVAL_112 = _EVAL_79;
  assign _EVAL_97 = _EVAL_2;
  assign _EVAL_215 = _EVAL_14;
  assign _EVAL_204 = _EVAL_89;
  assign _EVAL_122 = _EVAL_33;
  assign _EVAL_237 = _EVAL_223;
  assign _EVAL_168 = _EVAL_75;
  assign _EVAL_135 = _EVAL_77;
  assign _EVAL_71 = _EVAL_250;
  assign _EVAL_3 = _EVAL_149;
  assign _EVAL_243 = _EVAL_175;
  assign _EVAL_25 = _EVAL_199;
  assign _EVAL_192 = _EVAL_210;
  assign _EVAL_108 = _EVAL_227;
endmodule
