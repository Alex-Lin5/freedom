//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_77(
  input  [31:0] _EVAL,
  output [2:0]  _EVAL_0,
  output [1:0]  _EVAL_1,
  input         _EVAL_2,
  input  [4:0]  _EVAL_3,
  input  [31:0] _EVAL_4,
  input  [2:0]  _EVAL_5,
  output [2:0]  _EVAL_6,
  output [4:0]  _EVAL_7,
  output [2:0]  _EVAL_8,
  input         _EVAL_9,
  output [4:0]  _EVAL_10,
  output [3:0]  _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [4:0]  _EVAL_13,
  output [1:0]  _EVAL_14,
  output        _EVAL_15,
  output        _EVAL_16,
  output        _EVAL_17,
  input  [2:0]  _EVAL_18,
  input  [4:0]  _EVAL_19,
  input  [31:0] _EVAL_20,
  input         _EVAL_21,
  output [3:0]  _EVAL_22,
  input  [31:0] _EVAL_23,
  input  [3:0]  _EVAL_24,
  output [31:0] _EVAL_25,
  input         _EVAL_26,
  output [31:0] _EVAL_27,
  output [31:0] _EVAL_28,
  output [2:0]  _EVAL_29,
  output [2:0]  _EVAL_30,
  input         _EVAL_31,
  output [31:0] _EVAL_32,
  input  [2:0]  _EVAL_33,
  input  [1:0]  _EVAL_34,
  input         _EVAL_35,
  output [2:0]  _EVAL_36,
  output [31:0] _EVAL_37,
  input  [2:0]  _EVAL_38,
  output [2:0]  _EVAL_39,
  output [2:0]  _EVAL_40,
  input  [1:0]  _EVAL_41,
  output        _EVAL_42,
  input  [2:0]  _EVAL_43,
  output [4:0]  _EVAL_44,
  input  [2:0]  _EVAL_45
);
  wire  _EVAL_46;
  wire  rsource__EVAL;
  wire  rsource__EVAL_0;
  wire [4:0] rsource__EVAL_1;
  wire [2:0] rsource__EVAL_2;
  wire [4:0] rsource__EVAL_3;
  wire [2:0] rsource__EVAL_4;
  wire [2:0] rsource__EVAL_5;
  wire [3:0] rsource__EVAL_6;
  wire [2:0] rsource__EVAL_7;
  wire [4:0] rsource__EVAL_8;
  wire [2:0] rsource__EVAL_9;
  wire [2:0] rsource__EVAL_10;
  wire [1:0] rsource__EVAL_11;
  wire [2:0] rsource__EVAL_12;
  wire [3:0] rsource__EVAL_13;
  wire [31:0] rsource__EVAL_14;
  wire [2:0] rsource__EVAL_15;
  wire  rsource__EVAL_16;
  wire  rsource__EVAL_17;
  wire [31:0] rsource__EVAL_18;
  wire  rsource__EVAL_19;
  wire [31:0] rsource__EVAL_20;
  wire [4:0] rsource__EVAL_21;
  wire [31:0] rsource__EVAL_22;
  wire [31:0] rsource__EVAL_23;
  wire [4:0] rsource__EVAL_24;
  wire  rsource__EVAL_25;
  wire [31:0] rsource__EVAL_26;
  wire [1:0] rsource__EVAL_27;
  wire [31:0] rsource__EVAL_28;
  wire [31:0] rsource__EVAL_29;
  wire [2:0] rsource__EVAL_30;
  wire [2:0] rsource__EVAL_31;
  wire  rsource__EVAL_32;
  wire [2:0] rsource__EVAL_33;
  wire  rsource__EVAL_34;
  wire [2:0] rsource__EVAL_35;
  wire [1:0] rsource__EVAL_36;
  wire [2:0] rsource__EVAL_37;
  wire [4:0] rsource__EVAL_38;
  wire [1:0] rsource__EVAL_39;
  wire [2:0] rsource__EVAL_40;
  wire [31:0] rsource__EVAL_41;
  wire [2:0] rsource__EVAL_42;
  wire  rsource__EVAL_43;
  wire  rsource__EVAL_44;
  wire [3:0] rsource__EVAL_45;
  wire [31:0] _EVAL_47;
  wire [2:0] _EVAL_48;
  wire [2:0] _EVAL_49;
  wire [4:0] _EVAL_50;
  wire  _EVAL_51;
  wire [31:0] _EVAL_52;
  wire [2:0] _EVAL_53;
  wire [31:0] _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire [2:0] _EVAL_57;
  wire [4:0] _EVAL_58;
  wire [2:0] _EVAL_59;
  wire [31:0] _EVAL_60;
  wire  _EVAL_61;
  wire [3:0] _EVAL_62;
  wire  _EVAL_63;
  wire [2:0] _EVAL_64;
  wire [3:0] _EVAL_65;
  wire  _EVAL_66;
  wire [2:0] _EVAL_67;
  wire [2:0] _EVAL_68;
  wire [31:0] _EVAL_69;
  wire [4:0] _EVAL_70;
  wire [2:0] _EVAL_71;
  wire [31:0] _EVAL_72;
  wire [2:0] _EVAL_73;
  wire [4:0] _EVAL_74;
  wire  _EVAL_75;
  _EVAL_76 rsource (
    ._EVAL(rsource__EVAL),
    ._EVAL_0(rsource__EVAL_0),
    ._EVAL_1(rsource__EVAL_1),
    ._EVAL_2(rsource__EVAL_2),
    ._EVAL_3(rsource__EVAL_3),
    ._EVAL_4(rsource__EVAL_4),
    ._EVAL_5(rsource__EVAL_5),
    ._EVAL_6(rsource__EVAL_6),
    ._EVAL_7(rsource__EVAL_7),
    ._EVAL_8(rsource__EVAL_8),
    ._EVAL_9(rsource__EVAL_9),
    ._EVAL_10(rsource__EVAL_10),
    ._EVAL_11(rsource__EVAL_11),
    ._EVAL_12(rsource__EVAL_12),
    ._EVAL_13(rsource__EVAL_13),
    ._EVAL_14(rsource__EVAL_14),
    ._EVAL_15(rsource__EVAL_15),
    ._EVAL_16(rsource__EVAL_16),
    ._EVAL_17(rsource__EVAL_17),
    ._EVAL_18(rsource__EVAL_18),
    ._EVAL_19(rsource__EVAL_19),
    ._EVAL_20(rsource__EVAL_20),
    ._EVAL_21(rsource__EVAL_21),
    ._EVAL_22(rsource__EVAL_22),
    ._EVAL_23(rsource__EVAL_23),
    ._EVAL_24(rsource__EVAL_24),
    ._EVAL_25(rsource__EVAL_25),
    ._EVAL_26(rsource__EVAL_26),
    ._EVAL_27(rsource__EVAL_27),
    ._EVAL_28(rsource__EVAL_28),
    ._EVAL_29(rsource__EVAL_29),
    ._EVAL_30(rsource__EVAL_30),
    ._EVAL_31(rsource__EVAL_31),
    ._EVAL_32(rsource__EVAL_32),
    ._EVAL_33(rsource__EVAL_33),
    ._EVAL_34(rsource__EVAL_34),
    ._EVAL_35(rsource__EVAL_35),
    ._EVAL_36(rsource__EVAL_36),
    ._EVAL_37(rsource__EVAL_37),
    ._EVAL_38(rsource__EVAL_38),
    ._EVAL_39(rsource__EVAL_39),
    ._EVAL_40(rsource__EVAL_40),
    ._EVAL_41(rsource__EVAL_41),
    ._EVAL_42(rsource__EVAL_42),
    ._EVAL_43(rsource__EVAL_43),
    ._EVAL_44(rsource__EVAL_44),
    ._EVAL_45(rsource__EVAL_45)
  );
  assign _EVAL_62 = _EVAL_24;
  assign rsource__EVAL_18 = _EVAL_52;
  assign rsource__EVAL_8 = _EVAL_3;
  assign _EVAL_28 = _EVAL_60;
  assign _EVAL_75 = _EVAL_66;
  assign _EVAL_16 = _EVAL_75;
  assign _EVAL_64 = _EVAL_38;
  assign _EVAL_27 = rsource__EVAL_26;
  assign _EVAL_57 = _EVAL_18;
  assign _EVAL_25 = rsource__EVAL_29;
  assign rsource__EVAL_0 = _EVAL_26;
  assign _EVAL_17 = _EVAL_55;
  assign rsource__EVAL_13 = _EVAL_65;
  assign _EVAL_36 = _EVAL_68;
  assign _EVAL_48 = _EVAL_57;
  assign _EVAL_46 = _EVAL_9;
  assign _EVAL_70 = _EVAL_74;
  assign rsource__EVAL_34 = _EVAL_2;
  assign _EVAL_67 = _EVAL_59;
  assign _EVAL_56 = rsource__EVAL_17;
  assign _EVAL_14 = rsource__EVAL_27;
  assign rsource__EVAL_39 = _EVAL_41;
  assign _EVAL_51 = _EVAL_46;
  assign _EVAL_59 = _EVAL_33;
  assign rsource__EVAL_14 = _EVAL;
  assign _EVAL_30 = rsource__EVAL_12;
  assign _EVAL_11 = rsource__EVAL_45;
  assign _EVAL_7 = rsource__EVAL_21;
  assign _EVAL_55 = _EVAL_56;
  assign _EVAL_0 = rsource__EVAL_42;
  assign rsource__EVAL_36 = _EVAL_34;
  assign rsource__EVAL_35 = _EVAL_48;
  assign _EVAL_15 = rsource__EVAL_44;
  assign _EVAL_52 = _EVAL_72;
  assign _EVAL_72 = _EVAL_20;
  assign rsource__EVAL_40 = _EVAL_12;
  assign _EVAL_50 = _EVAL_13;
  assign rsource__EVAL_43 = _EVAL_21;
  assign _EVAL_32 = rsource__EVAL_23;
  assign _EVAL_44 = rsource__EVAL_24;
  assign _EVAL_58 = _EVAL_50;
  assign _EVAL_40 = rsource__EVAL_10;
  assign rsource__EVAL_19 = _EVAL_51;
  assign rsource__EVAL_30 = _EVAL_45;
  assign _EVAL_74 = rsource__EVAL_1;
  assign rsource__EVAL_9 = _EVAL_53;
  assign _EVAL_53 = _EVAL_64;
  assign _EVAL_37 = rsource__EVAL_28;
  assign rsource__EVAL_16 = _EVAL_61;
  assign _EVAL_65 = _EVAL_62;
  assign _EVAL_47 = rsource__EVAL_41;
  assign _EVAL_8 = rsource__EVAL_37;
  assign rsource__EVAL_38 = _EVAL_58;
  assign _EVAL_6 = _EVAL_71;
  assign _EVAL_39 = rsource__EVAL_31;
  assign _EVAL_1 = rsource__EVAL_11;
  assign _EVAL_42 = rsource__EVAL_25;
  assign _EVAL_54 = _EVAL_23;
  assign _EVAL_10 = _EVAL_70;
  assign _EVAL_69 = _EVAL_54;
  assign rsource__EVAL_20 = _EVAL_4;
  assign _EVAL_66 = rsource__EVAL_32;
  assign _EVAL_63 = _EVAL_31;
  assign rsource__EVAL_15 = _EVAL_67;
  assign _EVAL_29 = rsource__EVAL_4;
  assign _EVAL_73 = rsource__EVAL_5;
  assign _EVAL_68 = _EVAL_49;
  assign _EVAL_60 = _EVAL_47;
  assign rsource__EVAL = _EVAL_35;
  assign rsource__EVAL_2 = _EVAL_5;
  assign _EVAL_61 = _EVAL_63;
  assign _EVAL_49 = rsource__EVAL_33;
  assign _EVAL_22 = rsource__EVAL_6;
  assign rsource__EVAL_3 = _EVAL_19;
  assign rsource__EVAL_22 = _EVAL_69;
  assign rsource__EVAL_7 = _EVAL_43;
  assign _EVAL_71 = _EVAL_73;
endmodule
