//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_134(
  output        _EVAL,
  output        _EVAL_0,
  input  [31:0] _EVAL_1,
  input  [31:0] _EVAL_2,
  output        _EVAL_3,
  output        _EVAL_4,
  input         _EVAL_5,
  output        _EVAL_6,
  input         _EVAL_7,
  input  [3:0]  _EVAL_8,
  input         _EVAL_9,
  output [3:0]  _EVAL_10,
  output [31:0] _EVAL_11,
  output        _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  output        _EVAL_16,
  input         _EVAL_17,
  output        _EVAL_18,
  input         _EVAL_19,
  input  [2:0]  _EVAL_20,
  input         _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23,
  output        _EVAL_24,
  input         _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  input  [31:0] _EVAL_30,
  input  [2:0]  _EVAL_31,
  input         _EVAL_32,
  input         _EVAL_33,
  input  [31:0] _EVAL_34,
  output [2:0]  _EVAL_35,
  input         _EVAL_36,
  input         _EVAL_37,
  output [2:0]  _EVAL_38,
  output [4:0]  _EVAL_39,
  input         _EVAL_40,
  input         _EVAL_41,
  input         _EVAL_42,
  input         _EVAL_43,
  output [3:0]  _EVAL_44,
  output [31:0] _EVAL_45,
  output [31:0] _EVAL_46,
  output [2:0]  _EVAL_47,
  output [3:0]  _EVAL_48,
  input         _EVAL_49,
  input         _EVAL_50,
  input  [3:0]  _EVAL_51,
  output        _EVAL_52,
  input  [1:0]  _EVAL_53,
  input         _EVAL_54,
  output        _EVAL_55,
  input  [31:0] _EVAL_56,
  input         _EVAL_57,
  input  [2:0]  _EVAL_58,
  input         _EVAL_59,
  input  [2:0]  _EVAL_60,
  input  [3:0]  _EVAL_61,
  output        _EVAL_62,
  output [2:0]  _EVAL_63,
  input         _EVAL_64,
  input  [31:0] _EVAL_65,
  input  [4:0]  _EVAL_66,
  input         _EVAL_67,
  input         _EVAL_68
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] _EVAL_69;
  wire  dcache__EVAL;
  wire  dcache__EVAL_0;
  wire  dcache__EVAL_1;
  wire  dcache__EVAL_2;
  wire [31:0] dcache__EVAL_3;
  wire  dcache__EVAL_4;
  wire  dcache__EVAL_5;
  wire [3:0] dcache__EVAL_6;
  wire [1:0] dcache__EVAL_7;
  wire [29:0] dcache__EVAL_8;
  wire [31:0] dcache__EVAL_9;
  wire  dcache__EVAL_10;
  wire  dcache__EVAL_11;
  wire  dcache__EVAL_12;
  wire  dcache__EVAL_13;
  wire [1:0] dcache__EVAL_14;
  wire  dcache__EVAL_15;
  wire [31:0] dcache__EVAL_16;
  wire  dcache__EVAL_17;
  wire [2:0] dcache__EVAL_18;
  wire  dcache__EVAL_19;
  wire  dcache__EVAL_20;
  wire [1:0] dcache__EVAL_21;
  wire [31:0] dcache__EVAL_22;
  wire  dcache__EVAL_23;
  wire [6:0] dcache__EVAL_24;
  wire  dcache__EVAL_25;
  wire  dcache__EVAL_26;
  wire  dcache__EVAL_27;
  wire  dcache__EVAL_28;
  wire  dcache__EVAL_29;
  wire  dcache__EVAL_30;
  wire  dcache__EVAL_31;
  wire  dcache__EVAL_32;
  wire  dcache__EVAL_33;
  wire  dcache__EVAL_34;
  wire [2:0] dcache__EVAL_35;
  wire  dcache__EVAL_36;
  wire [29:0] dcache__EVAL_37;
  wire [31:0] dcache__EVAL_38;
  wire [31:0] dcache__EVAL_39;
  wire  dcache__EVAL_40;
  wire  dcache__EVAL_41;
  wire [31:0] dcache__EVAL_42;
  wire  dcache__EVAL_43;
  wire  dcache__EVAL_44;
  wire  dcache__EVAL_45;
  wire  dcache__EVAL_46;
  wire  dcache__EVAL_47;
  wire  dcache__EVAL_48;
  wire  dcache__EVAL_49;
  wire  dcache__EVAL_50;
  wire [2:0] dcache__EVAL_51;
  wire [31:0] dcache__EVAL_52;
  wire  dcache__EVAL_53;
  wire [31:0] dcache__EVAL_54;
  wire [1:0] dcache__EVAL_55;
  wire  dcache__EVAL_56;
  wire [31:0] dcache__EVAL_57;
  wire [31:0] dcache__EVAL_58;
  wire [29:0] dcache__EVAL_59;
  wire [1:0] dcache__EVAL_60;
  wire [29:0] dcache__EVAL_61;
  wire  dcache__EVAL_62;
  wire  dcache__EVAL_63;
  wire [3:0] dcache__EVAL_64;
  wire [1:0] dcache__EVAL_65;
  wire [1:0] dcache__EVAL_66;
  wire [1:0] dcache__EVAL_67;
  wire  dcache__EVAL_68;
  wire  dcache__EVAL_69;
  wire  dcache__EVAL_70;
  wire [29:0] dcache__EVAL_71;
  wire  dcache__EVAL_72;
  wire  dcache__EVAL_73;
  wire  dcache__EVAL_74;
  wire  dcache__EVAL_75;
  wire [31:0] dcache__EVAL_76;
  wire [6:0] dcache__EVAL_77;
  wire [29:0] dcache__EVAL_78;
  wire [3:0] dcache__EVAL_79;
  wire  dcache__EVAL_80;
  wire [29:0] dcache__EVAL_81;
  wire [1:0] dcache__EVAL_82;
  wire  dcache__EVAL_83;
  wire  dcache__EVAL_84;
  wire [31:0] dcache__EVAL_85;
  wire  dcache__EVAL_86;
  wire [3:0] dcache__EVAL_87;
  wire  dcache__EVAL_88;
  wire [1:0] dcache__EVAL_89;
  wire [31:0] dcache__EVAL_90;
  wire [29:0] dcache__EVAL_91;
  wire [31:0] dcache__EVAL_92;
  wire  dcache__EVAL_93;
  wire  dcache__EVAL_94;
  wire [3:0] dcache__EVAL_95;
  wire [1:0] dcache__EVAL_96;
  wire  dcache__EVAL_97;
  wire [4:0] dcache__EVAL_98;
  wire  dcache__EVAL_99;
  wire [31:0] dcache__EVAL_100;
  wire  dcache__EVAL_101;
  wire  dcache__EVAL_102;
  wire  dcache__EVAL_103;
  wire  dcache__EVAL_104;
  wire  dcache__EVAL_105;
  wire [2:0] dcache__EVAL_106;
  wire [1:0] dcache__EVAL_107;
  wire  dcache__EVAL_108;
  wire  dcache__EVAL_109;
  wire  dcache__EVAL_110;
  wire [1:0] dcache__EVAL_111;
  wire  dcache__EVAL_112;
  wire  dcache__EVAL_113;
  wire [31:0] dcache__EVAL_114;
  wire [3:0] dcache__EVAL_115;
  wire  dcache__EVAL_116;
  wire  dcache__EVAL_117;
  wire  dcache__EVAL_118;
  wire [31:0] dcache__EVAL_119;
  wire  dcache__EVAL_120;
  wire  dcache__EVAL_121;
  wire [1:0] dcache__EVAL_122;
  wire  dcache__EVAL_123;
  wire [4:0] dcache__EVAL_124;
  wire [31:0] dcache__EVAL_125;
  wire  dcache__EVAL_126;
  wire [2:0] dcache__EVAL_127;
  wire  dcache__EVAL_128;
  wire  _EVAL_71;
  wire [3:0] dtim_adapter__EVAL;
  wire  dtim_adapter__EVAL_0;
  wire [2:0] dtim_adapter__EVAL_1;
  wire  dtim_adapter__EVAL_2;
  wire  dtim_adapter__EVAL_3;
  wire  dtim_adapter__EVAL_4;
  wire  dtim_adapter__EVAL_5;
  wire  dtim_adapter__EVAL_6;
  wire [31:0] dtim_adapter__EVAL_7;
  wire [31:0] dtim_adapter__EVAL_8;
  wire  dtim_adapter__EVAL_9;
  wire [31:0] dtim_adapter__EVAL_10;
  wire [3:0] dtim_adapter__EVAL_11;
  wire [1:0] dtim_adapter__EVAL_12;
  wire  dtim_adapter__EVAL_13;
  wire [1:0] dtim_adapter__EVAL_14;
  wire [10:0] dtim_adapter__EVAL_15;
  wire  dtim_adapter__EVAL_16;
  wire [1:0] dtim_adapter__EVAL_17;
  wire  dtim_adapter__EVAL_18;
  wire  dtim_adapter__EVAL_19;
  wire [31:0] dtim_adapter__EVAL_20;
  wire [2:0] dtim_adapter__EVAL_21;
  wire [10:0] dtim_adapter__EVAL_22;
  wire [31:0] dtim_adapter__EVAL_23;
  wire [2:0] dtim_adapter__EVAL_24;
  wire [4:0] dtim_adapter__EVAL_25;
  wire [31:0] dtim_adapter__EVAL_26;
  wire [2:0] tlMasterXbar__EVAL;
  wire [2:0] tlMasterXbar__EVAL_0;
  wire  tlMasterXbar__EVAL_1;
  wire [3:0] tlMasterXbar__EVAL_2;
  wire  tlMasterXbar__EVAL_3;
  wire [31:0] tlMasterXbar__EVAL_4;
  wire [3:0] tlMasterXbar__EVAL_5;
  wire [2:0] tlMasterXbar__EVAL_6;
  wire [3:0] tlMasterXbar__EVAL_7;
  wire  tlMasterXbar__EVAL_8;
  wire  tlMasterXbar__EVAL_9;
  wire [3:0] tlMasterXbar__EVAL_10;
  wire  tlMasterXbar__EVAL_11;
  wire [3:0] tlMasterXbar__EVAL_12;
  wire  tlMasterXbar__EVAL_13;
  wire  tlMasterXbar__EVAL_14;
  wire  tlMasterXbar__EVAL_15;
  wire  tlMasterXbar__EVAL_16;
  wire [2:0] tlMasterXbar__EVAL_17;
  wire  tlMasterXbar__EVAL_18;
  wire [3:0] tlMasterXbar__EVAL_19;
  wire  tlMasterXbar__EVAL_20;
  wire  tlMasterXbar__EVAL_21;
  wire [3:0] tlMasterXbar__EVAL_22;
  wire [31:0] tlMasterXbar__EVAL_23;
  wire [31:0] tlMasterXbar__EVAL_24;
  wire  tlMasterXbar__EVAL_25;
  wire [1:0] tlMasterXbar__EVAL_26;
  wire [2:0] tlMasterXbar__EVAL_27;
  wire  tlMasterXbar__EVAL_28;
  wire  tlMasterXbar__EVAL_29;
  wire  tlMasterXbar__EVAL_30;
  wire  tlMasterXbar__EVAL_31;
  wire [31:0] tlMasterXbar__EVAL_32;
  wire  tlMasterXbar__EVAL_33;
  wire  tlMasterXbar__EVAL_34;
  wire [2:0] tlMasterXbar__EVAL_35;
  wire  tlMasterXbar__EVAL_36;
  wire [31:0] tlMasterXbar__EVAL_37;
  wire  tlMasterXbar__EVAL_38;
  wire  tlMasterXbar__EVAL_39;
  wire  tlMasterXbar__EVAL_40;
  wire [3:0] tlMasterXbar__EVAL_41;
  wire  tlMasterXbar__EVAL_42;
  wire [3:0] tlMasterXbar__EVAL_43;
  wire  tlMasterXbar__EVAL_44;
  wire  tlMasterXbar__EVAL_45;
  wire [2:0] tlMasterXbar__EVAL_46;
  wire [2:0] tlMasterXbar__EVAL_47;
  wire [31:0] tlMasterXbar__EVAL_48;
  wire  tlMasterXbar__EVAL_49;
  wire  tlMasterXbar__EVAL_50;
  wire  tlMasterXbar__EVAL_51;
  wire [31:0] tlMasterXbar__EVAL_52;
  wire  tlMasterXbar__EVAL_53;
  wire [1:0] tlMasterXbar__EVAL_54;
  wire [2:0] tlMasterXbar__EVAL_55;
  wire [31:0] tlMasterXbar__EVAL_56;
  wire  tlMasterXbar__EVAL_57;
  wire  _EVAL_72;
  wire [31:0] fragmenter_1__EVAL;
  wire [3:0] fragmenter_1__EVAL_0;
  wire  fragmenter_1__EVAL_1;
  wire  fragmenter_1__EVAL_2;
  wire [10:0] fragmenter_1__EVAL_3;
  wire  fragmenter_1__EVAL_4;
  wire [2:0] fragmenter_1__EVAL_5;
  wire [31:0] fragmenter_1__EVAL_6;
  wire  fragmenter_1__EVAL_7;
  wire [2:0] fragmenter_1__EVAL_8;
  wire [31:0] fragmenter_1__EVAL_9;
  wire  fragmenter_1__EVAL_10;
  wire [1:0] fragmenter_1__EVAL_11;
  wire [4:0] fragmenter_1__EVAL_12;
  wire [2:0] fragmenter_1__EVAL_13;
  wire  fragmenter_1__EVAL_14;
  wire  fragmenter_1__EVAL_15;
  wire [31:0] fragmenter_1__EVAL_16;
  wire [4:0] fragmenter_1__EVAL_17;
  wire [2:0] fragmenter_1__EVAL_18;
  wire [3:0] fragmenter_1__EVAL_19;
  wire  fragmenter_1__EVAL_20;
  wire [1:0] fragmenter_1__EVAL_21;
  wire  fragmenter_1__EVAL_22;
  wire [31:0] fragmenter_1__EVAL_23;
  wire [2:0] fragmenter_1__EVAL_24;
  wire [2:0] fragmenter_1__EVAL_25;
  wire [10:0] fragmenter_1__EVAL_26;
  wire [2:0] fragmenter_1__EVAL_27;
  wire [2:0] fragmenter_1__EVAL_28;
  wire  fragmenter_1__EVAL_29;
  wire [31:0] fragmenter_1__EVAL_30;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire [29:0] ptw__EVAL;
  wire  ptw__EVAL_0;
  wire [1:0] ptw__EVAL_1;
  wire [29:0] ptw__EVAL_2;
  wire [31:0] ptw__EVAL_3;
  wire  ptw__EVAL_4;
  wire [29:0] ptw__EVAL_5;
  wire  ptw__EVAL_6;
  wire  ptw__EVAL_7;
  wire [31:0] ptw__EVAL_8;
  wire  ptw__EVAL_9;
  wire  ptw__EVAL_10;
  wire [1:0] ptw__EVAL_11;
  wire  ptw__EVAL_12;
  wire  ptw__EVAL_13;
  wire  ptw__EVAL_14;
  wire  ptw__EVAL_15;
  wire  ptw__EVAL_16;
  wire  ptw__EVAL_17;
  wire  ptw__EVAL_18;
  wire [29:0] ptw__EVAL_19;
  wire [1:0] ptw__EVAL_20;
  wire  ptw__EVAL_21;
  wire  ptw__EVAL_22;
  wire  ptw__EVAL_23;
  wire  ptw__EVAL_24;
  wire  ptw__EVAL_25;
  wire  ptw__EVAL_26;
  wire  ptw__EVAL_27;
  wire  ptw__EVAL_28;
  wire  ptw__EVAL_29;
  wire  ptw__EVAL_30;
  wire  ptw__EVAL_31;
  wire  ptw__EVAL_32;
  wire  ptw__EVAL_33;
  wire [1:0] ptw__EVAL_34;
  wire  ptw__EVAL_35;
  wire  ptw__EVAL_36;
  wire  ptw__EVAL_37;
  wire  ptw__EVAL_38;
  wire [1:0] ptw__EVAL_39;
  wire [29:0] ptw__EVAL_40;
  wire [31:0] ptw__EVAL_41;
  wire  ptw__EVAL_42;
  wire  ptw__EVAL_43;
  wire [31:0] ptw__EVAL_44;
  wire  ptw__EVAL_45;
  wire  ptw__EVAL_46;
  wire  ptw__EVAL_47;
  wire [29:0] ptw__EVAL_48;
  wire [1:0] ptw__EVAL_49;
  wire [29:0] ptw__EVAL_50;
  wire  ptw__EVAL_51;
  wire  ptw__EVAL_52;
  wire  ptw__EVAL_53;
  wire [1:0] ptw__EVAL_54;
  wire  ptw__EVAL_55;
  wire  ptw__EVAL_56;
  wire  ptw__EVAL_57;
  wire  ptw__EVAL_58;
  wire  ptw__EVAL_59;
  wire  ptw__EVAL_60;
  wire [1:0] ptw__EVAL_61;
  wire  ptw__EVAL_62;
  wire [31:0] ptw__EVAL_63;
  wire [31:0] ptw__EVAL_64;
  wire [29:0] ptw__EVAL_65;
  wire  ptw__EVAL_66;
  wire  ptw__EVAL_67;
  wire  ptw__EVAL_68;
  wire [29:0] ptw__EVAL_69;
  wire  ptw__EVAL_70;
  wire [31:0] ptw__EVAL_71;
  wire  ptw__EVAL_72;
  wire  ptw__EVAL_73;
  wire [1:0] ptw__EVAL_74;
  wire [29:0] ptw__EVAL_75;
  wire  ptw__EVAL_76;
  wire [29:0] ptw__EVAL_77;
  wire [31:0] ptw__EVAL_78;
  wire  ptw__EVAL_79;
  wire  ptw__EVAL_80;
  wire [1:0] ptw__EVAL_81;
  wire [29:0] ptw__EVAL_82;
  wire  ptw__EVAL_83;
  wire  ptw__EVAL_84;
  wire  ptw__EVAL_85;
  wire  ptw__EVAL_86;
  wire [31:0] ptw__EVAL_87;
  wire  ptw__EVAL_88;
  wire [31:0] ptw__EVAL_89;
  wire [31:0] ptw__EVAL_90;
  wire  ptw__EVAL_91;
  wire [1:0] ptw__EVAL_92;
  wire [1:0] ptw__EVAL_93;
  wire [31:0] ptw__EVAL_94;
  wire [1:0] ptw__EVAL_95;
  wire  ptw__EVAL_96;
  wire [29:0] ptw__EVAL_97;
  wire  ptw__EVAL_98;
  wire  ptw__EVAL_99;
  wire [1:0] ptw__EVAL_100;
  wire [29:0] ptw__EVAL_101;
  wire  ptw__EVAL_102;
  wire [31:0] ptw__EVAL_103;
  wire  ptw__EVAL_104;
  wire [1:0] ptw__EVAL_105;
  wire [29:0] ptw__EVAL_106;
  wire  ptw__EVAL_107;
  wire [1:0] ptw__EVAL_108;
  wire  ptw__EVAL_109;
  wire [1:0] ptw__EVAL_110;
  wire [31:0] ptw__EVAL_111;
  wire [1:0] ptw__EVAL_112;
  wire [31:0] ptw__EVAL_113;
  wire  ptw__EVAL_114;
  wire [1:0] ptw__EVAL_115;
  wire  ptw__EVAL_116;
  wire  ptw__EVAL_117;
  wire [31:0] ptw__EVAL_118;
  wire  ptw__EVAL_119;
  wire [31:0] ptw__EVAL_120;
  wire [29:0] ptw__EVAL_121;
  wire [1:0] ptw__EVAL_122;
  wire  ptw__EVAL_123;
  wire  ptw__EVAL_124;
  wire [29:0] ptw__EVAL_125;
  wire [31:0] ptw__EVAL_126;
  wire  ptw__EVAL_127;
  wire  ptw__EVAL_128;
  wire [29:0] ptw__EVAL_129;
  wire  ptw__EVAL_130;
  wire  ptw__EVAL_131;
  wire [1:0] ptw__EVAL_132;
  wire  ptw__EVAL_133;
  wire [29:0] ptw__EVAL_134;
  wire  ptw__EVAL_135;
  wire  ptw__EVAL_136;
  wire [29:0] ptw__EVAL_137;
  wire [29:0] ptw__EVAL_138;
  wire [1:0] ptw__EVAL_139;
  wire [29:0] ptw__EVAL_140;
  wire  ptw__EVAL_141;
  wire  ptw__EVAL_142;
  wire [31:0] ptw__EVAL_143;
  wire  ptw__EVAL_144;
  wire  ptw__EVAL_145;
  wire  ptw__EVAL_146;
  wire [31:0] ptw__EVAL_147;
  wire  ptw__EVAL_148;
  wire [1:0] ptw__EVAL_149;
  wire  ptw__EVAL_150;
  wire [29:0] ptw__EVAL_151;
  wire  ptw__EVAL_152;
  wire [31:0] ptw__EVAL_153;
  wire  ptw__EVAL_154;
  wire  ptw__EVAL_155;
  wire [31:0] ptw__EVAL_156;
  wire [29:0] ptw__EVAL_157;
  wire  ptw__EVAL_158;
  wire [31:0] ptw__EVAL_159;
  wire  ptw__EVAL_160;
  wire  ptw__EVAL_161;
  wire [1:0] ptw__EVAL_162;
  wire [31:0] ptw__EVAL_163;
  wire  ptw__EVAL_164;
  wire [1:0] ptw__EVAL_165;
  wire  ptw__EVAL_166;
  wire  ptw__EVAL_167;
  wire [31:0] ptw__EVAL_168;
  wire  ptw__EVAL_169;
  wire  ptw__EVAL_170;
  wire  ptw__EVAL_171;
  wire [1:0] ptw__EVAL_172;
  wire  ptw__EVAL_173;
  wire [31:0] ptw__EVAL_174;
  wire  ptw__EVAL_175;
  wire  ptw__EVAL_176;
  wire [31:0] ptw__EVAL_177;
  wire [1:0] ptw__EVAL_178;
  wire  ptw__EVAL_179;
  wire  ptw__EVAL_180;
  wire  ptw__EVAL_181;
  wire [1:0] ptw__EVAL_182;
  wire [31:0] ptw__EVAL_183;
  wire [31:0] ptw__EVAL_184;
  wire  ptw__EVAL_185;
  wire  ptw__EVAL_186;
  wire  ptw__EVAL_187;
  wire [31:0] _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_78;
  wire  dcacheArb__EVAL;
  wire  dcacheArb__EVAL_0;
  wire  dcacheArb__EVAL_1;
  wire [31:0] dcacheArb__EVAL_2;
  wire [4:0] dcacheArb__EVAL_3;
  wire [3:0] dcacheArb__EVAL_4;
  wire [31:0] dcacheArb__EVAL_5;
  wire [31:0] dcacheArb__EVAL_6;
  wire  dcacheArb__EVAL_7;
  wire  dcacheArb__EVAL_8;
  wire  dcacheArb__EVAL_9;
  wire  dcacheArb__EVAL_10;
  wire  dcacheArb__EVAL_11;
  wire  dcacheArb__EVAL_12;
  wire  dcacheArb__EVAL_13;
  wire  dcacheArb__EVAL_14;
  wire  dcacheArb__EVAL_15;
  wire [31:0] dcacheArb__EVAL_16;
  wire  dcacheArb__EVAL_17;
  wire [31:0] dcacheArb__EVAL_18;
  wire [3:0] dcacheArb__EVAL_19;
  wire  dcacheArb__EVAL_20;
  wire  dcacheArb__EVAL_21;
  wire  dcacheArb__EVAL_22;
  wire [31:0] dcacheArb__EVAL_23;
  wire  dcacheArb__EVAL_24;
  wire [6:0] dcacheArb__EVAL_25;
  wire [1:0] dcacheArb__EVAL_26;
  wire [31:0] dcacheArb__EVAL_27;
  wire [31:0] dcacheArb__EVAL_28;
  wire  dcacheArb__EVAL_29;
  wire  dcacheArb__EVAL_30;
  wire  dcacheArb__EVAL_31;
  wire [6:0] dcacheArb__EVAL_32;
  wire  dcacheArb__EVAL_33;
  wire [1:0] dcacheArb__EVAL_34;
  wire  dcacheArb__EVAL_35;
  wire [6:0] dcacheArb__EVAL_36;
  wire [4:0] dcacheArb__EVAL_37;
  wire  dcacheArb__EVAL_38;
  wire [31:0] dcacheArb__EVAL_39;
  wire  dcacheArb__EVAL_40;
  wire  dcacheArb__EVAL_41;
  wire  dcacheArb__EVAL_42;
  wire  dcacheArb__EVAL_43;
  wire [4:0] dcacheArb__EVAL_44;
  wire  dcacheArb__EVAL_45;
  wire [4:0] dcacheArb__EVAL_46;
  wire [1:0] dcacheArb__EVAL_47;
  wire [1:0] dcacheArb__EVAL_48;
  wire  dcacheArb__EVAL_49;
  wire  dcacheArb__EVAL_50;
  wire  dcacheArb__EVAL_51;
  wire [1:0] dcacheArb__EVAL_52;
  wire  dcacheArb__EVAL_53;
  wire  dcacheArb__EVAL_54;
  wire [3:0] dcacheArb__EVAL_55;
  wire [31:0] dcacheArb__EVAL_56;
  wire  dcacheArb__EVAL_57;
  wire  dcacheArb__EVAL_58;
  wire  dcacheArb__EVAL_59;
  wire [4:0] dcacheArb__EVAL_60;
  wire [1:0] dcacheArb__EVAL_61;
  wire  dcacheArb__EVAL_62;
  wire  dcacheArb__EVAL_63;
  wire  dcacheArb__EVAL_64;
  wire  dcacheArb__EVAL_65;
  wire  dcacheArb__EVAL_66;
  wire  dcacheArb__EVAL_67;
  wire  dcacheArb__EVAL_68;
  wire  dcacheArb__EVAL_69;
  wire [6:0] dcacheArb__EVAL_70;
  wire  dcacheArb__EVAL_71;
  wire  dcacheArb__EVAL_72;
  wire  dcacheArb__EVAL_73;
  wire [31:0] dcacheArb__EVAL_74;
  wire [31:0] dcacheArb__EVAL_75;
  wire  dcacheArb__EVAL_76;
  wire  dcacheArb__EVAL_77;
  wire  dcacheArb__EVAL_78;
  wire [3:0] dcacheArb__EVAL_79;
  wire [3:0] dcacheArb__EVAL_80;
  wire [1:0] dcacheArb__EVAL_81;
  wire  dcacheArb__EVAL_82;
  wire  dcacheArb__EVAL_83;
  wire [31:0] dcacheArb__EVAL_84;
  wire [31:0] dcacheArb__EVAL_85;
  wire [3:0] _EVAL_80;
  wire  _EVAL_81;
  wire [31:0] _EVAL_82;
  wire [4:0] _EVAL_83;
  wire  frontend__EVAL;
  wire [29:0] frontend__EVAL_0;
  wire  frontend__EVAL_1;
  wire  frontend__EVAL_2;
  wire  frontend__EVAL_3;
  wire [29:0] frontend__EVAL_4;
  wire [31:0] frontend__EVAL_5;
  wire  frontend__EVAL_6;
  wire [1:0] frontend__EVAL_7;
  wire [2:0] frontend__EVAL_8;
  wire [31:0] frontend__EVAL_9;
  wire [4:0] frontend__EVAL_10;
  wire  frontend__EVAL_11;
  wire [31:0] frontend__EVAL_12;
  wire [31:0] frontend__EVAL_13;
  wire [31:0] frontend__EVAL_14;
  wire  frontend__EVAL_15;
  wire [31:0] frontend__EVAL_16;
  wire  frontend__EVAL_17;
  wire  frontend__EVAL_18;
  wire  frontend__EVAL_19;
  wire [31:0] frontend__EVAL_20;
  wire  frontend__EVAL_21;
  wire  frontend__EVAL_22;
  wire [31:0] frontend__EVAL_23;
  wire [1:0] frontend__EVAL_24;
  wire  frontend__EVAL_25;
  wire [1:0] frontend__EVAL_26;
  wire  frontend__EVAL_27;
  wire [31:0] frontend__EVAL_28;
  wire [7:0] frontend__EVAL_29;
  wire [31:0] frontend__EVAL_30;
  wire [29:0] frontend__EVAL_31;
  wire [3:0] frontend__EVAL_32;
  wire  frontend__EVAL_33;
  wire  frontend__EVAL_34;
  wire  frontend__EVAL_35;
  wire  frontend__EVAL_36;
  wire [29:0] frontend__EVAL_37;
  wire [31:0] frontend__EVAL_38;
  wire  frontend__EVAL_39;
  wire [31:0] frontend__EVAL_40;
  wire  frontend__EVAL_41;
  wire  frontend__EVAL_42;
  wire [4:0] frontend__EVAL_43;
  wire [29:0] frontend__EVAL_44;
  wire  frontend__EVAL_45;
  wire [24:0] frontend__EVAL_46;
  wire  frontend__EVAL_47;
  wire  frontend__EVAL_48;
  wire  frontend__EVAL_49;
  wire  frontend__EVAL_50;
  wire [31:0] frontend__EVAL_51;
  wire [1:0] frontend__EVAL_52;
  wire  frontend__EVAL_53;
  wire  frontend__EVAL_54;
  wire [31:0] frontend__EVAL_55;
  wire  frontend__EVAL_56;
  wire  frontend__EVAL_57;
  wire [7:0] frontend__EVAL_58;
  wire  frontend__EVAL_59;
  wire  frontend__EVAL_60;
  wire [10:0] frontend__EVAL_61;
  wire [31:0] frontend__EVAL_62;
  wire [1:0] frontend__EVAL_63;
  wire  frontend__EVAL_64;
  wire  frontend__EVAL_65;
  wire  frontend__EVAL_66;
  wire  frontend__EVAL_67;
  wire  frontend__EVAL_68;
  wire [31:0] frontend__EVAL_69;
  wire  frontend__EVAL_70;
  wire [31:0] frontend__EVAL_71;
  wire [3:0] frontend__EVAL_72;
  wire [31:0] frontend__EVAL_73;
  wire [2:0] frontend__EVAL_74;
  wire  frontend__EVAL_75;
  wire [29:0] frontend__EVAL_76;
  wire  frontend__EVAL_77;
  wire [1:0] frontend__EVAL_78;
  wire  frontend__EVAL_79;
  wire [29:0] frontend__EVAL_80;
  wire  frontend__EVAL_81;
  wire  frontend__EVAL_82;
  wire  frontend__EVAL_83;
  wire [1:0] frontend__EVAL_84;
  wire  frontend__EVAL_85;
  wire [10:0] frontend__EVAL_86;
  wire [29:0] frontend__EVAL_87;
  wire  frontend__EVAL_88;
  wire  frontend__EVAL_89;
  wire [1:0] frontend__EVAL_90;
  wire  frontend__EVAL_91;
  wire [31:0] frontend__EVAL_92;
  wire  frontend__EVAL_93;
  wire [1:0] frontend__EVAL_94;
  wire  frontend__EVAL_95;
  wire  frontend__EVAL_96;
  wire  frontend__EVAL_97;
  wire  frontend__EVAL_98;
  wire  frontend__EVAL_99;
  wire  frontend__EVAL_100;
  wire  frontend__EVAL_101;
  wire [31:0] frontend__EVAL_102;
  wire [31:0] frontend__EVAL_103;
  wire  frontend__EVAL_104;
  wire [2:0] frontend__EVAL_105;
  wire  frontend__EVAL_106;
  wire [1:0] frontend__EVAL_107;
  wire [1:0] frontend__EVAL_108;
  wire [31:0] frontend__EVAL_109;
  wire [1:0] frontend__EVAL_110;
  wire  frontend__EVAL_111;
  wire  frontend__EVAL_112;
  wire  frontend__EVAL_113;
  wire  frontend__EVAL_114;
  wire [1:0] frontend__EVAL_115;
  wire  frontend__EVAL_116;
  wire  frontend__EVAL_117;
  wire  frontend__EVAL_118;
  wire  frontend__EVAL_119;
  wire  frontend__EVAL_120;
  wire  _EVAL_85;
  wire  _EVAL_86;
  reg  _EVAL_87;
  wire [31:0] _EVAL_88;
  wire  tlSlaveXbar__EVAL;
  wire [2:0] tlSlaveXbar__EVAL_0;
  wire [31:0] tlSlaveXbar__EVAL_1;
  wire [31:0] tlSlaveXbar__EVAL_2;
  wire  tlSlaveXbar__EVAL_3;
  wire [2:0] tlSlaveXbar__EVAL_4;
  wire [4:0] tlSlaveXbar__EVAL_5;
  wire [31:0] tlSlaveXbar__EVAL_6;
  wire [24:0] tlSlaveXbar__EVAL_7;
  wire [31:0] tlSlaveXbar__EVAL_8;
  wire [2:0] tlSlaveXbar__EVAL_9;
  wire [4:0] tlSlaveXbar__EVAL_10;
  wire [2:0] tlSlaveXbar__EVAL_11;
  wire [4:0] tlSlaveXbar__EVAL_12;
  wire [31:0] tlSlaveXbar__EVAL_13;
  wire [31:0] tlSlaveXbar__EVAL_14;
  wire  tlSlaveXbar__EVAL_15;
  wire  tlSlaveXbar__EVAL_16;
  wire [2:0] tlSlaveXbar__EVAL_17;
  wire [2:0] tlSlaveXbar__EVAL_18;
  wire [2:0] tlSlaveXbar__EVAL_19;
  wire [2:0] tlSlaveXbar__EVAL_20;
  wire [2:0] tlSlaveXbar__EVAL_21;
  wire  tlSlaveXbar__EVAL_22;
  wire  tlSlaveXbar__EVAL_23;
  wire [4:0] tlSlaveXbar__EVAL_24;
  wire [4:0] tlSlaveXbar__EVAL_25;
  wire [2:0] tlSlaveXbar__EVAL_26;
  wire [2:0] tlSlaveXbar__EVAL_27;
  wire  tlSlaveXbar__EVAL_28;
  wire  tlSlaveXbar__EVAL_29;
  wire  tlSlaveXbar__EVAL_30;
  wire  tlSlaveXbar__EVAL_31;
  wire [31:0] tlSlaveXbar__EVAL_32;
  wire [3:0] tlSlaveXbar__EVAL_33;
  wire  tlSlaveXbar__EVAL_34;
  wire  tlSlaveXbar__EVAL_35;
  wire [3:0] tlSlaveXbar__EVAL_36;
  wire [3:0] tlSlaveXbar__EVAL_37;
  wire  tlSlaveXbar__EVAL_38;
  wire [31:0] tlSlaveXbar__EVAL_39;
  wire  tlSlaveXbar__EVAL_40;
  wire [2:0] tlSlaveXbar__EVAL_41;
  wire [2:0] tlSlaveXbar__EVAL_42;
  wire [4:0] tlSlaveXbar__EVAL_43;
  wire [2:0] tlSlaveXbar__EVAL_44;
  wire  core__EVAL;
  wire  core__EVAL_0;
  wire [31:0] core__EVAL_1;
  wire [6:0] core__EVAL_2;
  wire  core__EVAL_3;
  wire  core__EVAL_4;
  wire  core__EVAL_5;
  wire  core__EVAL_6;
  wire  core__EVAL_7;
  wire  core__EVAL_8;
  wire [4:0] core__EVAL_9;
  wire  core__EVAL_10;
  wire [1:0] core__EVAL_11;
  wire  core__EVAL_12;
  wire  core__EVAL_13;
  wire  core__EVAL_14;
  wire [31:0] core__EVAL_15;
  wire [3:0] core__EVAL_16;
  wire  core__EVAL_17;
  wire  core__EVAL_18;
  wire  core__EVAL_19;
  wire [31:0] core__EVAL_20;
  wire  core__EVAL_21;
  wire [1:0] core__EVAL_22;
  wire  core__EVAL_23;
  wire  core__EVAL_24;
  wire [29:0] core__EVAL_25;
  wire [1:0] core__EVAL_26;
  wire [31:0] core__EVAL_27;
  wire  core__EVAL_28;
  wire [31:0] core__EVAL_29;
  wire [29:0] core__EVAL_30;
  wire  core__EVAL_31;
  wire  core__EVAL_32;
  wire [1:0] core__EVAL_33;
  wire [1:0] core__EVAL_34;
  wire [1:0] core__EVAL_35;
  wire [31:0] core__EVAL_36;
  wire  core__EVAL_37;
  wire [29:0] core__EVAL_38;
  wire  core__EVAL_39;
  wire  core__EVAL_40;
  wire  core__EVAL_41;
  wire  core__EVAL_42;
  wire [4:0] core__EVAL_43;
  wire [31:0] core__EVAL_44;
  wire [4:0] core__EVAL_45;
  wire [1:0] core__EVAL_46;
  wire  core__EVAL_47;
  wire [31:0] core__EVAL_48;
  wire [1:0] core__EVAL_49;
  wire  core__EVAL_50;
  wire [31:0] core__EVAL_51;
  wire  core__EVAL_52;
  wire  core__EVAL_53;
  wire [1:0] core__EVAL_54;
  wire  core__EVAL_55;
  wire  core__EVAL_56;
  wire  core__EVAL_57;
  wire  core__EVAL_58;
  wire  core__EVAL_59;
  wire [4:0] core__EVAL_60;
  wire  core__EVAL_61;
  wire [31:0] core__EVAL_62;
  wire  core__EVAL_63;
  wire [1:0] core__EVAL_64;
  wire  core__EVAL_65;
  wire [31:0] core__EVAL_66;
  wire  core__EVAL_67;
  wire [1:0] core__EVAL_68;
  wire [31:0] core__EVAL_69;
  wire [1:0] core__EVAL_70;
  wire [7:0] core__EVAL_71;
  wire [31:0] core__EVAL_72;
  wire  core__EVAL_73;
  wire  core__EVAL_74;
  wire [31:0] core__EVAL_75;
  wire [6:0] core__EVAL_76;
  wire  core__EVAL_77;
  wire  core__EVAL_78;
  wire  core__EVAL_79;
  wire  core__EVAL_80;
  wire  core__EVAL_81;
  wire  core__EVAL_82;
  wire  core__EVAL_83;
  wire  core__EVAL_84;
  wire  core__EVAL_85;
  wire  core__EVAL_86;
  wire  core__EVAL_87;
  wire  core__EVAL_88;
  wire [1:0] core__EVAL_89;
  wire  core__EVAL_90;
  wire [31:0] core__EVAL_91;
  wire  core__EVAL_92;
  wire  core__EVAL_93;
  wire  core__EVAL_94;
  wire [31:0] core__EVAL_95;
  wire  core__EVAL_96;
  wire  core__EVAL_97;
  wire  core__EVAL_98;
  wire  core__EVAL_99;
  wire  core__EVAL_100;
  wire  core__EVAL_101;
  wire  core__EVAL_102;
  wire  core__EVAL_103;
  wire [31:0] core__EVAL_104;
  wire  core__EVAL_105;
  wire  core__EVAL_106;
  wire  core__EVAL_107;
  wire [31:0] core__EVAL_108;
  wire  core__EVAL_109;
  wire [1:0] core__EVAL_110;
  wire  core__EVAL_111;
  wire [31:0] core__EVAL_112;
  wire [31:0] core__EVAL_113;
  wire  core__EVAL_114;
  wire  core__EVAL_115;
  wire  core__EVAL_116;
  wire  core__EVAL_117;
  wire  core__EVAL_118;
  wire  core__EVAL_119;
  wire  core__EVAL_120;
  wire  core__EVAL_121;
  wire  core__EVAL_122;
  wire  core__EVAL_123;
  wire  core__EVAL_124;
  wire [31:0] core__EVAL_125;
  wire  core__EVAL_126;
  wire  core__EVAL_127;
  wire [7:0] core__EVAL_128;
  wire  core__EVAL_129;
  wire  core__EVAL_130;
  wire  core__EVAL_131;
  wire  core__EVAL_132;
  wire [29:0] core__EVAL_133;
  wire  core__EVAL_134;
  wire  core__EVAL_135;
  wire [29:0] core__EVAL_136;
  wire  core__EVAL_137;
  wire [29:0] core__EVAL_138;
  wire  core__EVAL_139;
  wire  core__EVAL_140;
  wire  core__EVAL_141;
  wire [1:0] core__EVAL_142;
  wire  core__EVAL_143;
  wire  core__EVAL_144;
  wire  core__EVAL_145;
  wire [31:0] core__EVAL_146;
  wire  core__EVAL_147;
  wire [31:0] core__EVAL_148;
  wire  core__EVAL_149;
  wire  core__EVAL_150;
  wire  core__EVAL_151;
  wire [31:0] core__EVAL_152;
  wire [3:0] core__EVAL_153;
  wire  core__EVAL_154;
  wire [29:0] core__EVAL_155;
  wire [29:0] core__EVAL_156;
  wire  core__EVAL_157;
  wire  core__EVAL_158;
  wire  core__EVAL_159;
  wire  core__EVAL_160;
  wire  core__EVAL_161;
  reg [3:0] _EVAL_91;
  wire  fragmenter__EVAL;
  wire [2:0] fragmenter__EVAL_0;
  wire [2:0] fragmenter__EVAL_1;
  wire [2:0] fragmenter__EVAL_2;
  wire [2:0] fragmenter__EVAL_3;
  wire  fragmenter__EVAL_4;
  wire [24:0] fragmenter__EVAL_5;
  wire  fragmenter__EVAL_6;
  wire [3:0] fragmenter__EVAL_7;
  wire  fragmenter__EVAL_8;
  wire [1:0] fragmenter__EVAL_9;
  wire [31:0] fragmenter__EVAL_10;
  wire  fragmenter__EVAL_11;
  wire [4:0] fragmenter__EVAL_12;
  wire [31:0] fragmenter__EVAL_13;
  wire [2:0] fragmenter__EVAL_14;
  wire [31:0] fragmenter__EVAL_15;
  wire [24:0] fragmenter__EVAL_16;
  wire  fragmenter__EVAL_17;
  wire [31:0] fragmenter__EVAL_18;
  wire [2:0] fragmenter__EVAL_19;
  wire [3:0] fragmenter__EVAL_20;
  wire [10:0] fragmenter__EVAL_21;
  wire [4:0] fragmenter__EVAL_22;
  wire  fragmenter__EVAL_23;
  wire  fragmenter__EVAL_24;
  wire  fragmenter__EVAL_25;
  wire [1:0] fragmenter__EVAL_26;
  wire [10:0] fragmenter__EVAL_27;
  wire  fragmenter__EVAL_28;
  wire [31:0] _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire [31:0] _EVAL_97;
  _EVAL_110 dcache (
    ._EVAL(dcache__EVAL),
    ._EVAL_0(dcache__EVAL_0),
    ._EVAL_1(dcache__EVAL_1),
    ._EVAL_2(dcache__EVAL_2),
    ._EVAL_3(dcache__EVAL_3),
    ._EVAL_4(dcache__EVAL_4),
    ._EVAL_5(dcache__EVAL_5),
    ._EVAL_6(dcache__EVAL_6),
    ._EVAL_7(dcache__EVAL_7),
    ._EVAL_8(dcache__EVAL_8),
    ._EVAL_9(dcache__EVAL_9),
    ._EVAL_10(dcache__EVAL_10),
    ._EVAL_11(dcache__EVAL_11),
    ._EVAL_12(dcache__EVAL_12),
    ._EVAL_13(dcache__EVAL_13),
    ._EVAL_14(dcache__EVAL_14),
    ._EVAL_15(dcache__EVAL_15),
    ._EVAL_16(dcache__EVAL_16),
    ._EVAL_17(dcache__EVAL_17),
    ._EVAL_18(dcache__EVAL_18),
    ._EVAL_19(dcache__EVAL_19),
    ._EVAL_20(dcache__EVAL_20),
    ._EVAL_21(dcache__EVAL_21),
    ._EVAL_22(dcache__EVAL_22),
    ._EVAL_23(dcache__EVAL_23),
    ._EVAL_24(dcache__EVAL_24),
    ._EVAL_25(dcache__EVAL_25),
    ._EVAL_26(dcache__EVAL_26),
    ._EVAL_27(dcache__EVAL_27),
    ._EVAL_28(dcache__EVAL_28),
    ._EVAL_29(dcache__EVAL_29),
    ._EVAL_30(dcache__EVAL_30),
    ._EVAL_31(dcache__EVAL_31),
    ._EVAL_32(dcache__EVAL_32),
    ._EVAL_33(dcache__EVAL_33),
    ._EVAL_34(dcache__EVAL_34),
    ._EVAL_35(dcache__EVAL_35),
    ._EVAL_36(dcache__EVAL_36),
    ._EVAL_37(dcache__EVAL_37),
    ._EVAL_38(dcache__EVAL_38),
    ._EVAL_39(dcache__EVAL_39),
    ._EVAL_40(dcache__EVAL_40),
    ._EVAL_41(dcache__EVAL_41),
    ._EVAL_42(dcache__EVAL_42),
    ._EVAL_43(dcache__EVAL_43),
    ._EVAL_44(dcache__EVAL_44),
    ._EVAL_45(dcache__EVAL_45),
    ._EVAL_46(dcache__EVAL_46),
    ._EVAL_47(dcache__EVAL_47),
    ._EVAL_48(dcache__EVAL_48),
    ._EVAL_49(dcache__EVAL_49),
    ._EVAL_50(dcache__EVAL_50),
    ._EVAL_51(dcache__EVAL_51),
    ._EVAL_52(dcache__EVAL_52),
    ._EVAL_53(dcache__EVAL_53),
    ._EVAL_54(dcache__EVAL_54),
    ._EVAL_55(dcache__EVAL_55),
    ._EVAL_56(dcache__EVAL_56),
    ._EVAL_57(dcache__EVAL_57),
    ._EVAL_58(dcache__EVAL_58),
    ._EVAL_59(dcache__EVAL_59),
    ._EVAL_60(dcache__EVAL_60),
    ._EVAL_61(dcache__EVAL_61),
    ._EVAL_62(dcache__EVAL_62),
    ._EVAL_63(dcache__EVAL_63),
    ._EVAL_64(dcache__EVAL_64),
    ._EVAL_65(dcache__EVAL_65),
    ._EVAL_66(dcache__EVAL_66),
    ._EVAL_67(dcache__EVAL_67),
    ._EVAL_68(dcache__EVAL_68),
    ._EVAL_69(dcache__EVAL_69),
    ._EVAL_70(dcache__EVAL_70),
    ._EVAL_71(dcache__EVAL_71),
    ._EVAL_72(dcache__EVAL_72),
    ._EVAL_73(dcache__EVAL_73),
    ._EVAL_74(dcache__EVAL_74),
    ._EVAL_75(dcache__EVAL_75),
    ._EVAL_76(dcache__EVAL_76),
    ._EVAL_77(dcache__EVAL_77),
    ._EVAL_78(dcache__EVAL_78),
    ._EVAL_79(dcache__EVAL_79),
    ._EVAL_80(dcache__EVAL_80),
    ._EVAL_81(dcache__EVAL_81),
    ._EVAL_82(dcache__EVAL_82),
    ._EVAL_83(dcache__EVAL_83),
    ._EVAL_84(dcache__EVAL_84),
    ._EVAL_85(dcache__EVAL_85),
    ._EVAL_86(dcache__EVAL_86),
    ._EVAL_87(dcache__EVAL_87),
    ._EVAL_88(dcache__EVAL_88),
    ._EVAL_89(dcache__EVAL_89),
    ._EVAL_90(dcache__EVAL_90),
    ._EVAL_91(dcache__EVAL_91),
    ._EVAL_92(dcache__EVAL_92),
    ._EVAL_93(dcache__EVAL_93),
    ._EVAL_94(dcache__EVAL_94),
    ._EVAL_95(dcache__EVAL_95),
    ._EVAL_96(dcache__EVAL_96),
    ._EVAL_97(dcache__EVAL_97),
    ._EVAL_98(dcache__EVAL_98),
    ._EVAL_99(dcache__EVAL_99),
    ._EVAL_100(dcache__EVAL_100),
    ._EVAL_101(dcache__EVAL_101),
    ._EVAL_102(dcache__EVAL_102),
    ._EVAL_103(dcache__EVAL_103),
    ._EVAL_104(dcache__EVAL_104),
    ._EVAL_105(dcache__EVAL_105),
    ._EVAL_106(dcache__EVAL_106),
    ._EVAL_107(dcache__EVAL_107),
    ._EVAL_108(dcache__EVAL_108),
    ._EVAL_109(dcache__EVAL_109),
    ._EVAL_110(dcache__EVAL_110),
    ._EVAL_111(dcache__EVAL_111),
    ._EVAL_112(dcache__EVAL_112),
    ._EVAL_113(dcache__EVAL_113),
    ._EVAL_114(dcache__EVAL_114),
    ._EVAL_115(dcache__EVAL_115),
    ._EVAL_116(dcache__EVAL_116),
    ._EVAL_117(dcache__EVAL_117),
    ._EVAL_118(dcache__EVAL_118),
    ._EVAL_119(dcache__EVAL_119),
    ._EVAL_120(dcache__EVAL_120),
    ._EVAL_121(dcache__EVAL_121),
    ._EVAL_122(dcache__EVAL_122),
    ._EVAL_123(dcache__EVAL_123),
    ._EVAL_124(dcache__EVAL_124),
    ._EVAL_125(dcache__EVAL_125),
    ._EVAL_126(dcache__EVAL_126),
    ._EVAL_127(dcache__EVAL_127),
    ._EVAL_128(dcache__EVAL_128)
  );
  _EVAL_118 dtim_adapter (
    ._EVAL(dtim_adapter__EVAL),
    ._EVAL_0(dtim_adapter__EVAL_0),
    ._EVAL_1(dtim_adapter__EVAL_1),
    ._EVAL_2(dtim_adapter__EVAL_2),
    ._EVAL_3(dtim_adapter__EVAL_3),
    ._EVAL_4(dtim_adapter__EVAL_4),
    ._EVAL_5(dtim_adapter__EVAL_5),
    ._EVAL_6(dtim_adapter__EVAL_6),
    ._EVAL_7(dtim_adapter__EVAL_7),
    ._EVAL_8(dtim_adapter__EVAL_8),
    ._EVAL_9(dtim_adapter__EVAL_9),
    ._EVAL_10(dtim_adapter__EVAL_10),
    ._EVAL_11(dtim_adapter__EVAL_11),
    ._EVAL_12(dtim_adapter__EVAL_12),
    ._EVAL_13(dtim_adapter__EVAL_13),
    ._EVAL_14(dtim_adapter__EVAL_14),
    ._EVAL_15(dtim_adapter__EVAL_15),
    ._EVAL_16(dtim_adapter__EVAL_16),
    ._EVAL_17(dtim_adapter__EVAL_17),
    ._EVAL_18(dtim_adapter__EVAL_18),
    ._EVAL_19(dtim_adapter__EVAL_19),
    ._EVAL_20(dtim_adapter__EVAL_20),
    ._EVAL_21(dtim_adapter__EVAL_21),
    ._EVAL_22(dtim_adapter__EVAL_22),
    ._EVAL_23(dtim_adapter__EVAL_23),
    ._EVAL_24(dtim_adapter__EVAL_24),
    ._EVAL_25(dtim_adapter__EVAL_25),
    ._EVAL_26(dtim_adapter__EVAL_26)
  );
  _EVAL_103 tlMasterXbar (
    ._EVAL(tlMasterXbar__EVAL),
    ._EVAL_0(tlMasterXbar__EVAL_0),
    ._EVAL_1(tlMasterXbar__EVAL_1),
    ._EVAL_2(tlMasterXbar__EVAL_2),
    ._EVAL_3(tlMasterXbar__EVAL_3),
    ._EVAL_4(tlMasterXbar__EVAL_4),
    ._EVAL_5(tlMasterXbar__EVAL_5),
    ._EVAL_6(tlMasterXbar__EVAL_6),
    ._EVAL_7(tlMasterXbar__EVAL_7),
    ._EVAL_8(tlMasterXbar__EVAL_8),
    ._EVAL_9(tlMasterXbar__EVAL_9),
    ._EVAL_10(tlMasterXbar__EVAL_10),
    ._EVAL_11(tlMasterXbar__EVAL_11),
    ._EVAL_12(tlMasterXbar__EVAL_12),
    ._EVAL_13(tlMasterXbar__EVAL_13),
    ._EVAL_14(tlMasterXbar__EVAL_14),
    ._EVAL_15(tlMasterXbar__EVAL_15),
    ._EVAL_16(tlMasterXbar__EVAL_16),
    ._EVAL_17(tlMasterXbar__EVAL_17),
    ._EVAL_18(tlMasterXbar__EVAL_18),
    ._EVAL_19(tlMasterXbar__EVAL_19),
    ._EVAL_20(tlMasterXbar__EVAL_20),
    ._EVAL_21(tlMasterXbar__EVAL_21),
    ._EVAL_22(tlMasterXbar__EVAL_22),
    ._EVAL_23(tlMasterXbar__EVAL_23),
    ._EVAL_24(tlMasterXbar__EVAL_24),
    ._EVAL_25(tlMasterXbar__EVAL_25),
    ._EVAL_26(tlMasterXbar__EVAL_26),
    ._EVAL_27(tlMasterXbar__EVAL_27),
    ._EVAL_28(tlMasterXbar__EVAL_28),
    ._EVAL_29(tlMasterXbar__EVAL_29),
    ._EVAL_30(tlMasterXbar__EVAL_30),
    ._EVAL_31(tlMasterXbar__EVAL_31),
    ._EVAL_32(tlMasterXbar__EVAL_32),
    ._EVAL_33(tlMasterXbar__EVAL_33),
    ._EVAL_34(tlMasterXbar__EVAL_34),
    ._EVAL_35(tlMasterXbar__EVAL_35),
    ._EVAL_36(tlMasterXbar__EVAL_36),
    ._EVAL_37(tlMasterXbar__EVAL_37),
    ._EVAL_38(tlMasterXbar__EVAL_38),
    ._EVAL_39(tlMasterXbar__EVAL_39),
    ._EVAL_40(tlMasterXbar__EVAL_40),
    ._EVAL_41(tlMasterXbar__EVAL_41),
    ._EVAL_42(tlMasterXbar__EVAL_42),
    ._EVAL_43(tlMasterXbar__EVAL_43),
    ._EVAL_44(tlMasterXbar__EVAL_44),
    ._EVAL_45(tlMasterXbar__EVAL_45),
    ._EVAL_46(tlMasterXbar__EVAL_46),
    ._EVAL_47(tlMasterXbar__EVAL_47),
    ._EVAL_48(tlMasterXbar__EVAL_48),
    ._EVAL_49(tlMasterXbar__EVAL_49),
    ._EVAL_50(tlMasterXbar__EVAL_50),
    ._EVAL_51(tlMasterXbar__EVAL_51),
    ._EVAL_52(tlMasterXbar__EVAL_52),
    ._EVAL_53(tlMasterXbar__EVAL_53),
    ._EVAL_54(tlMasterXbar__EVAL_54),
    ._EVAL_55(tlMasterXbar__EVAL_55),
    ._EVAL_56(tlMasterXbar__EVAL_56),
    ._EVAL_57(tlMasterXbar__EVAL_57)
  );
  _EVAL_120 fragmenter_1 (
    ._EVAL(fragmenter_1__EVAL),
    ._EVAL_0(fragmenter_1__EVAL_0),
    ._EVAL_1(fragmenter_1__EVAL_1),
    ._EVAL_2(fragmenter_1__EVAL_2),
    ._EVAL_3(fragmenter_1__EVAL_3),
    ._EVAL_4(fragmenter_1__EVAL_4),
    ._EVAL_5(fragmenter_1__EVAL_5),
    ._EVAL_6(fragmenter_1__EVAL_6),
    ._EVAL_7(fragmenter_1__EVAL_7),
    ._EVAL_8(fragmenter_1__EVAL_8),
    ._EVAL_9(fragmenter_1__EVAL_9),
    ._EVAL_10(fragmenter_1__EVAL_10),
    ._EVAL_11(fragmenter_1__EVAL_11),
    ._EVAL_12(fragmenter_1__EVAL_12),
    ._EVAL_13(fragmenter_1__EVAL_13),
    ._EVAL_14(fragmenter_1__EVAL_14),
    ._EVAL_15(fragmenter_1__EVAL_15),
    ._EVAL_16(fragmenter_1__EVAL_16),
    ._EVAL_17(fragmenter_1__EVAL_17),
    ._EVAL_18(fragmenter_1__EVAL_18),
    ._EVAL_19(fragmenter_1__EVAL_19),
    ._EVAL_20(fragmenter_1__EVAL_20),
    ._EVAL_21(fragmenter_1__EVAL_21),
    ._EVAL_22(fragmenter_1__EVAL_22),
    ._EVAL_23(fragmenter_1__EVAL_23),
    ._EVAL_24(fragmenter_1__EVAL_24),
    ._EVAL_25(fragmenter_1__EVAL_25),
    ._EVAL_26(fragmenter_1__EVAL_26),
    ._EVAL_27(fragmenter_1__EVAL_27),
    ._EVAL_28(fragmenter_1__EVAL_28),
    ._EVAL_29(fragmenter_1__EVAL_29),
    ._EVAL_30(fragmenter_1__EVAL_30)
  );
  _EVAL_124 ptw (
    ._EVAL(ptw__EVAL),
    ._EVAL_0(ptw__EVAL_0),
    ._EVAL_1(ptw__EVAL_1),
    ._EVAL_2(ptw__EVAL_2),
    ._EVAL_3(ptw__EVAL_3),
    ._EVAL_4(ptw__EVAL_4),
    ._EVAL_5(ptw__EVAL_5),
    ._EVAL_6(ptw__EVAL_6),
    ._EVAL_7(ptw__EVAL_7),
    ._EVAL_8(ptw__EVAL_8),
    ._EVAL_9(ptw__EVAL_9),
    ._EVAL_10(ptw__EVAL_10),
    ._EVAL_11(ptw__EVAL_11),
    ._EVAL_12(ptw__EVAL_12),
    ._EVAL_13(ptw__EVAL_13),
    ._EVAL_14(ptw__EVAL_14),
    ._EVAL_15(ptw__EVAL_15),
    ._EVAL_16(ptw__EVAL_16),
    ._EVAL_17(ptw__EVAL_17),
    ._EVAL_18(ptw__EVAL_18),
    ._EVAL_19(ptw__EVAL_19),
    ._EVAL_20(ptw__EVAL_20),
    ._EVAL_21(ptw__EVAL_21),
    ._EVAL_22(ptw__EVAL_22),
    ._EVAL_23(ptw__EVAL_23),
    ._EVAL_24(ptw__EVAL_24),
    ._EVAL_25(ptw__EVAL_25),
    ._EVAL_26(ptw__EVAL_26),
    ._EVAL_27(ptw__EVAL_27),
    ._EVAL_28(ptw__EVAL_28),
    ._EVAL_29(ptw__EVAL_29),
    ._EVAL_30(ptw__EVAL_30),
    ._EVAL_31(ptw__EVAL_31),
    ._EVAL_32(ptw__EVAL_32),
    ._EVAL_33(ptw__EVAL_33),
    ._EVAL_34(ptw__EVAL_34),
    ._EVAL_35(ptw__EVAL_35),
    ._EVAL_36(ptw__EVAL_36),
    ._EVAL_37(ptw__EVAL_37),
    ._EVAL_38(ptw__EVAL_38),
    ._EVAL_39(ptw__EVAL_39),
    ._EVAL_40(ptw__EVAL_40),
    ._EVAL_41(ptw__EVAL_41),
    ._EVAL_42(ptw__EVAL_42),
    ._EVAL_43(ptw__EVAL_43),
    ._EVAL_44(ptw__EVAL_44),
    ._EVAL_45(ptw__EVAL_45),
    ._EVAL_46(ptw__EVAL_46),
    ._EVAL_47(ptw__EVAL_47),
    ._EVAL_48(ptw__EVAL_48),
    ._EVAL_49(ptw__EVAL_49),
    ._EVAL_50(ptw__EVAL_50),
    ._EVAL_51(ptw__EVAL_51),
    ._EVAL_52(ptw__EVAL_52),
    ._EVAL_53(ptw__EVAL_53),
    ._EVAL_54(ptw__EVAL_54),
    ._EVAL_55(ptw__EVAL_55),
    ._EVAL_56(ptw__EVAL_56),
    ._EVAL_57(ptw__EVAL_57),
    ._EVAL_58(ptw__EVAL_58),
    ._EVAL_59(ptw__EVAL_59),
    ._EVAL_60(ptw__EVAL_60),
    ._EVAL_61(ptw__EVAL_61),
    ._EVAL_62(ptw__EVAL_62),
    ._EVAL_63(ptw__EVAL_63),
    ._EVAL_64(ptw__EVAL_64),
    ._EVAL_65(ptw__EVAL_65),
    ._EVAL_66(ptw__EVAL_66),
    ._EVAL_67(ptw__EVAL_67),
    ._EVAL_68(ptw__EVAL_68),
    ._EVAL_69(ptw__EVAL_69),
    ._EVAL_70(ptw__EVAL_70),
    ._EVAL_71(ptw__EVAL_71),
    ._EVAL_72(ptw__EVAL_72),
    ._EVAL_73(ptw__EVAL_73),
    ._EVAL_74(ptw__EVAL_74),
    ._EVAL_75(ptw__EVAL_75),
    ._EVAL_76(ptw__EVAL_76),
    ._EVAL_77(ptw__EVAL_77),
    ._EVAL_78(ptw__EVAL_78),
    ._EVAL_79(ptw__EVAL_79),
    ._EVAL_80(ptw__EVAL_80),
    ._EVAL_81(ptw__EVAL_81),
    ._EVAL_82(ptw__EVAL_82),
    ._EVAL_83(ptw__EVAL_83),
    ._EVAL_84(ptw__EVAL_84),
    ._EVAL_85(ptw__EVAL_85),
    ._EVAL_86(ptw__EVAL_86),
    ._EVAL_87(ptw__EVAL_87),
    ._EVAL_88(ptw__EVAL_88),
    ._EVAL_89(ptw__EVAL_89),
    ._EVAL_90(ptw__EVAL_90),
    ._EVAL_91(ptw__EVAL_91),
    ._EVAL_92(ptw__EVAL_92),
    ._EVAL_93(ptw__EVAL_93),
    ._EVAL_94(ptw__EVAL_94),
    ._EVAL_95(ptw__EVAL_95),
    ._EVAL_96(ptw__EVAL_96),
    ._EVAL_97(ptw__EVAL_97),
    ._EVAL_98(ptw__EVAL_98),
    ._EVAL_99(ptw__EVAL_99),
    ._EVAL_100(ptw__EVAL_100),
    ._EVAL_101(ptw__EVAL_101),
    ._EVAL_102(ptw__EVAL_102),
    ._EVAL_103(ptw__EVAL_103),
    ._EVAL_104(ptw__EVAL_104),
    ._EVAL_105(ptw__EVAL_105),
    ._EVAL_106(ptw__EVAL_106),
    ._EVAL_107(ptw__EVAL_107),
    ._EVAL_108(ptw__EVAL_108),
    ._EVAL_109(ptw__EVAL_109),
    ._EVAL_110(ptw__EVAL_110),
    ._EVAL_111(ptw__EVAL_111),
    ._EVAL_112(ptw__EVAL_112),
    ._EVAL_113(ptw__EVAL_113),
    ._EVAL_114(ptw__EVAL_114),
    ._EVAL_115(ptw__EVAL_115),
    ._EVAL_116(ptw__EVAL_116),
    ._EVAL_117(ptw__EVAL_117),
    ._EVAL_118(ptw__EVAL_118),
    ._EVAL_119(ptw__EVAL_119),
    ._EVAL_120(ptw__EVAL_120),
    ._EVAL_121(ptw__EVAL_121),
    ._EVAL_122(ptw__EVAL_122),
    ._EVAL_123(ptw__EVAL_123),
    ._EVAL_124(ptw__EVAL_124),
    ._EVAL_125(ptw__EVAL_125),
    ._EVAL_126(ptw__EVAL_126),
    ._EVAL_127(ptw__EVAL_127),
    ._EVAL_128(ptw__EVAL_128),
    ._EVAL_129(ptw__EVAL_129),
    ._EVAL_130(ptw__EVAL_130),
    ._EVAL_131(ptw__EVAL_131),
    ._EVAL_132(ptw__EVAL_132),
    ._EVAL_133(ptw__EVAL_133),
    ._EVAL_134(ptw__EVAL_134),
    ._EVAL_135(ptw__EVAL_135),
    ._EVAL_136(ptw__EVAL_136),
    ._EVAL_137(ptw__EVAL_137),
    ._EVAL_138(ptw__EVAL_138),
    ._EVAL_139(ptw__EVAL_139),
    ._EVAL_140(ptw__EVAL_140),
    ._EVAL_141(ptw__EVAL_141),
    ._EVAL_142(ptw__EVAL_142),
    ._EVAL_143(ptw__EVAL_143),
    ._EVAL_144(ptw__EVAL_144),
    ._EVAL_145(ptw__EVAL_145),
    ._EVAL_146(ptw__EVAL_146),
    ._EVAL_147(ptw__EVAL_147),
    ._EVAL_148(ptw__EVAL_148),
    ._EVAL_149(ptw__EVAL_149),
    ._EVAL_150(ptw__EVAL_150),
    ._EVAL_151(ptw__EVAL_151),
    ._EVAL_152(ptw__EVAL_152),
    ._EVAL_153(ptw__EVAL_153),
    ._EVAL_154(ptw__EVAL_154),
    ._EVAL_155(ptw__EVAL_155),
    ._EVAL_156(ptw__EVAL_156),
    ._EVAL_157(ptw__EVAL_157),
    ._EVAL_158(ptw__EVAL_158),
    ._EVAL_159(ptw__EVAL_159),
    ._EVAL_160(ptw__EVAL_160),
    ._EVAL_161(ptw__EVAL_161),
    ._EVAL_162(ptw__EVAL_162),
    ._EVAL_163(ptw__EVAL_163),
    ._EVAL_164(ptw__EVAL_164),
    ._EVAL_165(ptw__EVAL_165),
    ._EVAL_166(ptw__EVAL_166),
    ._EVAL_167(ptw__EVAL_167),
    ._EVAL_168(ptw__EVAL_168),
    ._EVAL_169(ptw__EVAL_169),
    ._EVAL_170(ptw__EVAL_170),
    ._EVAL_171(ptw__EVAL_171),
    ._EVAL_172(ptw__EVAL_172),
    ._EVAL_173(ptw__EVAL_173),
    ._EVAL_174(ptw__EVAL_174),
    ._EVAL_175(ptw__EVAL_175),
    ._EVAL_176(ptw__EVAL_176),
    ._EVAL_177(ptw__EVAL_177),
    ._EVAL_178(ptw__EVAL_178),
    ._EVAL_179(ptw__EVAL_179),
    ._EVAL_180(ptw__EVAL_180),
    ._EVAL_181(ptw__EVAL_181),
    ._EVAL_182(ptw__EVAL_182),
    ._EVAL_183(ptw__EVAL_183),
    ._EVAL_184(ptw__EVAL_184),
    ._EVAL_185(ptw__EVAL_185),
    ._EVAL_186(ptw__EVAL_186),
    ._EVAL_187(ptw__EVAL_187)
  );
  _EVAL_121 dcacheArb (
    ._EVAL(dcacheArb__EVAL),
    ._EVAL_0(dcacheArb__EVAL_0),
    ._EVAL_1(dcacheArb__EVAL_1),
    ._EVAL_2(dcacheArb__EVAL_2),
    ._EVAL_3(dcacheArb__EVAL_3),
    ._EVAL_4(dcacheArb__EVAL_4),
    ._EVAL_5(dcacheArb__EVAL_5),
    ._EVAL_6(dcacheArb__EVAL_6),
    ._EVAL_7(dcacheArb__EVAL_7),
    ._EVAL_8(dcacheArb__EVAL_8),
    ._EVAL_9(dcacheArb__EVAL_9),
    ._EVAL_10(dcacheArb__EVAL_10),
    ._EVAL_11(dcacheArb__EVAL_11),
    ._EVAL_12(dcacheArb__EVAL_12),
    ._EVAL_13(dcacheArb__EVAL_13),
    ._EVAL_14(dcacheArb__EVAL_14),
    ._EVAL_15(dcacheArb__EVAL_15),
    ._EVAL_16(dcacheArb__EVAL_16),
    ._EVAL_17(dcacheArb__EVAL_17),
    ._EVAL_18(dcacheArb__EVAL_18),
    ._EVAL_19(dcacheArb__EVAL_19),
    ._EVAL_20(dcacheArb__EVAL_20),
    ._EVAL_21(dcacheArb__EVAL_21),
    ._EVAL_22(dcacheArb__EVAL_22),
    ._EVAL_23(dcacheArb__EVAL_23),
    ._EVAL_24(dcacheArb__EVAL_24),
    ._EVAL_25(dcacheArb__EVAL_25),
    ._EVAL_26(dcacheArb__EVAL_26),
    ._EVAL_27(dcacheArb__EVAL_27),
    ._EVAL_28(dcacheArb__EVAL_28),
    ._EVAL_29(dcacheArb__EVAL_29),
    ._EVAL_30(dcacheArb__EVAL_30),
    ._EVAL_31(dcacheArb__EVAL_31),
    ._EVAL_32(dcacheArb__EVAL_32),
    ._EVAL_33(dcacheArb__EVAL_33),
    ._EVAL_34(dcacheArb__EVAL_34),
    ._EVAL_35(dcacheArb__EVAL_35),
    ._EVAL_36(dcacheArb__EVAL_36),
    ._EVAL_37(dcacheArb__EVAL_37),
    ._EVAL_38(dcacheArb__EVAL_38),
    ._EVAL_39(dcacheArb__EVAL_39),
    ._EVAL_40(dcacheArb__EVAL_40),
    ._EVAL_41(dcacheArb__EVAL_41),
    ._EVAL_42(dcacheArb__EVAL_42),
    ._EVAL_43(dcacheArb__EVAL_43),
    ._EVAL_44(dcacheArb__EVAL_44),
    ._EVAL_45(dcacheArb__EVAL_45),
    ._EVAL_46(dcacheArb__EVAL_46),
    ._EVAL_47(dcacheArb__EVAL_47),
    ._EVAL_48(dcacheArb__EVAL_48),
    ._EVAL_49(dcacheArb__EVAL_49),
    ._EVAL_50(dcacheArb__EVAL_50),
    ._EVAL_51(dcacheArb__EVAL_51),
    ._EVAL_52(dcacheArb__EVAL_52),
    ._EVAL_53(dcacheArb__EVAL_53),
    ._EVAL_54(dcacheArb__EVAL_54),
    ._EVAL_55(dcacheArb__EVAL_55),
    ._EVAL_56(dcacheArb__EVAL_56),
    ._EVAL_57(dcacheArb__EVAL_57),
    ._EVAL_58(dcacheArb__EVAL_58),
    ._EVAL_59(dcacheArb__EVAL_59),
    ._EVAL_60(dcacheArb__EVAL_60),
    ._EVAL_61(dcacheArb__EVAL_61),
    ._EVAL_62(dcacheArb__EVAL_62),
    ._EVAL_63(dcacheArb__EVAL_63),
    ._EVAL_64(dcacheArb__EVAL_64),
    ._EVAL_65(dcacheArb__EVAL_65),
    ._EVAL_66(dcacheArb__EVAL_66),
    ._EVAL_67(dcacheArb__EVAL_67),
    ._EVAL_68(dcacheArb__EVAL_68),
    ._EVAL_69(dcacheArb__EVAL_69),
    ._EVAL_70(dcacheArb__EVAL_70),
    ._EVAL_71(dcacheArb__EVAL_71),
    ._EVAL_72(dcacheArb__EVAL_72),
    ._EVAL_73(dcacheArb__EVAL_73),
    ._EVAL_74(dcacheArb__EVAL_74),
    ._EVAL_75(dcacheArb__EVAL_75),
    ._EVAL_76(dcacheArb__EVAL_76),
    ._EVAL_77(dcacheArb__EVAL_77),
    ._EVAL_78(dcacheArb__EVAL_78),
    ._EVAL_79(dcacheArb__EVAL_79),
    ._EVAL_80(dcacheArb__EVAL_80),
    ._EVAL_81(dcacheArb__EVAL_81),
    ._EVAL_82(dcacheArb__EVAL_82),
    ._EVAL_83(dcacheArb__EVAL_83),
    ._EVAL_84(dcacheArb__EVAL_84),
    ._EVAL_85(dcacheArb__EVAL_85)
  );
  _EVAL_115 frontend (
    ._EVAL(frontend__EVAL),
    ._EVAL_0(frontend__EVAL_0),
    ._EVAL_1(frontend__EVAL_1),
    ._EVAL_2(frontend__EVAL_2),
    ._EVAL_3(frontend__EVAL_3),
    ._EVAL_4(frontend__EVAL_4),
    ._EVAL_5(frontend__EVAL_5),
    ._EVAL_6(frontend__EVAL_6),
    ._EVAL_7(frontend__EVAL_7),
    ._EVAL_8(frontend__EVAL_8),
    ._EVAL_9(frontend__EVAL_9),
    ._EVAL_10(frontend__EVAL_10),
    ._EVAL_11(frontend__EVAL_11),
    ._EVAL_12(frontend__EVAL_12),
    ._EVAL_13(frontend__EVAL_13),
    ._EVAL_14(frontend__EVAL_14),
    ._EVAL_15(frontend__EVAL_15),
    ._EVAL_16(frontend__EVAL_16),
    ._EVAL_17(frontend__EVAL_17),
    ._EVAL_18(frontend__EVAL_18),
    ._EVAL_19(frontend__EVAL_19),
    ._EVAL_20(frontend__EVAL_20),
    ._EVAL_21(frontend__EVAL_21),
    ._EVAL_22(frontend__EVAL_22),
    ._EVAL_23(frontend__EVAL_23),
    ._EVAL_24(frontend__EVAL_24),
    ._EVAL_25(frontend__EVAL_25),
    ._EVAL_26(frontend__EVAL_26),
    ._EVAL_27(frontend__EVAL_27),
    ._EVAL_28(frontend__EVAL_28),
    ._EVAL_29(frontend__EVAL_29),
    ._EVAL_30(frontend__EVAL_30),
    ._EVAL_31(frontend__EVAL_31),
    ._EVAL_32(frontend__EVAL_32),
    ._EVAL_33(frontend__EVAL_33),
    ._EVAL_34(frontend__EVAL_34),
    ._EVAL_35(frontend__EVAL_35),
    ._EVAL_36(frontend__EVAL_36),
    ._EVAL_37(frontend__EVAL_37),
    ._EVAL_38(frontend__EVAL_38),
    ._EVAL_39(frontend__EVAL_39),
    ._EVAL_40(frontend__EVAL_40),
    ._EVAL_41(frontend__EVAL_41),
    ._EVAL_42(frontend__EVAL_42),
    ._EVAL_43(frontend__EVAL_43),
    ._EVAL_44(frontend__EVAL_44),
    ._EVAL_45(frontend__EVAL_45),
    ._EVAL_46(frontend__EVAL_46),
    ._EVAL_47(frontend__EVAL_47),
    ._EVAL_48(frontend__EVAL_48),
    ._EVAL_49(frontend__EVAL_49),
    ._EVAL_50(frontend__EVAL_50),
    ._EVAL_51(frontend__EVAL_51),
    ._EVAL_52(frontend__EVAL_52),
    ._EVAL_53(frontend__EVAL_53),
    ._EVAL_54(frontend__EVAL_54),
    ._EVAL_55(frontend__EVAL_55),
    ._EVAL_56(frontend__EVAL_56),
    ._EVAL_57(frontend__EVAL_57),
    ._EVAL_58(frontend__EVAL_58),
    ._EVAL_59(frontend__EVAL_59),
    ._EVAL_60(frontend__EVAL_60),
    ._EVAL_61(frontend__EVAL_61),
    ._EVAL_62(frontend__EVAL_62),
    ._EVAL_63(frontend__EVAL_63),
    ._EVAL_64(frontend__EVAL_64),
    ._EVAL_65(frontend__EVAL_65),
    ._EVAL_66(frontend__EVAL_66),
    ._EVAL_67(frontend__EVAL_67),
    ._EVAL_68(frontend__EVAL_68),
    ._EVAL_69(frontend__EVAL_69),
    ._EVAL_70(frontend__EVAL_70),
    ._EVAL_71(frontend__EVAL_71),
    ._EVAL_72(frontend__EVAL_72),
    ._EVAL_73(frontend__EVAL_73),
    ._EVAL_74(frontend__EVAL_74),
    ._EVAL_75(frontend__EVAL_75),
    ._EVAL_76(frontend__EVAL_76),
    ._EVAL_77(frontend__EVAL_77),
    ._EVAL_78(frontend__EVAL_78),
    ._EVAL_79(frontend__EVAL_79),
    ._EVAL_80(frontend__EVAL_80),
    ._EVAL_81(frontend__EVAL_81),
    ._EVAL_82(frontend__EVAL_82),
    ._EVAL_83(frontend__EVAL_83),
    ._EVAL_84(frontend__EVAL_84),
    ._EVAL_85(frontend__EVAL_85),
    ._EVAL_86(frontend__EVAL_86),
    ._EVAL_87(frontend__EVAL_87),
    ._EVAL_88(frontend__EVAL_88),
    ._EVAL_89(frontend__EVAL_89),
    ._EVAL_90(frontend__EVAL_90),
    ._EVAL_91(frontend__EVAL_91),
    ._EVAL_92(frontend__EVAL_92),
    ._EVAL_93(frontend__EVAL_93),
    ._EVAL_94(frontend__EVAL_94),
    ._EVAL_95(frontend__EVAL_95),
    ._EVAL_96(frontend__EVAL_96),
    ._EVAL_97(frontend__EVAL_97),
    ._EVAL_98(frontend__EVAL_98),
    ._EVAL_99(frontend__EVAL_99),
    ._EVAL_100(frontend__EVAL_100),
    ._EVAL_101(frontend__EVAL_101),
    ._EVAL_102(frontend__EVAL_102),
    ._EVAL_103(frontend__EVAL_103),
    ._EVAL_104(frontend__EVAL_104),
    ._EVAL_105(frontend__EVAL_105),
    ._EVAL_106(frontend__EVAL_106),
    ._EVAL_107(frontend__EVAL_107),
    ._EVAL_108(frontend__EVAL_108),
    ._EVAL_109(frontend__EVAL_109),
    ._EVAL_110(frontend__EVAL_110),
    ._EVAL_111(frontend__EVAL_111),
    ._EVAL_112(frontend__EVAL_112),
    ._EVAL_113(frontend__EVAL_113),
    ._EVAL_114(frontend__EVAL_114),
    ._EVAL_115(frontend__EVAL_115),
    ._EVAL_116(frontend__EVAL_116),
    ._EVAL_117(frontend__EVAL_117),
    ._EVAL_118(frontend__EVAL_118),
    ._EVAL_119(frontend__EVAL_119),
    ._EVAL_120(frontend__EVAL_120)
  );
  _EVAL_104 tlSlaveXbar (
    ._EVAL(tlSlaveXbar__EVAL),
    ._EVAL_0(tlSlaveXbar__EVAL_0),
    ._EVAL_1(tlSlaveXbar__EVAL_1),
    ._EVAL_2(tlSlaveXbar__EVAL_2),
    ._EVAL_3(tlSlaveXbar__EVAL_3),
    ._EVAL_4(tlSlaveXbar__EVAL_4),
    ._EVAL_5(tlSlaveXbar__EVAL_5),
    ._EVAL_6(tlSlaveXbar__EVAL_6),
    ._EVAL_7(tlSlaveXbar__EVAL_7),
    ._EVAL_8(tlSlaveXbar__EVAL_8),
    ._EVAL_9(tlSlaveXbar__EVAL_9),
    ._EVAL_10(tlSlaveXbar__EVAL_10),
    ._EVAL_11(tlSlaveXbar__EVAL_11),
    ._EVAL_12(tlSlaveXbar__EVAL_12),
    ._EVAL_13(tlSlaveXbar__EVAL_13),
    ._EVAL_14(tlSlaveXbar__EVAL_14),
    ._EVAL_15(tlSlaveXbar__EVAL_15),
    ._EVAL_16(tlSlaveXbar__EVAL_16),
    ._EVAL_17(tlSlaveXbar__EVAL_17),
    ._EVAL_18(tlSlaveXbar__EVAL_18),
    ._EVAL_19(tlSlaveXbar__EVAL_19),
    ._EVAL_20(tlSlaveXbar__EVAL_20),
    ._EVAL_21(tlSlaveXbar__EVAL_21),
    ._EVAL_22(tlSlaveXbar__EVAL_22),
    ._EVAL_23(tlSlaveXbar__EVAL_23),
    ._EVAL_24(tlSlaveXbar__EVAL_24),
    ._EVAL_25(tlSlaveXbar__EVAL_25),
    ._EVAL_26(tlSlaveXbar__EVAL_26),
    ._EVAL_27(tlSlaveXbar__EVAL_27),
    ._EVAL_28(tlSlaveXbar__EVAL_28),
    ._EVAL_29(tlSlaveXbar__EVAL_29),
    ._EVAL_30(tlSlaveXbar__EVAL_30),
    ._EVAL_31(tlSlaveXbar__EVAL_31),
    ._EVAL_32(tlSlaveXbar__EVAL_32),
    ._EVAL_33(tlSlaveXbar__EVAL_33),
    ._EVAL_34(tlSlaveXbar__EVAL_34),
    ._EVAL_35(tlSlaveXbar__EVAL_35),
    ._EVAL_36(tlSlaveXbar__EVAL_36),
    ._EVAL_37(tlSlaveXbar__EVAL_37),
    ._EVAL_38(tlSlaveXbar__EVAL_38),
    ._EVAL_39(tlSlaveXbar__EVAL_39),
    ._EVAL_40(tlSlaveXbar__EVAL_40),
    ._EVAL_41(tlSlaveXbar__EVAL_41),
    ._EVAL_42(tlSlaveXbar__EVAL_42),
    ._EVAL_43(tlSlaveXbar__EVAL_43),
    ._EVAL_44(tlSlaveXbar__EVAL_44)
  );
  _EVAL_133 core (
    ._EVAL(core__EVAL),
    ._EVAL_0(core__EVAL_0),
    ._EVAL_1(core__EVAL_1),
    ._EVAL_2(core__EVAL_2),
    ._EVAL_3(core__EVAL_3),
    ._EVAL_4(core__EVAL_4),
    ._EVAL_5(core__EVAL_5),
    ._EVAL_6(core__EVAL_6),
    ._EVAL_7(core__EVAL_7),
    ._EVAL_8(core__EVAL_8),
    ._EVAL_9(core__EVAL_9),
    ._EVAL_10(core__EVAL_10),
    ._EVAL_11(core__EVAL_11),
    ._EVAL_12(core__EVAL_12),
    ._EVAL_13(core__EVAL_13),
    ._EVAL_14(core__EVAL_14),
    ._EVAL_15(core__EVAL_15),
    ._EVAL_16(core__EVAL_16),
    ._EVAL_17(core__EVAL_17),
    ._EVAL_18(core__EVAL_18),
    ._EVAL_19(core__EVAL_19),
    ._EVAL_20(core__EVAL_20),
    ._EVAL_21(core__EVAL_21),
    ._EVAL_22(core__EVAL_22),
    ._EVAL_23(core__EVAL_23),
    ._EVAL_24(core__EVAL_24),
    ._EVAL_25(core__EVAL_25),
    ._EVAL_26(core__EVAL_26),
    ._EVAL_27(core__EVAL_27),
    ._EVAL_28(core__EVAL_28),
    ._EVAL_29(core__EVAL_29),
    ._EVAL_30(core__EVAL_30),
    ._EVAL_31(core__EVAL_31),
    ._EVAL_32(core__EVAL_32),
    ._EVAL_33(core__EVAL_33),
    ._EVAL_34(core__EVAL_34),
    ._EVAL_35(core__EVAL_35),
    ._EVAL_36(core__EVAL_36),
    ._EVAL_37(core__EVAL_37),
    ._EVAL_38(core__EVAL_38),
    ._EVAL_39(core__EVAL_39),
    ._EVAL_40(core__EVAL_40),
    ._EVAL_41(core__EVAL_41),
    ._EVAL_42(core__EVAL_42),
    ._EVAL_43(core__EVAL_43),
    ._EVAL_44(core__EVAL_44),
    ._EVAL_45(core__EVAL_45),
    ._EVAL_46(core__EVAL_46),
    ._EVAL_47(core__EVAL_47),
    ._EVAL_48(core__EVAL_48),
    ._EVAL_49(core__EVAL_49),
    ._EVAL_50(core__EVAL_50),
    ._EVAL_51(core__EVAL_51),
    ._EVAL_52(core__EVAL_52),
    ._EVAL_53(core__EVAL_53),
    ._EVAL_54(core__EVAL_54),
    ._EVAL_55(core__EVAL_55),
    ._EVAL_56(core__EVAL_56),
    ._EVAL_57(core__EVAL_57),
    ._EVAL_58(core__EVAL_58),
    ._EVAL_59(core__EVAL_59),
    ._EVAL_60(core__EVAL_60),
    ._EVAL_61(core__EVAL_61),
    ._EVAL_62(core__EVAL_62),
    ._EVAL_63(core__EVAL_63),
    ._EVAL_64(core__EVAL_64),
    ._EVAL_65(core__EVAL_65),
    ._EVAL_66(core__EVAL_66),
    ._EVAL_67(core__EVAL_67),
    ._EVAL_68(core__EVAL_68),
    ._EVAL_69(core__EVAL_69),
    ._EVAL_70(core__EVAL_70),
    ._EVAL_71(core__EVAL_71),
    ._EVAL_72(core__EVAL_72),
    ._EVAL_73(core__EVAL_73),
    ._EVAL_74(core__EVAL_74),
    ._EVAL_75(core__EVAL_75),
    ._EVAL_76(core__EVAL_76),
    ._EVAL_77(core__EVAL_77),
    ._EVAL_78(core__EVAL_78),
    ._EVAL_79(core__EVAL_79),
    ._EVAL_80(core__EVAL_80),
    ._EVAL_81(core__EVAL_81),
    ._EVAL_82(core__EVAL_82),
    ._EVAL_83(core__EVAL_83),
    ._EVAL_84(core__EVAL_84),
    ._EVAL_85(core__EVAL_85),
    ._EVAL_86(core__EVAL_86),
    ._EVAL_87(core__EVAL_87),
    ._EVAL_88(core__EVAL_88),
    ._EVAL_89(core__EVAL_89),
    ._EVAL_90(core__EVAL_90),
    ._EVAL_91(core__EVAL_91),
    ._EVAL_92(core__EVAL_92),
    ._EVAL_93(core__EVAL_93),
    ._EVAL_94(core__EVAL_94),
    ._EVAL_95(core__EVAL_95),
    ._EVAL_96(core__EVAL_96),
    ._EVAL_97(core__EVAL_97),
    ._EVAL_98(core__EVAL_98),
    ._EVAL_99(core__EVAL_99),
    ._EVAL_100(core__EVAL_100),
    ._EVAL_101(core__EVAL_101),
    ._EVAL_102(core__EVAL_102),
    ._EVAL_103(core__EVAL_103),
    ._EVAL_104(core__EVAL_104),
    ._EVAL_105(core__EVAL_105),
    ._EVAL_106(core__EVAL_106),
    ._EVAL_107(core__EVAL_107),
    ._EVAL_108(core__EVAL_108),
    ._EVAL_109(core__EVAL_109),
    ._EVAL_110(core__EVAL_110),
    ._EVAL_111(core__EVAL_111),
    ._EVAL_112(core__EVAL_112),
    ._EVAL_113(core__EVAL_113),
    ._EVAL_114(core__EVAL_114),
    ._EVAL_115(core__EVAL_115),
    ._EVAL_116(core__EVAL_116),
    ._EVAL_117(core__EVAL_117),
    ._EVAL_118(core__EVAL_118),
    ._EVAL_119(core__EVAL_119),
    ._EVAL_120(core__EVAL_120),
    ._EVAL_121(core__EVAL_121),
    ._EVAL_122(core__EVAL_122),
    ._EVAL_123(core__EVAL_123),
    ._EVAL_124(core__EVAL_124),
    ._EVAL_125(core__EVAL_125),
    ._EVAL_126(core__EVAL_126),
    ._EVAL_127(core__EVAL_127),
    ._EVAL_128(core__EVAL_128),
    ._EVAL_129(core__EVAL_129),
    ._EVAL_130(core__EVAL_130),
    ._EVAL_131(core__EVAL_131),
    ._EVAL_132(core__EVAL_132),
    ._EVAL_133(core__EVAL_133),
    ._EVAL_134(core__EVAL_134),
    ._EVAL_135(core__EVAL_135),
    ._EVAL_136(core__EVAL_136),
    ._EVAL_137(core__EVAL_137),
    ._EVAL_138(core__EVAL_138),
    ._EVAL_139(core__EVAL_139),
    ._EVAL_140(core__EVAL_140),
    ._EVAL_141(core__EVAL_141),
    ._EVAL_142(core__EVAL_142),
    ._EVAL_143(core__EVAL_143),
    ._EVAL_144(core__EVAL_144),
    ._EVAL_145(core__EVAL_145),
    ._EVAL_146(core__EVAL_146),
    ._EVAL_147(core__EVAL_147),
    ._EVAL_148(core__EVAL_148),
    ._EVAL_149(core__EVAL_149),
    ._EVAL_150(core__EVAL_150),
    ._EVAL_151(core__EVAL_151),
    ._EVAL_152(core__EVAL_152),
    ._EVAL_153(core__EVAL_153),
    ._EVAL_154(core__EVAL_154),
    ._EVAL_155(core__EVAL_155),
    ._EVAL_156(core__EVAL_156),
    ._EVAL_157(core__EVAL_157),
    ._EVAL_158(core__EVAL_158),
    ._EVAL_159(core__EVAL_159),
    ._EVAL_160(core__EVAL_160),
    ._EVAL_161(core__EVAL_161)
  );
  _EVAL_117 fragmenter (
    ._EVAL(fragmenter__EVAL),
    ._EVAL_0(fragmenter__EVAL_0),
    ._EVAL_1(fragmenter__EVAL_1),
    ._EVAL_2(fragmenter__EVAL_2),
    ._EVAL_3(fragmenter__EVAL_3),
    ._EVAL_4(fragmenter__EVAL_4),
    ._EVAL_5(fragmenter__EVAL_5),
    ._EVAL_6(fragmenter__EVAL_6),
    ._EVAL_7(fragmenter__EVAL_7),
    ._EVAL_8(fragmenter__EVAL_8),
    ._EVAL_9(fragmenter__EVAL_9),
    ._EVAL_10(fragmenter__EVAL_10),
    ._EVAL_11(fragmenter__EVAL_11),
    ._EVAL_12(fragmenter__EVAL_12),
    ._EVAL_13(fragmenter__EVAL_13),
    ._EVAL_14(fragmenter__EVAL_14),
    ._EVAL_15(fragmenter__EVAL_15),
    ._EVAL_16(fragmenter__EVAL_16),
    ._EVAL_17(fragmenter__EVAL_17),
    ._EVAL_18(fragmenter__EVAL_18),
    ._EVAL_19(fragmenter__EVAL_19),
    ._EVAL_20(fragmenter__EVAL_20),
    ._EVAL_21(fragmenter__EVAL_21),
    ._EVAL_22(fragmenter__EVAL_22),
    ._EVAL_23(fragmenter__EVAL_23),
    ._EVAL_24(fragmenter__EVAL_24),
    ._EVAL_25(fragmenter__EVAL_25),
    ._EVAL_26(fragmenter__EVAL_26),
    ._EVAL_27(fragmenter__EVAL_27),
    ._EVAL_28(fragmenter__EVAL_28)
  );
  assign ptw__EVAL_21 = core__EVAL_145;
  assign tlSlaveXbar__EVAL_8 = _EVAL_56;
  assign core__EVAL_57 = dcacheArb__EVAL_38;
  assign frontend__EVAL_80 = ptw__EVAL_151;
  assign _EVAL_55 = tlSlaveXbar__EVAL_22;
  assign fragmenter_1__EVAL_21 = dtim_adapter__EVAL_12;
  assign fragmenter__EVAL_13 = frontend__EVAL_20;
  assign tlSlaveXbar__EVAL_30 = fragmenter__EVAL_11;
  assign core__EVAL_53 = _EVAL_27;
  assign _EVAL_69 = _EVAL_82;
  assign dtim_adapter__EVAL_1 = fragmenter_1__EVAL_8;
  assign ptw__EVAL_60 = core__EVAL_37;
  assign core__EVAL_2 = dcacheArb__EVAL_70;
  assign dcache__EVAL_77 = dcacheArb__EVAL_25;
  assign dcache__EVAL_96 = ptw__EVAL_93;
  assign dcache__EVAL_126 = ptw__EVAL_32;
  assign frontend__EVAL_92 = fragmenter__EVAL_15;
  assign core__EVAL_154 = _EVAL_57;
  assign ptw__EVAL_186 = core__EVAL_78;
  assign core__EVAL_4 = dcacheArb__EVAL_53;
  assign frontend__EVAL_108 = ptw__EVAL_39;
  assign fragmenter__EVAL_5 = tlSlaveXbar__EVAL_7;
  assign dcacheArb__EVAL_75 = dtim_adapter__EVAL_7;
  assign ptw__EVAL_67 = core__EVAL_88;
  assign ptw__EVAL_3 = core__EVAL_36;
  assign frontend__EVAL_41 = ptw__EVAL_38;
  assign dcache__EVAL_15 = dcacheArb__EVAL_8;
  assign frontend__EVAL_32 = fragmenter__EVAL_20;
  assign frontend__EVAL_118 = core__EVAL_61;
  assign frontend__EVAL_69 = _EVAL_88;
  assign core__EVAL_18 = frontend__EVAL_6;
  assign frontend__EVAL_44 = ptw__EVAL_157;
  assign ptw__EVAL_56 = core__EVAL_98;
  assign ptw__EVAL_47 = core__EVAL_124;
  assign dcache__EVAL_67 = ptw__EVAL_182;
  assign _EVAL_80 = _EVAL_83[3:0];
  assign tlMasterXbar__EVAL_33 = _EVAL_14;
  assign frontend__EVAL_115 = ptw__EVAL_112;
  assign tlMasterXbar__EVAL_54 = _EVAL_53;
  assign dcacheArb__EVAL_10 = core__EVAL_139;
  assign dcache__EVAL_7 = ptw__EVAL_81;
  assign core__EVAL_140 = dcacheArb__EVAL_35;
  assign ptw__EVAL_41 = core__EVAL_95;
  assign tlMasterXbar__EVAL_6 = dcache__EVAL_127;
  assign frontend__EVAL_38 = ptw__EVAL_159;
  assign tlMasterXbar__EVAL_50 = frontend__EVAL_99;
  assign core__EVAL_71 = frontend__EVAL_58;
  assign dtim_adapter__EVAL_10 = dcacheArb__EVAL_56;
  assign _EVAL_39 = tlSlaveXbar__EVAL_5;
  assign core__EVAL_105 = frontend__EVAL_68;
  assign dcache__EVAL_36 = dcacheArb__EVAL_57;
  assign ptw__EVAL_87 = core__EVAL_66;
  assign tlSlaveXbar__EVAL_37 = _EVAL_51;
  assign ptw__EVAL_19 = core__EVAL_138;
  assign _EVAL_11 = tlSlaveXbar__EVAL_13;
  assign fragmenter__EVAL_18 = tlSlaveXbar__EVAL_32;
  assign frontend__EVAL_28 = ptw__EVAL_78;
  assign frontend__EVAL_75 = ptw__EVAL_96;
  assign frontend__EVAL_117 = ptw__EVAL_16;
  assign dcache__EVAL_80 = ptw__EVAL_53;
  assign _EVAL_0 = tlMasterXbar__EVAL_53;
  assign ptw__EVAL_129 = core__EVAL_38;
  assign dcacheArb__EVAL_40 = _EVAL_37;
  assign dcache__EVAL_103 = ptw__EVAL_80;
  assign core__EVAL_106 = dcacheArb__EVAL_11;
  assign dtim_adapter__EVAL_13 = dcacheArb__EVAL_22;
  assign dcache__EVAL_91 = ptw__EVAL_106;
  assign dtim_adapter__EVAL_15 = fragmenter_1__EVAL_26;
  assign frontend__EVAL_76 = ptw__EVAL_77;
  assign ptw__EVAL_156 = core__EVAL_27;
  assign tlSlaveXbar__EVAL_39 = _EVAL_65;
  assign core__EVAL_118 = dcacheArb__EVAL_63;
  assign _EVAL_46 = tlMasterXbar__EVAL_24;
  assign core__EVAL_90 = _EVAL_67;
  assign frontend__EVAL_50 = ptw__EVAL_127;
  assign fragmenter_1__EVAL_14 = dtim_adapter__EVAL_19;
  assign dcacheArb__EVAL_6 = dcache__EVAL_119;
  assign fragmenter__EVAL_3 = frontend__EVAL_105;
  assign dcache__EVAL_62 = ptw__EVAL_28;
  assign frontend__EVAL_83 = core__EVAL_79;
  assign frontend__EVAL_23 = core__EVAL_112;
  assign core__EVAL_12 = _EVAL_41;
  assign core__EVAL_81 = dcacheArb__EVAL_62;
  assign ptw__EVAL_140 = core__EVAL_25;
  assign tlMasterXbar__EVAL_34 = _EVAL_29;
  assign dcache__EVAL_111 = dcacheArb__EVAL_52;
  assign dcacheArb__EVAL_80 = core__EVAL_153;
  assign fragmenter__EVAL_28 = frontend__EVAL_101;
  assign _EVAL_95 = ~_EVAL_85;
  assign frontend__EVAL_33 = ptw__EVAL_130;
  assign _EVAL_72 = _EVAL_71 & core__EVAL_19;
  assign dcache__EVAL_110 = ptw__EVAL_117;
  assign ptw__EVAL_66 = core__EVAL_21;
  assign frontend__EVAL_72 = tlMasterXbar__EVAL_5;
  assign _EVAL_4 = tlMasterXbar__EVAL_16;
  assign _EVAL_35 = tlMasterXbar__EVAL_47;
  assign frontend__EVAL_93 = ptw__EVAL_13;
  assign ptw__EVAL_92 = core__EVAL_89;
  assign tlSlaveXbar__EVAL_18 = fragmenter_1__EVAL_25;
  assign fragmenter_1__EVAL_6 = tlSlaveXbar__EVAL_14;
  assign frontend__EVAL_0 = ptw__EVAL_134;
  assign frontend__EVAL_42 = ptw__EVAL_84;
  assign frontend__EVAL_85 = ptw__EVAL_128;
  assign dcache__EVAL_32 = dcacheArb__EVAL_82;
  assign core__EVAL_44 = _EVAL_69;
  assign frontend__EVAL_114 = ptw__EVAL_73;
  assign fragmenter__EVAL_7 = tlSlaveXbar__EVAL_33;
  assign ptw__EVAL_90 = core__EVAL_75;
  assign core__EVAL_119 = frontend__EVAL_56;
  assign _EVAL_16 = _EVAL_91 >= 4'h8;
  assign ptw__EVAL_104 = core__EVAL_87;
  assign core__EVAL_160 = dcacheArb__EVAL_50;
  assign dcacheArb__EVAL_13 = dcache__EVAL_83;
  assign dcacheArb__EVAL_18 = dcache__EVAL_3;
  assign fragmenter__EVAL_23 = tlSlaveXbar__EVAL_35;
  assign tlMasterXbar__EVAL_52 = dcache__EVAL_9;
  assign _EVAL_78 = _EVAL_74;
  assign core__EVAL_135 = _EVAL_17;
  assign dcacheArb__EVAL_66 = dcache__EVAL_50;
  assign ptw__EVAL_48 = core__EVAL_30;
  assign _EVAL_10 = tlMasterXbar__EVAL_43;
  assign tlMasterXbar__EVAL_10 = dcache__EVAL_79;
  assign dcache__EVAL_35 = tlMasterXbar__EVAL_35;
  assign frontend__EVAL_66 = ptw__EVAL_51;
  assign dcache__EVAL_51 = tlMasterXbar__EVAL_27;
  assign dcache__EVAL_23 = ptw__EVAL_158;
  assign frontend__EVAL_36 = ptw__EVAL_160;
  assign fragmenter_1__EVAL_28 = tlSlaveXbar__EVAL_41;
  assign frontend__EVAL_61 = fragmenter__EVAL_21;
  assign dcacheArb__EVAL_17 = dcache__EVAL_11;
  assign dtim_adapter__EVAL_5 = _EVAL_37;
  assign ptw__EVAL_178 = core__EVAL_49;
  assign dcache__EVAL_63 = ptw__EVAL_57;
  assign tlSlaveXbar__EVAL_10 = fragmenter__EVAL_22;
  assign dcacheArb__EVAL_1 = core__EVAL_127;
  assign frontend__EVAL_96 = ptw__EVAL_141;
  assign dcache__EVAL_59 = ptw__EVAL_5;
  assign ptw__EVAL_43 = core__EVAL_58;
  assign frontend__EVAL_45 = core__EVAL_129;
  assign frontend__EVAL_119 = ptw__EVAL_83;
  assign dcacheArb__EVAL_27 = core__EVAL_51;
  assign _EVAL_18 = tlMasterXbar__EVAL_36;
  assign dcache__EVAL_82 = tlMasterXbar__EVAL_26;
  assign frontend__EVAL_57 = ptw__EVAL_145;
  assign tlMasterXbar__EVAL_0 = dcache__EVAL_18;
  assign core__EVAL_100 = _EVAL_78;
  assign ptw__EVAL_181 = core__EVAL_143;
  assign core__EVAL_116 = dcacheArb__EVAL_15;
  assign core__EVAL_141 = dcacheArb__EVAL_12;
  assign dcache__EVAL = ptw__EVAL_37;
  assign _EVAL_71 = _EVAL_76 & _EVAL_94;
  assign tlSlaveXbar__EVAL_15 = fragmenter_1__EVAL_4;
  assign fragmenter__EVAL_27 = frontend__EVAL_86;
  assign frontend__EVAL_49 = ptw__EVAL_171;
  assign ptw__EVAL_114 = core__EVAL;
  assign frontend__EVAL_77 = _EVAL_54;
  assign fragmenter_1__EVAL_22 = tlSlaveXbar__EVAL_40;
  assign tlSlaveXbar__EVAL_2 = fragmenter__EVAL_10;
  assign ptw__EVAL_71 = core__EVAL_20;
  assign _EVAL_24 = tlMasterXbar__EVAL_8;
  assign dtim_adapter__EVAL_20 = fragmenter_1__EVAL_16;
  assign dcacheArb__EVAL_83 = dcache__EVAL_28;
  assign frontend__EVAL_79 = ptw__EVAL_152;
  assign core__EVAL_48 = frontend__EVAL_73;
  assign ptw__EVAL_11 = core__EVAL_34;
  assign dtim_adapter__EVAL_16 = _EVAL_54;
  assign tlMasterXbar__EVAL_55 = _EVAL_60;
  assign dcacheArb__EVAL_60 = dtim_adapter__EVAL_25;
  assign tlMasterXbar__EVAL_4 = dcache__EVAL_38;
  assign fragmenter__EVAL_1 = tlSlaveXbar__EVAL_4;
  assign _EVAL_47 = tlSlaveXbar__EVAL_42;
  assign dcache__EVAL_39 = ptw__EVAL_147;
  assign _EVAL_81 = _EVAL_96;
  assign tlSlaveXbar__EVAL_12 = _EVAL_66;
  assign frontend__EVAL_90 = ptw__EVAL_20;
  assign _EVAL_48 = tlMasterXbar__EVAL_22;
  assign dcache__EVAL_14 = ptw__EVAL_132;
  assign frontend__EVAL_91 = ptw__EVAL_164;
  assign frontend__EVAL_26 = core__EVAL_110;
  assign frontend__EVAL_120 = ptw__EVAL_99;
  assign core__EVAL_45 = frontend__EVAL_10;
  assign ptw__EVAL_35 = _EVAL_54;
  assign frontend__EVAL_64 = core__EVAL_97;
  assign core__EVAL_46 = dcacheArb__EVAL_47;
  assign frontend__EVAL_24 = ptw__EVAL_74;
  assign ptw__EVAL_100 = core__EVAL_26;
  assign _EVAL_73 = _EVAL_72 & _EVAL_95;
  assign dtim_adapter__EVAL_26 = fragmenter_1__EVAL;
  assign dcache__EVAL_55 = ptw__EVAL_139;
  assign core__EVAL_63 = _EVAL_28;
  assign frontend__EVAL_113 = core__EVAL_121;
  assign dcache__EVAL_75 = ptw__EVAL_79;
  assign dcache__EVAL_112 = _EVAL_37;
  assign tlMasterXbar__EVAL_31 = dcache__EVAL_13;
  assign fragmenter__EVAL_6 = _EVAL_54;
  assign dtim_adapter__EVAL_9 = fragmenter_1__EVAL_1;
  assign core__EVAL_82 = _EVAL_64;
  assign frontend__EVAL_104 = core__EVAL_130;
  assign dcache__EVAL_122 = dcacheArb__EVAL_48;
  assign ptw__EVAL_55 = core__EVAL_41;
  assign dcache__EVAL_125 = ptw__EVAL_183;
  assign tlMasterXbar__EVAL_19 = _EVAL_61;
  assign frontend__EVAL_71 = ptw__EVAL_168;
  assign dcacheArb__EVAL_49 = dcache__EVAL_2;
  assign frontend__EVAL_11 = ptw__EVAL_155;
  assign frontend__EVAL_81 = ptw__EVAL_31;
  assign ptw__EVAL_119 = core__EVAL_93;
  assign dcache__EVAL_49 = ptw__EVAL_24;
  assign tlSlaveXbar__EVAL_19 = fragmenter__EVAL_0;
  assign dcacheArb__EVAL_46 = dcache__EVAL_124;
  assign ptw__EVAL_166 = core__EVAL_159;
  assign dcache__EVAL_84 = ptw__EVAL_52;
  assign frontend__EVAL_30 = ptw__EVAL_64;
  assign ptw__EVAL_122 = core__EVAL_142;
  assign core__EVAL_126 = dcacheArb__EVAL_45;
  assign tlMasterXbar__EVAL_15 = _EVAL_37;
  assign tlMasterXbar__EVAL_28 = dcache__EVAL_72;
  assign tlMasterXbar__EVAL_25 = _EVAL_19;
  assign dcache__EVAL_16 = dcacheArb__EVAL_2;
  assign dcacheArb__EVAL_85 = dtim_adapter__EVAL_23;
  assign core__EVAL_72 = frontend__EVAL_14;
  assign dcache__EVAL_47 = ptw__EVAL_161;
  assign dcache__EVAL_98 = dcacheArb__EVAL_37;
  assign fragmenter_1__EVAL_20 = dtim_adapter__EVAL_18;
  assign dcache__EVAL_52 = dcacheArb__EVAL_23;
  assign tlMasterXbar__EVAL_48 = frontend__EVAL_62;
  assign ptw__EVAL_85 = core__EVAL_13;
  assign core__EVAL_158 = 1'h0;
  assign frontend__EVAL_51 = tlMasterXbar__EVAL_23;
  assign _EVAL_63 = tlMasterXbar__EVAL_46;
  assign dcache__EVAL_45 = dcacheArb__EVAL_24;
  assign dcache__EVAL_40 = ptw__EVAL_15;
  assign fragmenter_1__EVAL_27 = tlSlaveXbar__EVAL_0;
  assign ptw__EVAL_142 = core__EVAL_86;
  assign core__EVAL_47 = frontend__EVAL_27;
  assign dcache__EVAL_121 = ptw__EVAL_124;
  assign fragmenter_1__EVAL_7 = tlSlaveXbar__EVAL_28;
  assign tlMasterXbar__EVAL_18 = dcache__EVAL_20;
  assign tlSlaveXbar__EVAL_3 = _EVAL_54;
  assign frontend__EVAL_1 = ptw__EVAL_33;
  assign frontend__EVAL_22 = ptw__EVAL_25;
  assign dcache__EVAL_85 = ptw__EVAL_103;
  assign dcache__EVAL_93 = _EVAL_54;
  assign ptw__EVAL_70 = core__EVAL_17;
  assign dcache__EVAL_78 = ptw__EVAL_2;
  assign frontend__EVAL_17 = ptw__EVAL_116;
  assign dcache__EVAL_60 = ptw__EVAL_165;
  assign dcacheArb__EVAL_21 = dcache__EVAL_31;
  assign dcache__EVAL_30 = ptw__EVAL_91;
  assign dcacheArb__EVAL_16 = dcache__EVAL_54;
  assign _EVAL = tlMasterXbar__EVAL_1;
  assign frontend__EVAL_13 = ptw__EVAL_153;
  assign _EVAL_45 = tlMasterXbar__EVAL_56;
  assign frontend__EVAL_65 = core__EVAL_5;
  assign core__EVAL_84 = _EVAL_7;
  assign frontend__EVAL_109 = core__EVAL_29;
  assign dcache__EVAL_41 = ptw__EVAL_10;
  assign core__EVAL_23 = dcacheArb__EVAL_33;
  assign dcache__EVAL_118 = tlMasterXbar__EVAL_13;
  assign dcacheArb__EVAL_55 = core__EVAL_16;
  assign frontend__EVAL_100 = _EVAL_37;
  assign core__EVAL_122 = _EVAL_43;
  assign dcacheArb__EVAL_79 = dtim_adapter__EVAL_11;
  assign fragmenter__EVAL_14 = tlSlaveXbar__EVAL_27;
  assign fragmenter__EVAL_12 = tlSlaveXbar__EVAL_24;
  assign core__EVAL_157 = _EVAL_81;
  assign frontend__EVAL_89 = ptw__EVAL_150;
  assign tlSlaveXbar__EVAL_38 = fragmenter_1__EVAL_2;
  assign _EVAL_52 = _EVAL_87;
  assign ptw__EVAL_185 = core__EVAL_120;
  assign frontend__EVAL_53 = ptw__EVAL_18;
  assign frontend__EVAL_5 = core__EVAL_15;
  assign dcache__EVAL_19 = _EVAL_57;
  assign core__EVAL_59 = frontend__EVAL_98;
  assign core__EVAL_109 = dcacheArb__EVAL_65;
  assign fragmenter__EVAL_9 = frontend__EVAL_84;
  assign tlSlaveXbar__EVAL_26 = fragmenter__EVAL_19;
  assign ptw__EVAL_6 = core__EVAL_114;
  assign dcacheArb__EVAL = dcache__EVAL_25;
  assign frontend__EVAL_95 = ptw__EVAL_123;
  assign _EVAL_12 = core__EVAL_99;
  assign dcacheArb__EVAL_74 = core__EVAL_146;
  assign frontend__EVAL_18 = core__EVAL_24;
  assign dcache__EVAL_43 = ptw__EVAL_176;
  assign dcacheArb__EVAL_67 = dtim_adapter__EVAL_0;
  assign tlSlaveXbar__EVAL_11 = _EVAL_58;
  assign dcache__EVAL_66 = ptw__EVAL_95;
  assign frontend__EVAL_9 = ptw__EVAL_126;
  assign dtim_adapter__EVAL_3 = dcacheArb__EVAL_7;
  assign dcache__EVAL_94 = tlMasterXbar__EVAL_44;
  assign dcacheArb__EVAL_29 = dcache__EVAL_128;
  assign ptw__EVAL_107 = core__EVAL_161;
  assign dcache__EVAL_108 = ptw__EVAL_154;
  assign _EVAL_97 = _EVAL_30;
  assign fragmenter_1__EVAL_3 = dtim_adapter__EVAL_22;
  assign core__EVAL_8 = _EVAL_68;
  assign tlSlaveXbar__EVAL_16 = _EVAL_23;
  assign frontend__EVAL_74 = tlMasterXbar__EVAL_17;
  assign fragmenter__EVAL_17 = tlSlaveXbar__EVAL_31;
  assign tlSlaveXbar__EVAL_29 = fragmenter__EVAL_24;
  assign ptw__EVAL_12 = core__EVAL_67;
  assign core__EVAL_92 = _EVAL_37;
  assign frontend__EVAL_102 = ptw__EVAL_163;
  assign dcacheArb__EVAL_26 = core__EVAL_68;
  assign _EVAL_44 = tlMasterXbar__EVAL_7;
  assign frontend__EVAL_31 = ptw__EVAL_75;
  assign dcacheArb__EVAL_68 = dcache__EVAL_69;
  assign dcacheArb__EVAL_34 = dcache__EVAL_107;
  assign core__EVAL_131 = _EVAL_50;
  assign dcacheArb__EVAL_32 = core__EVAL_76;
  assign dcache__EVAL_21 = ptw__EVAL_172;
  assign dcache__EVAL_58 = ptw__EVAL_44;
  assign dcache__EVAL_81 = ptw__EVAL_40;
  assign dcacheArb__EVAL_58 = dcache__EVAL_33;
  assign tlSlaveXbar__EVAL_23 = _EVAL_37;
  assign tlMasterXbar__EVAL_29 = dcache__EVAL_56;
  assign core__EVAL_149 = frontend__EVAL_112;
  assign ptw__EVAL_26 = core__EVAL_102;
  assign dcache__EVAL_46 = ptw__EVAL_68;
  assign ptw__EVAL_101 = core__EVAL_136;
  assign core__EVAL_1 = dcacheArb__EVAL_28;
  assign dcache__EVAL_48 = ptw__EVAL_98;
  assign dcache__EVAL_22 = ptw__EVAL_118;
  assign dcacheArb__EVAL_36 = dcache__EVAL_24;
  assign dcache__EVAL_87 = tlMasterXbar__EVAL_12;
  assign frontend__EVAL_43 = core__EVAL_60;
  assign dcache__EVAL_105 = ptw__EVAL_42;
  assign tlMasterXbar__EVAL_38 = dcache__EVAL_26;
  assign frontend__EVAL_29 = core__EVAL_128;
  assign frontend__EVAL_97 = tlMasterXbar__EVAL_45;
  assign dcacheArb__EVAL_44 = core__EVAL_9;
  assign core__EVAL_43 = dcacheArb__EVAL_3;
  assign frontend__EVAL_40 = core__EVAL_148;
  assign frontend__EVAL = tlMasterXbar__EVAL_42;
  assign dcacheArb__EVAL_72 = dcache__EVAL_86;
  assign fragmenter_1__EVAL_12 = tlSlaveXbar__EVAL_43;
  assign dcache__EVAL_10 = ptw__EVAL_59;
  assign tlMasterXbar__EVAL_21 = _EVAL_54;
  assign _EVAL_94 = ~frontend__EVAL_39;
  assign ptw__EVAL_7 = core__EVAL_14;
  assign ptw__EVAL_45 = core__EVAL_94;
  assign dcache__EVAL_104 = ptw__EVAL_30;
  assign tlMasterXbar__EVAL_14 = _EVAL_15;
  assign core__EVAL_103 = _EVAL_21;
  assign _EVAL_3 = tlMasterXbar__EVAL_3;
  assign dcacheArb__EVAL_64 = core__EVAL_123;
  assign dcache__EVAL_113 = tlMasterXbar__EVAL_51;
  assign ptw__EVAL_120 = core__EVAL_125;
  assign dcache__EVAL_90 = ptw__EVAL_8;
  assign core__EVAL_152 = dcacheArb__EVAL_84;
  assign core__EVAL_115 = _EVAL_13;
  assign dcache__EVAL_73 = ptw__EVAL_14;
  assign ptw__EVAL_54 = core__EVAL_11;
  assign _EVAL_6 = tlSlaveXbar__EVAL;
  assign dcache__EVAL_120 = ptw__EVAL_4;
  assign frontend__EVAL_35 = ptw__EVAL_0;
  assign dtim_adapter__EVAL_2 = dcacheArb__EVAL_42;
  assign core__EVAL_117 = _EVAL_42;
  assign dcacheArb__EVAL_81 = dtim_adapter__EVAL_14;
  assign core__EVAL_150 = dcacheArb__EVAL_59;
  assign dcacheArb__EVAL_41 = dcache__EVAL_27;
  assign dcacheArb__EVAL_76 = dcache__EVAL_102;
  assign frontend__EVAL_63 = ptw__EVAL_162;
  assign frontend__EVAL_3 = fragmenter__EVAL_8;
  assign ptw__EVAL_34 = core__EVAL_35;
  assign core__EVAL_22 = frontend__EVAL_7;
  assign core__EVAL_107 = frontend__EVAL_48;
  assign ptw__EVAL_170 = core__EVAL_96;
  assign core__EVAL_80 = _EVAL_25;
  assign core__EVAL_0 = _EVAL_33;
  assign ptw__EVAL_82 = core__EVAL_155;
  assign core__EVAL_32 = dcacheArb__EVAL_9;
  assign ptw__EVAL_167 = core__EVAL_134;
  assign frontend__EVAL_15 = core__EVAL_65;
  assign ptw__EVAL_175 = core__EVAL_77;
  assign fragmenter_1__EVAL_0 = tlSlaveXbar__EVAL_36;
  assign tlMasterXbar__EVAL_2 = dcache__EVAL_95;
  assign core__EVAL_113 = _EVAL_75;
  assign ptw__EVAL_149 = core__EVAL_64;
  assign dcache__EVAL_92 = ptw__EVAL_63;
  assign frontend__EVAL_4 = ptw__EVAL_138;
  assign frontend__EVAL_25 = ptw__EVAL_146;
  assign _EVAL_38 = tlSlaveXbar__EVAL_20;
  assign tlSlaveXbar__EVAL_21 = _EVAL_31;
  assign ptw__EVAL_94 = core__EVAL_104;
  assign dcacheArb__EVAL_73 = dcache__EVAL_34;
  assign dcacheArb__EVAL_61 = core__EVAL_33;
  assign dcache__EVAL_71 = ptw__EVAL_97;
  assign core__EVAL_31 = _EVAL_40;
  assign dtim_adapter__EVAL = fragmenter_1__EVAL_19;
  assign _EVAL_76 = ~dcache__EVAL_102;
  assign _EVAL_86 = ~_EVAL_72;
  assign frontend__EVAL_60 = ptw__EVAL_173;
  assign dcache__EVAL_76 = ptw__EVAL_113;
  assign tlSlaveXbar__EVAL_6 = fragmenter_1__EVAL_30;
  assign frontend__EVAL_34 = ptw__EVAL_148;
  assign _EVAL_82 = _EVAL_2;
  assign dcacheArb__EVAL_20 = dcache__EVAL_70;
  assign ptw__EVAL_29 = core__EVAL_73;
  assign frontend__EVAL_54 = core__EVAL_52;
  assign frontend__EVAL_2 = fragmenter__EVAL_25;
  assign tlMasterXbar__EVAL_41 = _EVAL_8;
  assign dtim_adapter__EVAL_17 = fragmenter_1__EVAL_11;
  assign fragmenter__EVAL_4 = _EVAL_37;
  assign _EVAL_75 = _EVAL_93;
  assign frontend__EVAL_21 = ptw__EVAL_187;
  assign frontend__EVAL_106 = core__EVAL_101;
  assign dcache__EVAL_74 = ptw__EVAL_17;
  assign tlSlaveXbar__EVAL_34 = _EVAL_59;
  assign dcacheArb__EVAL_14 = dtim_adapter__EVAL_6;
  assign core__EVAL_42 = dcacheArb__EVAL_78;
  assign dcache__EVAL_1 = ptw__EVAL_62;
  assign dcacheArb__EVAL_43 = core__EVAL_56;
  assign fragmenter_1__EVAL_9 = dtim_adapter__EVAL_8;
  assign core__EVAL_83 = dcacheArb__EVAL_54;
  assign dcacheArb__EVAL_0 = dcache__EVAL_116;
  assign tlMasterXbar__EVAL = dcache__EVAL_106;
  assign dcache__EVAL_57 = ptw__EVAL_111;
  assign tlMasterXbar__EVAL_57 = frontend__EVAL_47;
  assign dcache__EVAL_123 = ptw__EVAL_136;
  assign dcacheArb__EVAL_39 = dcache__EVAL_100;
  assign dcache__EVAL_17 = ptw__EVAL_27;
  assign _EVAL_74 = _EVAL_22;
  assign tlMasterXbar__EVAL_37 = _EVAL_1;
  assign dcache__EVAL_61 = ptw__EVAL_121;
  assign _EVAL_85 = _EVAL_91 >= 4'h8;
  assign frontend__EVAL_12 = ptw__EVAL_174;
  assign dcache__EVAL_12 = ptw__EVAL_86;
  assign _EVAL_62 = tlMasterXbar__EVAL_9;
  assign tlMasterXbar__EVAL_49 = dcache__EVAL_4;
  assign dtim_adapter__EVAL_4 = fragmenter_1__EVAL_29;
  assign dtim_adapter__EVAL_21 = fragmenter_1__EVAL_13;
  assign frontend__EVAL_67 = ptw__EVAL_180;
  assign tlSlaveXbar__EVAL_17 = fragmenter_1__EVAL_24;
  assign tlMasterXbar__EVAL_40 = _EVAL_5;
  assign frontend__EVAL_116 = tlMasterXbar__EVAL_30;
  assign frontend__EVAL_8 = fragmenter__EVAL_2;
  assign frontend__EVAL_59 = ptw__EVAL_23;
  assign fragmenter_1__EVAL_15 = _EVAL_37;
  assign core__EVAL_74 = _EVAL_54;
  assign frontend__EVAL_88 = ptw__EVAL_76;
  assign core__EVAL_39 = dcacheArb__EVAL_77;
  assign dcache__EVAL_42 = tlMasterXbar__EVAL_32;
  assign frontend__EVAL_94 = fragmenter__EVAL_26;
  assign ptw__EVAL_49 = core__EVAL_70;
  assign fragmenter_1__EVAL_18 = dtim_adapter__EVAL_24;
  assign ptw__EVAL_102 = core__EVAL_50;
  assign dcache__EVAL_115 = dcacheArb__EVAL_19;
  assign frontend__EVAL_107 = ptw__EVAL_108;
  assign core__EVAL_3 = _EVAL_49;
  assign tlSlaveXbar__EVAL_25 = fragmenter_1__EVAL_17;
  assign ptw__EVAL_131 = core__EVAL_10;
  assign dcache__EVAL_68 = ptw__EVAL_133;
  assign frontend__EVAL_78 = ptw__EVAL_105;
  assign ptw__EVAL_109 = core__EVAL_55;
  assign core__EVAL_111 = _EVAL_32;
  assign frontend__EVAL_55 = ptw__EVAL_143;
  assign _EVAL_93 = _EVAL_34;
  assign core__EVAL_151 = _EVAL_9;
  assign core__EVAL_85 = dcacheArb__EVAL_71;
  assign dcache__EVAL_29 = ptw__EVAL_135;
  assign ptw__EVAL_50 = core__EVAL_133;
  assign dcacheArb__EVAL_31 = core__EVAL_144;
  assign dcache__EVAL_37 = ptw__EVAL_137;
  assign tlSlaveXbar__EVAL_44 = _EVAL_20;
  assign frontend__EVAL_52 = ptw__EVAL_110;
  assign tlMasterXbar__EVAL_39 = dcache__EVAL_53;
  assign _EVAL_88 = _EVAL_97;
  assign frontend__EVAL_70 = _EVAL_57;
  assign dcache__EVAL_0 = ptw__EVAL_9;
  assign dcache__EVAL_65 = ptw__EVAL_115;
  assign frontend__EVAL_46 = fragmenter__EVAL_16;
  assign core__EVAL_69 = dcacheArb__EVAL_5;
  assign ptw__EVAL_144 = core__EVAL_28;
  assign _EVAL_83 = _EVAL_91 + 4'h1;
  assign ptw__EVAL_184 = core__EVAL_108;
  assign ptw__EVAL_46 = core__EVAL_137;
  assign ptw__EVAL_72 = _EVAL_37;
  assign fragmenter__EVAL = frontend__EVAL_111;
  assign dcacheArb__EVAL_69 = dcache__EVAL_117;
  assign dcache__EVAL_6 = dcacheArb__EVAL_4;
  assign core__EVAL_147 = _EVAL_26;
  assign ptw__EVAL_169 = core__EVAL_6;
  assign frontend__EVAL_87 = ptw__EVAL_125;
  assign ptw__EVAL_61 = core__EVAL_54;
  assign fragmenter_1__EVAL_5 = tlSlaveXbar__EVAL_9;
  assign dcache__EVAL_8 = ptw__EVAL_69;
  assign frontend__EVAL_82 = ptw__EVAL_22;
  assign dcache__EVAL_44 = tlMasterXbar__EVAL_20;
  assign fragmenter_1__EVAL_23 = tlSlaveXbar__EVAL_1;
  assign frontend__EVAL_110 = ptw__EVAL_1;
  assign _EVAL_96 = _EVAL_36;
  assign dcache__EVAL_88 = dcacheArb__EVAL_51;
  assign dcache__EVAL_109 = ptw__EVAL_179;
  assign ptw__EVAL_65 = core__EVAL_156;
  assign dcacheArb__EVAL_30 = dcache__EVAL_99;
  assign fragmenter_1__EVAL_10 = _EVAL_54;
  assign ptw__EVAL_89 = core__EVAL_62;
  assign dcache__EVAL_97 = tlMasterXbar__EVAL_11;
  assign frontend__EVAL_16 = ptw__EVAL_177;
  assign frontend__EVAL_37 = ptw__EVAL;
  always @(posedge _EVAL_37) begin
    if (_EVAL_54) begin
      _EVAL_87 <= 1'h0;
    end else begin
      _EVAL_87 <= core__EVAL_7;
    end
    if (_EVAL_54) begin
      _EVAL_91 <= 4'h0;
    end else if (_EVAL_73) begin
      _EVAL_91 <= _EVAL_80;
    end else if (_EVAL_86) begin
      _EVAL_91 <= 4'h0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_87 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_91 = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
