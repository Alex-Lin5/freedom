//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_112(
  input  [1:0]  _EVAL,
  input         _EVAL_0,
  output        _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  output        _EVAL_6,
  output [31:0] _EVAL_7,
  output [1:0]  _EVAL_8,
  input  [7:0]  _EVAL_9,
  output [4:0]  _EVAL_10,
  output        _EVAL_11,
  output        _EVAL_12,
  input         _EVAL_13,
  output        _EVAL_14,
  input         _EVAL_15,
  output [31:0] _EVAL_16,
  output        _EVAL_17,
  input  [31:0] _EVAL_18,
  input         _EVAL_19,
  output [4:0]  _EVAL_20,
  input  [31:0] _EVAL_21,
  input  [4:0]  _EVAL_22,
  output [7:0]  _EVAL_23
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] _EVAL_24;
  reg  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  reg  _EVAL_32;
  reg [1:0] _EVAL_33;
  reg  _EVAL_34;
  reg [31:0] _EVAL_35;
  wire  _EVAL_36;
  reg  _EVAL_37;
  reg  _EVAL_38;
  reg  _EVAL_41;
  reg [31:0] _EVAL_42;
  reg  _EVAL_43;
  reg [31:0] _EVAL_44;
  reg [4:0] _EVAL_48;
  wire  _EVAL_49;
  reg [7:0] _EVAL_52;
  reg [4:0] _EVAL_53;
  wire  _EVAL_55;
  wire  _EVAL_56;
  reg [4:0] _EVAL_57;
  reg  _EVAL_58;
  reg  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  reg [7:0] _EVAL_66;
  wire  _EVAL_70;
  reg  _EVAL_71;
  reg [1:0] _EVAL_74;
  reg  _EVAL_75;
  reg  _EVAL_77;
  wire  _EVAL_78;
  reg [7:0] _EVAL_80;
  wire  _EVAL_81;
  reg  _EVAL_84;
  wire  _EVAL_85;
  reg  _EVAL_86;
  reg  _EVAL_88;
  reg  _EVAL_89;
  wire  _EVAL_90;
  reg  _EVAL_91;
  reg  _EVAL_92;
  wire  _EVAL_95;
  reg  _EVAL_96;
  wire [1:0] _EVAL_99;
  wire  _EVAL_100;
  reg [4:0] _EVAL_101;
  wire  _EVAL_102;
  reg  _EVAL_104;
  wire  _EVAL_106;
  reg [1:0] _EVAL_108;
  wire  _EVAL_109;
  reg [31:0] _EVAL_111;
  reg [31:0] _EVAL_112;
  reg [31:0] _EVAL_114;
  reg [31:0] _EVAL_115;
  reg [7:0] _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_122;
  wire  _EVAL_123;
  reg  _EVAL_124;
  reg  _EVAL_125;
  reg [31:0] _EVAL_127;
  reg  _EVAL_129;
  wire  _EVAL_130;
  reg  _EVAL_133;
  reg [7:0] _EVAL_134;
  reg  _EVAL_135;
  reg [4:0] _EVAL_136;
  reg [1:0] _EVAL_137;
  reg [1:0] _EVAL_138;
  reg [31:0] _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_142;
  wire  _EVAL_144;
  wire [2:0] _EVAL_146;
  assign _EVAL_146 = {_EVAL_37,_EVAL_75,_EVAL_88};
  assign _EVAL_14 = _EVAL_36 ? _EVAL_15 : _EVAL_25;
  assign _EVAL_119 = ~_EVAL_37;
  assign _EVAL_8 = _EVAL_36 ? _EVAL : _EVAL_33;
  assign _EVAL_90 = _EVAL_64 & _EVAL_36;
  assign _EVAL_56 = _EVAL_19 ? _EVAL_85 : _EVAL_90;
  assign _EVAL_10 = {_EVAL_146,_EVAL_99};
  assign _EVAL_81 = _EVAL_102 & _EVAL_109;
  assign _EVAL_142 = _EVAL_64 & _EVAL_59;
  assign _EVAL_12 = _EVAL_5 | _EVAL_96;
  assign _EVAL_95 = _EVAL_19 ? _EVAL_27 : _EVAL_26;
  assign _EVAL_11 = ~_EVAL_37;
  assign _EVAL_26 = _EVAL_142 & _EVAL_28;
  assign _EVAL_17 = _EVAL_36 ? _EVAL_3 : _EVAL_32;
  assign _EVAL_106 = _EVAL_64 & _EVAL_37;
  assign _EVAL_28 = ~_EVAL_88;
  assign _EVAL_144 = _EVAL_64 & _EVAL_96;
  assign _EVAL_60 = _EVAL_64 | _EVAL_96;
  assign _EVAL_55 = _EVAL_64 & _EVAL_75;
  assign _EVAL_16 = _EVAL_36 ? _EVAL_18 : _EVAL_112;
  assign _EVAL_27 = _EVAL_75 | _EVAL_102;
  assign _EVAL_6 = _EVAL_36 ? _EVAL_4 : _EVAL_41;
  assign _EVAL_64 = _EVAL_11 & _EVAL_5;
  assign _EVAL_140 = _EVAL_19 ? _EVAL_29 : _EVAL_61;
  assign _EVAL_123 = _EVAL_102 | _EVAL_75;
  assign _EVAL_78 = _EVAL_19 ? _EVAL_100 : _EVAL_81;
  assign _EVAL_122 = _EVAL_142 | _EVAL_88;
  assign _EVAL_100 = _EVAL_37 | _EVAL_55;
  assign _EVAL_99 = {_EVAL_59,_EVAL_96};
  assign _EVAL_65 = _EVAL_55 | _EVAL_37;
  assign _EVAL_36 = ~_EVAL_96;
  assign _EVAL_85 = _EVAL_59 | _EVAL_144;
  assign _EVAL_1 = _EVAL_36 ? _EVAL_13 : _EVAL_92;
  assign _EVAL_130 = _EVAL_55 & _EVAL_119;
  assign _EVAL_29 = _EVAL_88 | _EVAL_142;
  assign _EVAL_61 = _EVAL_144 & _EVAL_70;
  assign _EVAL_20 = _EVAL_36 ? _EVAL_22 : _EVAL_136;
  assign _EVAL_23 = _EVAL_36 ? _EVAL_9 : _EVAL_66;
  assign _EVAL_49 = _EVAL_19 ? _EVAL_106 : _EVAL_130;
  assign _EVAL_109 = ~_EVAL_75;
  assign _EVAL_63 = _EVAL_144 | _EVAL_59;
  assign _EVAL_102 = _EVAL_64 & _EVAL_88;
  assign _EVAL_70 = ~_EVAL_59;
  assign _EVAL_7 = _EVAL_36 ? _EVAL_21 : _EVAL_35;
  always @(posedge _EVAL_2) begin
    if (_EVAL_140) begin
      if (_EVAL_88) begin
        _EVAL_24 <= _EVAL_42;
      end else begin
        _EVAL_24 <= _EVAL_21;
      end
    end
    if (_EVAL_56) begin
      if (_EVAL_59) begin
        _EVAL_25 <= _EVAL_34;
      end else begin
        _EVAL_25 <= _EVAL_15;
      end
    end
    if (_EVAL_56) begin
      if (_EVAL_59) begin
        _EVAL_32 <= _EVAL_91;
      end else begin
        _EVAL_32 <= _EVAL_3;
      end
    end
    if (_EVAL_56) begin
      if (_EVAL_59) begin
        _EVAL_33 <= _EVAL_74;
      end else begin
        _EVAL_33 <= _EVAL;
      end
    end
    if (_EVAL_140) begin
      if (_EVAL_88) begin
        _EVAL_34 <= _EVAL_58;
      end else begin
        _EVAL_34 <= _EVAL_15;
      end
    end
    if (_EVAL_56) begin
      if (_EVAL_59) begin
        _EVAL_35 <= _EVAL_24;
      end else begin
        _EVAL_35 <= _EVAL_21;
      end
    end
    if (_EVAL_0) begin
      _EVAL_37 <= 1'h0;
    end else if (_EVAL_19) begin
      _EVAL_37 <= _EVAL_106;
    end else begin
      _EVAL_37 <= _EVAL_65;
    end
    if (_EVAL_49) begin
      _EVAL_38 <= _EVAL_13;
    end
    if (_EVAL_56) begin
      if (_EVAL_59) begin
        _EVAL_41 <= _EVAL_86;
      end else begin
        _EVAL_41 <= _EVAL_4;
      end
    end
    if (_EVAL_95) begin
      if (_EVAL_75) begin
        _EVAL_42 <= _EVAL_115;
      end else begin
        _EVAL_42 <= _EVAL_21;
      end
    end
    if (_EVAL_95) begin
      if (_EVAL_75) begin
        _EVAL_43 <= _EVAL_133;
      end else begin
        _EVAL_43 <= _EVAL_3;
      end
    end
    if (_EVAL_78) begin
      if (_EVAL_37) begin
        _EVAL_44 <= _EVAL_139;
      end else begin
        _EVAL_44 <= _EVAL_18;
      end
    end
    if (_EVAL_95) begin
      if (_EVAL_75) begin
        _EVAL_48 <= _EVAL_101;
      end else begin
        _EVAL_48 <= _EVAL_22;
      end
    end
    if (_EVAL_140) begin
      if (_EVAL_88) begin
        _EVAL_52 <= _EVAL_134;
      end else begin
        _EVAL_52 <= _EVAL_9;
      end
    end
    if (_EVAL_140) begin
      if (_EVAL_88) begin
        _EVAL_53 <= _EVAL_48;
      end else begin
        _EVAL_53 <= _EVAL_22;
      end
    end
    if (_EVAL_49) begin
      _EVAL_57 <= _EVAL_22;
    end
    if (_EVAL_95) begin
      if (_EVAL_75) begin
        _EVAL_58 <= _EVAL_89;
      end else begin
        _EVAL_58 <= _EVAL_15;
      end
    end
    if (_EVAL_0) begin
      _EVAL_59 <= 1'h0;
    end else if (_EVAL_19) begin
      _EVAL_59 <= _EVAL_29;
    end else begin
      _EVAL_59 <= _EVAL_63;
    end
    if (_EVAL_56) begin
      if (_EVAL_59) begin
        _EVAL_66 <= _EVAL_52;
      end else begin
        _EVAL_66 <= _EVAL_9;
      end
    end
    if (_EVAL_49) begin
      _EVAL_71 <= _EVAL_3;
    end
    if (_EVAL_140) begin
      if (_EVAL_88) begin
        _EVAL_74 <= _EVAL_108;
      end else begin
        _EVAL_74 <= _EVAL;
      end
    end
    if (_EVAL_0) begin
      _EVAL_75 <= 1'h0;
    end else if (_EVAL_19) begin
      _EVAL_75 <= _EVAL_100;
    end else begin
      _EVAL_75 <= _EVAL_123;
    end
    if (_EVAL_95) begin
      if (_EVAL_75) begin
        _EVAL_77 <= _EVAL_135;
      end else begin
        _EVAL_77 <= _EVAL_4;
      end
    end
    if (_EVAL_78) begin
      if (_EVAL_37) begin
        _EVAL_80 <= _EVAL_118;
      end else begin
        _EVAL_80 <= _EVAL_9;
      end
    end
    if (_EVAL_49) begin
      _EVAL_84 <= _EVAL_15;
    end
    if (_EVAL_140) begin
      if (_EVAL_88) begin
        _EVAL_86 <= _EVAL_77;
      end else begin
        _EVAL_86 <= _EVAL_4;
      end
    end
    if (_EVAL_0) begin
      _EVAL_88 <= 1'h0;
    end else if (_EVAL_19) begin
      _EVAL_88 <= _EVAL_27;
    end else begin
      _EVAL_88 <= _EVAL_122;
    end
    if (_EVAL_78) begin
      if (_EVAL_37) begin
        _EVAL_89 <= _EVAL_84;
      end else begin
        _EVAL_89 <= _EVAL_15;
      end
    end
    if (_EVAL_140) begin
      if (_EVAL_88) begin
        _EVAL_91 <= _EVAL_43;
      end else begin
        _EVAL_91 <= _EVAL_3;
      end
    end
    if (_EVAL_56) begin
      if (_EVAL_59) begin
        _EVAL_92 <= _EVAL_129;
      end else begin
        _EVAL_92 <= _EVAL_13;
      end
    end
    if (_EVAL_0) begin
      _EVAL_96 <= 1'h0;
    end else if (_EVAL_19) begin
      _EVAL_96 <= _EVAL_85;
    end else begin
      _EVAL_96 <= _EVAL_60;
    end
    if (_EVAL_78) begin
      if (_EVAL_37) begin
        _EVAL_101 <= _EVAL_57;
      end else begin
        _EVAL_101 <= _EVAL_22;
      end
    end
    if (_EVAL_78) begin
      if (_EVAL_37) begin
        _EVAL_104 <= _EVAL_38;
      end else begin
        _EVAL_104 <= _EVAL_13;
      end
    end
    if (_EVAL_95) begin
      if (_EVAL_75) begin
        _EVAL_108 <= _EVAL_138;
      end else begin
        _EVAL_108 <= _EVAL;
      end
    end
    if (_EVAL_95) begin
      if (_EVAL_75) begin
        _EVAL_111 <= _EVAL_44;
      end else begin
        _EVAL_111 <= _EVAL_18;
      end
    end
    if (_EVAL_56) begin
      if (_EVAL_59) begin
        _EVAL_112 <= _EVAL_114;
      end else begin
        _EVAL_112 <= _EVAL_18;
      end
    end
    if (_EVAL_140) begin
      if (_EVAL_88) begin
        _EVAL_114 <= _EVAL_111;
      end else begin
        _EVAL_114 <= _EVAL_18;
      end
    end
    if (_EVAL_78) begin
      if (_EVAL_37) begin
        _EVAL_115 <= _EVAL_127;
      end else begin
        _EVAL_115 <= _EVAL_21;
      end
    end
    if (_EVAL_49) begin
      _EVAL_118 <= _EVAL_9;
    end
    if (_EVAL_95) begin
      if (_EVAL_75) begin
        _EVAL_124 <= _EVAL_104;
      end else begin
        _EVAL_124 <= _EVAL_13;
      end
    end
    if (_EVAL_49) begin
      _EVAL_125 <= _EVAL_4;
    end
    if (_EVAL_49) begin
      _EVAL_127 <= _EVAL_21;
    end
    if (_EVAL_140) begin
      if (_EVAL_88) begin
        _EVAL_129 <= _EVAL_124;
      end else begin
        _EVAL_129 <= _EVAL_13;
      end
    end
    if (_EVAL_78) begin
      if (_EVAL_37) begin
        _EVAL_133 <= _EVAL_71;
      end else begin
        _EVAL_133 <= _EVAL_3;
      end
    end
    if (_EVAL_95) begin
      if (_EVAL_75) begin
        _EVAL_134 <= _EVAL_80;
      end else begin
        _EVAL_134 <= _EVAL_9;
      end
    end
    if (_EVAL_78) begin
      if (_EVAL_37) begin
        _EVAL_135 <= _EVAL_125;
      end else begin
        _EVAL_135 <= _EVAL_4;
      end
    end
    if (_EVAL_56) begin
      if (_EVAL_59) begin
        _EVAL_136 <= _EVAL_53;
      end else begin
        _EVAL_136 <= _EVAL_22;
      end
    end
    if (_EVAL_49) begin
      _EVAL_137 <= _EVAL;
    end
    if (_EVAL_78) begin
      if (_EVAL_37) begin
        _EVAL_138 <= _EVAL_137;
      end else begin
        _EVAL_138 <= _EVAL;
      end
    end
    if (_EVAL_49) begin
      _EVAL_139 <= _EVAL_18;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_24 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_25 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_32 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_33 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_34 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_35 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_37 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_38 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_41 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_42 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_43 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_44 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_48 = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_52 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_53 = _RAND_14[4:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_57 = _RAND_15[4:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_58 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _EVAL_59 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _EVAL_66 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  _EVAL_71 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  _EVAL_74 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  _EVAL_75 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  _EVAL_77 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  _EVAL_80 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  _EVAL_84 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  _EVAL_86 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  _EVAL_88 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  _EVAL_89 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  _EVAL_91 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  _EVAL_92 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  _EVAL_96 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  _EVAL_101 = _RAND_31[4:0];
  _RAND_32 = {1{`RANDOM}};
  _EVAL_104 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  _EVAL_108 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  _EVAL_111 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  _EVAL_112 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  _EVAL_114 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  _EVAL_115 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  _EVAL_118 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  _EVAL_124 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  _EVAL_125 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  _EVAL_127 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  _EVAL_129 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  _EVAL_133 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  _EVAL_134 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  _EVAL_135 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  _EVAL_136 = _RAND_46[4:0];
  _RAND_47 = {1{`RANDOM}};
  _EVAL_137 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  _EVAL_138 = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  _EVAL_139 = _RAND_49[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
