//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_11(
  input  [3:0]  _EVAL,
  input  [31:0] _EVAL_0,
  output [1:0]  _EVAL_1,
  output        _EVAL_2,
  input  [1:0]  _EVAL_3,
  input         _EVAL_4,
  output        _EVAL_5,
  output [2:0]  _EVAL_6,
  input  [3:0]  _EVAL_7,
  output [3:0]  _EVAL_8,
  input  [3:0]  _EVAL_9,
  output [3:0]  _EVAL_10,
  input         _EVAL_11,
  output [2:0]  _EVAL_12,
  input         _EVAL_13,
  output [3:0]  _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  output        _EVAL_17,
  input         _EVAL_18,
  input  [3:0]  _EVAL_19,
  output        _EVAL_20,
  output        _EVAL_21,
  output [3:0]  _EVAL_22,
  input         _EVAL_23,
  output        _EVAL_24,
  input  [2:0]  _EVAL_25,
  input         _EVAL_26,
  output [3:0]  _EVAL_27,
  input  [31:0] _EVAL_28,
  output [2:0]  _EVAL_29,
  output [31:0] _EVAL_30,
  input         _EVAL_31,
  output [1:0]  _EVAL_32,
  input  [31:0] _EVAL_33,
  output        _EVAL_34,
  input  [3:0]  _EVAL_35,
  input         _EVAL_36,
  input         _EVAL_37,
  output        _EVAL_38,
  input         _EVAL_39,
  input  [3:0]  _EVAL_40,
  input         _EVAL_41,
  input  [2:0]  _EVAL_42,
  output [31:0] _EVAL_43,
  output [3:0]  _EVAL_44,
  output        _EVAL_45,
  output [31:0] _EVAL_46,
  input  [1:0]  _EVAL_47,
  input  [2:0]  _EVAL_48,
  output [3:0]  _EVAL_49,
  input         _EVAL_50,
  input  [3:0]  _EVAL_51,
  output [2:0]  _EVAL_52,
  input  [3:0]  _EVAL_53,
  input         _EVAL_54,
  input  [2:0]  _EVAL_55,
  output        _EVAL_56,
  output [1:0]  _EVAL_57,
  output        _EVAL_58,
  input         _EVAL_59,
  input         _EVAL_60,
  input  [2:0]  _EVAL_61,
  output [1:0]  _EVAL_62,
  input         _EVAL_63,
  output [31:0] _EVAL_64,
  input         _EVAL_65,
  input  [1:0]  _EVAL_66,
  output        _EVAL_67,
  output        _EVAL_68,
  output        _EVAL_69,
  output        _EVAL_70,
  input  [31:0] _EVAL_71,
  input  [31:0] _EVAL_72
);
  wire  bundleOut_0_a_sink__EVAL;
  wire  bundleOut_0_a_sink__EVAL_0;
  wire  bundleOut_0_a_sink__EVAL_1;
  wire [3:0] bundleOut_0_a_sink__EVAL_2;
  wire [31:0] bundleOut_0_a_sink__EVAL_3;
  wire  bundleOut_0_a_sink__EVAL_4;
  wire [3:0] bundleOut_0_a_sink__EVAL_5;
  wire  bundleOut_0_a_sink__EVAL_6;
  wire [2:0] bundleOut_0_a_sink__EVAL_7;
  wire  bundleOut_0_a_sink__EVAL_8;
  wire  bundleOut_0_a_sink__EVAL_9;
  wire [3:0] bundleOut_0_a_sink__EVAL_10;
  wire  bundleOut_0_a_sink__EVAL_11;
  wire [2:0] bundleOut_0_a_sink__EVAL_12;
  wire  bundleOut_0_a_sink__EVAL_13;
  wire [31:0] bundleOut_0_a_sink__EVAL_14;
  wire [3:0] bundleOut_0_a_sink__EVAL_15;
  wire [2:0] bundleOut_0_a_sink__EVAL_16;
  wire  bundleOut_0_a_sink__EVAL_17;
  wire  bundleOut_0_a_sink__EVAL_18;
  wire  bundleOut_0_a_sink__EVAL_19;
  wire  bundleOut_0_a_sink__EVAL_20;
  wire [31:0] bundleOut_0_a_sink__EVAL_21;
  wire [31:0] bundleOut_0_a_sink__EVAL_22;
  wire  bundleOut_0_a_sink__EVAL_23;
  wire [31:0] bundleOut_0_a_sink__EVAL_24;
  wire  bundleOut_0_a_sink__EVAL_25;
  wire [3:0] bundleOut_0_a_sink__EVAL_26;
  wire [2:0] bundleOut_0_a_sink__EVAL_27;
  wire  bundleOut_0_a_sink__EVAL_28;
  wire [1:0] bundleOut_0_a_sink__EVAL_29;
  wire  bundleOut_0_a_sink__EVAL_30;
  wire [3:0] bundleOut_0_a_sink__EVAL_31;
  wire [2:0] bundleOut_0_a_sink__EVAL_32;
  wire  bundleOut_0_a_sink__EVAL_33;
  wire  bundleOut_0_a_sink__EVAL_34;
  wire [1:0] bundleOut_0_a_sink__EVAL_35;
  wire [3:0] bundleOut_0_a_sink__EVAL_36;
  wire [2:0] bundleOut_0_a_sink__EVAL_37;
  wire  bundleOut_0_a_sink__EVAL_38;
  wire [31:0] bundleOut_0_a_sink__EVAL_39;
  wire  bundleOut_0_a_sink__EVAL_40;
  wire [3:0] bundleOut_0_a_sink__EVAL_41;
  wire [3:0] bundleOut_0_a_sink__EVAL_42;
  wire [1:0] bundleIn_0_d_source__EVAL;
  wire [1:0] bundleIn_0_d_source__EVAL_0;
  wire [1:0] bundleIn_0_d_source__EVAL_1;
  wire [2:0] bundleIn_0_d_source__EVAL_2;
  wire  bundleIn_0_d_source__EVAL_3;
  wire  bundleIn_0_d_source__EVAL_4;
  wire [2:0] bundleIn_0_d_source__EVAL_5;
  wire  bundleIn_0_d_source__EVAL_6;
  wire [1:0] bundleIn_0_d_source__EVAL_7;
  wire  bundleIn_0_d_source__EVAL_8;
  wire [31:0] bundleIn_0_d_source__EVAL_9;
  wire  bundleIn_0_d_source__EVAL_10;
  wire  bundleIn_0_d_source__EVAL_11;
  wire [3:0] bundleIn_0_d_source__EVAL_12;
  wire  bundleIn_0_d_source__EVAL_13;
  wire  bundleIn_0_d_source__EVAL_14;
  wire [1:0] bundleIn_0_d_source__EVAL_15;
  wire  bundleIn_0_d_source__EVAL_16;
  wire [3:0] bundleIn_0_d_source__EVAL_17;
  wire [31:0] bundleIn_0_d_source__EVAL_18;
  wire  bundleIn_0_d_source__EVAL_19;
  wire  bundleIn_0_d_source__EVAL_20;
  wire  bundleIn_0_d_source__EVAL_21;
  wire [3:0] bundleIn_0_d_source__EVAL_22;
  wire  bundleIn_0_d_source__EVAL_23;
  wire [31:0] bundleIn_0_d_source__EVAL_24;
  wire [3:0] bundleIn_0_d_source__EVAL_25;
  wire [3:0] bundleIn_0_d_source__EVAL_26;
  wire [3:0] bundleIn_0_d_source__EVAL_27;
  wire [2:0] bundleIn_0_d_source__EVAL_28;
  wire  bundleIn_0_d_source__EVAL_29;
  wire  bundleIn_0_d_source__EVAL_30;
  _EVAL_8 bundleOut_0_a_sink (
    ._EVAL(bundleOut_0_a_sink__EVAL),
    ._EVAL_0(bundleOut_0_a_sink__EVAL_0),
    ._EVAL_1(bundleOut_0_a_sink__EVAL_1),
    ._EVAL_2(bundleOut_0_a_sink__EVAL_2),
    ._EVAL_3(bundleOut_0_a_sink__EVAL_3),
    ._EVAL_4(bundleOut_0_a_sink__EVAL_4),
    ._EVAL_5(bundleOut_0_a_sink__EVAL_5),
    ._EVAL_6(bundleOut_0_a_sink__EVAL_6),
    ._EVAL_7(bundleOut_0_a_sink__EVAL_7),
    ._EVAL_8(bundleOut_0_a_sink__EVAL_8),
    ._EVAL_9(bundleOut_0_a_sink__EVAL_9),
    ._EVAL_10(bundleOut_0_a_sink__EVAL_10),
    ._EVAL_11(bundleOut_0_a_sink__EVAL_11),
    ._EVAL_12(bundleOut_0_a_sink__EVAL_12),
    ._EVAL_13(bundleOut_0_a_sink__EVAL_13),
    ._EVAL_14(bundleOut_0_a_sink__EVAL_14),
    ._EVAL_15(bundleOut_0_a_sink__EVAL_15),
    ._EVAL_16(bundleOut_0_a_sink__EVAL_16),
    ._EVAL_17(bundleOut_0_a_sink__EVAL_17),
    ._EVAL_18(bundleOut_0_a_sink__EVAL_18),
    ._EVAL_19(bundleOut_0_a_sink__EVAL_19),
    ._EVAL_20(bundleOut_0_a_sink__EVAL_20),
    ._EVAL_21(bundleOut_0_a_sink__EVAL_21),
    ._EVAL_22(bundleOut_0_a_sink__EVAL_22),
    ._EVAL_23(bundleOut_0_a_sink__EVAL_23),
    ._EVAL_24(bundleOut_0_a_sink__EVAL_24),
    ._EVAL_25(bundleOut_0_a_sink__EVAL_25),
    ._EVAL_26(bundleOut_0_a_sink__EVAL_26),
    ._EVAL_27(bundleOut_0_a_sink__EVAL_27),
    ._EVAL_28(bundleOut_0_a_sink__EVAL_28),
    ._EVAL_29(bundleOut_0_a_sink__EVAL_29),
    ._EVAL_30(bundleOut_0_a_sink__EVAL_30),
    ._EVAL_31(bundleOut_0_a_sink__EVAL_31),
    ._EVAL_32(bundleOut_0_a_sink__EVAL_32),
    ._EVAL_33(bundleOut_0_a_sink__EVAL_33),
    ._EVAL_34(bundleOut_0_a_sink__EVAL_34),
    ._EVAL_35(bundleOut_0_a_sink__EVAL_35),
    ._EVAL_36(bundleOut_0_a_sink__EVAL_36),
    ._EVAL_37(bundleOut_0_a_sink__EVAL_37),
    ._EVAL_38(bundleOut_0_a_sink__EVAL_38),
    ._EVAL_39(bundleOut_0_a_sink__EVAL_39),
    ._EVAL_40(bundleOut_0_a_sink__EVAL_40),
    ._EVAL_41(bundleOut_0_a_sink__EVAL_41),
    ._EVAL_42(bundleOut_0_a_sink__EVAL_42)
  );
  _EVAL_10 bundleIn_0_d_source (
    ._EVAL(bundleIn_0_d_source__EVAL),
    ._EVAL_0(bundleIn_0_d_source__EVAL_0),
    ._EVAL_1(bundleIn_0_d_source__EVAL_1),
    ._EVAL_2(bundleIn_0_d_source__EVAL_2),
    ._EVAL_3(bundleIn_0_d_source__EVAL_3),
    ._EVAL_4(bundleIn_0_d_source__EVAL_4),
    ._EVAL_5(bundleIn_0_d_source__EVAL_5),
    ._EVAL_6(bundleIn_0_d_source__EVAL_6),
    ._EVAL_7(bundleIn_0_d_source__EVAL_7),
    ._EVAL_8(bundleIn_0_d_source__EVAL_8),
    ._EVAL_9(bundleIn_0_d_source__EVAL_9),
    ._EVAL_10(bundleIn_0_d_source__EVAL_10),
    ._EVAL_11(bundleIn_0_d_source__EVAL_11),
    ._EVAL_12(bundleIn_0_d_source__EVAL_12),
    ._EVAL_13(bundleIn_0_d_source__EVAL_13),
    ._EVAL_14(bundleIn_0_d_source__EVAL_14),
    ._EVAL_15(bundleIn_0_d_source__EVAL_15),
    ._EVAL_16(bundleIn_0_d_source__EVAL_16),
    ._EVAL_17(bundleIn_0_d_source__EVAL_17),
    ._EVAL_18(bundleIn_0_d_source__EVAL_18),
    ._EVAL_19(bundleIn_0_d_source__EVAL_19),
    ._EVAL_20(bundleIn_0_d_source__EVAL_20),
    ._EVAL_21(bundleIn_0_d_source__EVAL_21),
    ._EVAL_22(bundleIn_0_d_source__EVAL_22),
    ._EVAL_23(bundleIn_0_d_source__EVAL_23),
    ._EVAL_24(bundleIn_0_d_source__EVAL_24),
    ._EVAL_25(bundleIn_0_d_source__EVAL_25),
    ._EVAL_26(bundleIn_0_d_source__EVAL_26),
    ._EVAL_27(bundleIn_0_d_source__EVAL_27),
    ._EVAL_28(bundleIn_0_d_source__EVAL_28),
    ._EVAL_29(bundleIn_0_d_source__EVAL_29),
    ._EVAL_30(bundleIn_0_d_source__EVAL_30)
  );
  assign bundleOut_0_a_sink__EVAL_10 = _EVAL_53;
  assign _EVAL_34 = bundleOut_0_a_sink__EVAL_9;
  assign bundleOut_0_a_sink__EVAL_1 = _EVAL_63;
  assign _EVAL_69 = bundleIn_0_d_source__EVAL_6;
  assign _EVAL_52 = bundleOut_0_a_sink__EVAL_12;
  assign bundleOut_0_a_sink__EVAL_38 = _EVAL_15;
  assign bundleOut_0_a_sink__EVAL_15 = _EVAL_7;
  assign _EVAL_44 = bundleIn_0_d_source__EVAL_17;
  assign _EVAL_64 = bundleOut_0_a_sink__EVAL_39;
  assign _EVAL_62 = bundleOut_0_a_sink__EVAL_29;
  assign _EVAL_14 = bundleIn_0_d_source__EVAL_26;
  assign bundleOut_0_a_sink__EVAL_31 = _EVAL_51;
  assign bundleOut_0_a_sink__EVAL_19 = _EVAL_26;
  assign bundleOut_0_a_sink__EVAL_21 = _EVAL_71;
  assign _EVAL_32 = bundleIn_0_d_source__EVAL_15;
  assign bundleOut_0_a_sink__EVAL_35 = _EVAL_3;
  assign bundleIn_0_d_source__EVAL_18 = _EVAL_0;
  assign bundleIn_0_d_source__EVAL_25 = _EVAL_9;
  assign _EVAL_1 = bundleIn_0_d_source__EVAL_1;
  assign bundleIn_0_d_source__EVAL_28 = _EVAL_61;
  assign _EVAL_2 = bundleOut_0_a_sink__EVAL_25;
  assign _EVAL_10 = bundleOut_0_a_sink__EVAL_2;
  assign _EVAL_8 = bundleOut_0_a_sink__EVAL_5;
  assign _EVAL_22 = bundleOut_0_a_sink__EVAL_41;
  assign _EVAL_58 = bundleIn_0_d_source__EVAL_13;
  assign _EVAL_67 = bundleIn_0_d_source__EVAL_30;
  assign bundleOut_0_a_sink__EVAL_20 = _EVAL_13;
  assign bundleOut_0_a_sink__EVAL_18 = _EVAL_59;
  assign bundleOut_0_a_sink__EVAL_4 = _EVAL_18;
  assign bundleIn_0_d_source__EVAL_20 = _EVAL_16;
  assign bundleOut_0_a_sink__EVAL_22 = _EVAL_72;
  assign bundleIn_0_d_source__EVAL_3 = _EVAL_65;
  assign _EVAL_56 = bundleOut_0_a_sink__EVAL_33;
  assign _EVAL_43 = bundleIn_0_d_source__EVAL_9;
  assign bundleIn_0_d_source__EVAL_4 = _EVAL_31;
  assign bundleOut_0_a_sink__EVAL_36 = _EVAL_40;
  assign bundleOut_0_a_sink__EVAL_37 = _EVAL_25;
  assign bundleIn_0_d_source__EVAL_12 = _EVAL;
  assign _EVAL_38 = bundleOut_0_a_sink__EVAL_17;
  assign bundleOut_0_a_sink__EVAL_34 = _EVAL_50;
  assign bundleIn_0_d_source__EVAL_23 = _EVAL_13;
  assign bundleIn_0_d_source__EVAL = _EVAL_66;
  assign _EVAL_12 = bundleOut_0_a_sink__EVAL_32;
  assign bundleOut_0_a_sink__EVAL_23 = _EVAL_36;
  assign bundleOut_0_a_sink__EVAL_30 = _EVAL_11;
  assign _EVAL_27 = bundleIn_0_d_source__EVAL_22;
  assign bundleIn_0_d_source__EVAL_14 = _EVAL_63;
  assign _EVAL_46 = bundleIn_0_d_source__EVAL_24;
  assign bundleOut_0_a_sink__EVAL_24 = _EVAL_33;
  assign _EVAL_29 = bundleIn_0_d_source__EVAL_2;
  assign _EVAL_24 = bundleIn_0_d_source__EVAL_29;
  assign bundleOut_0_a_sink__EVAL_27 = _EVAL_48;
  assign bundleOut_0_a_sink__EVAL_6 = _EVAL_37;
  assign _EVAL_30 = bundleOut_0_a_sink__EVAL_14;
  assign bundleOut_0_a_sink__EVAL_16 = _EVAL_42;
  assign bundleOut_0_a_sink__EVAL_7 = _EVAL_55;
  assign bundleOut_0_a_sink__EVAL_13 = _EVAL_39;
  assign bundleIn_0_d_source__EVAL_21 = _EVAL_60;
  assign bundleOut_0_a_sink__EVAL_11 = _EVAL_4;
  assign _EVAL_6 = bundleIn_0_d_source__EVAL_5;
  assign _EVAL_45 = bundleOut_0_a_sink__EVAL;
  assign _EVAL_49 = bundleIn_0_d_source__EVAL_27;
  assign bundleOut_0_a_sink__EVAL_26 = _EVAL_19;
  assign _EVAL_57 = bundleIn_0_d_source__EVAL_7;
  assign bundleOut_0_a_sink__EVAL_40 = _EVAL_54;
  assign _EVAL_70 = bundleOut_0_a_sink__EVAL_8;
  assign bundleOut_0_a_sink__EVAL_42 = _EVAL_35;
  assign bundleOut_0_a_sink__EVAL_3 = _EVAL_28;
  assign _EVAL_5 = bundleIn_0_d_source__EVAL_8;
  assign bundleOut_0_a_sink__EVAL_28 = _EVAL_23;
  assign _EVAL_17 = bundleIn_0_d_source__EVAL_19;
  assign _EVAL_68 = bundleIn_0_d_source__EVAL_10;
  assign bundleIn_0_d_source__EVAL_11 = _EVAL_41;
  assign _EVAL_20 = bundleOut_0_a_sink__EVAL_0;
  assign bundleIn_0_d_source__EVAL_0 = _EVAL_47;
  assign _EVAL_21 = bundleIn_0_d_source__EVAL_16;
endmodule
