//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_184(
  output        _EVAL,
  input  [9:0]  _EVAL_0,
  output [31:0] _EVAL_1,
  input         _EVAL_2,
  output [9:0]  _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input  [7:0]  _EVAL_6,
  output [3:0]  _EVAL_7,
  output [1:0]  _EVAL_8,
  output [7:0]  _EVAL_9,
  input         _EVAL_10,
  input  [8:0]  _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  output        _EVAL_15,
  input  [31:0] _EVAL_16,
  output        _EVAL_17,
  output [2:0]  _EVAL_18,
  output [31:0] _EVAL_19,
  input         _EVAL_20,
  input  [11:0] _EVAL_21,
  input         _EVAL_22,
  output [2:0]  _EVAL_23,
  output        _EVAL_24,
  input  [3:0]  _EVAL_25,
  output        _EVAL_26,
  input         _EVAL_27,
  input         _EVAL_28,
  output [31:0] _EVAL_29,
  input         _EVAL_30,
  input         _EVAL_31,
  input         _EVAL_32,
  input  [31:0] _EVAL_33,
  output        _EVAL_34,
  input  [1:0]  _EVAL_35,
  output [2:0]  _EVAL_36,
  input         _EVAL_37,
  input         _EVAL_38,
  input  [2:0]  _EVAL_39,
  output        _EVAL_40,
  input         _EVAL_41,
  input  [2:0]  _EVAL_42,
  input         _EVAL_43,
  input         _EVAL_44,
  output        _EVAL_45,
  output        _EVAL_46,
  input         _EVAL_47,
  output [1:0]  _EVAL_48
);
  wire [1:0] dmiXing__EVAL;
  wire [31:0] dmiXing__EVAL_0;
  wire  dmiXing__EVAL_1;
  wire [31:0] dmiXing__EVAL_2;
  wire  dmiXing__EVAL_3;
  wire  dmiXing__EVAL_4;
  wire [2:0] dmiXing__EVAL_5;
  wire [1:0] dmiXing__EVAL_6;
  wire  dmiXing__EVAL_7;
  wire [31:0] dmiXing__EVAL_8;
  wire  dmiXing__EVAL_9;
  wire [2:0] dmiXing__EVAL_10;
  wire  dmiXing__EVAL_11;
  wire  dmiXing__EVAL_12;
  wire  dmiXing__EVAL_13;
  wire [1:0] dmiXing__EVAL_14;
  wire  dmiXing__EVAL_15;
  wire  dmiXing__EVAL_16;
  wire  dmiXing__EVAL_17;
  wire [2:0] dmiXing__EVAL_18;
  wire [3:0] dmiXing__EVAL_19;
  wire  dmiXing__EVAL_20;
  wire [2:0] dmiXing__EVAL_21;
  wire  dmiXing__EVAL_22;
  wire [8:0] dmiXing__EVAL_23;
  wire [31:0] dmiXing__EVAL_24;
  wire [2:0] dmiXing__EVAL_25;
  wire [8:0] dmiXing__EVAL_26;
  wire  dmiXing__EVAL_27;
  wire  dmactive_synced_dmactive_synced_dmactiveSync__EVAL;
  wire  dmactive_synced_dmactive_synced_dmactiveSync__EVAL_0;
  wire  dmactive_synced_dmactive_synced_dmactiveSync__EVAL_1;
  wire  dmactive_synced_dmactive_synced_dmactiveSync__EVAL_2;
  wire  dmInner__EVAL;
  wire [2:0] dmInner__EVAL_0;
  wire  dmInner__EVAL_1;
  wire  dmInner__EVAL_2;
  wire [2:0] dmInner__EVAL_3;
  wire  dmInner__EVAL_4;
  wire [3:0] dmInner__EVAL_5;
  wire [9:0] dmInner__EVAL_6;
  wire [31:0] dmInner__EVAL_7;
  wire [7:0] dmInner__EVAL_8;
  wire [2:0] dmInner__EVAL_9;
  wire  dmInner__EVAL_10;
  wire [9:0] dmInner__EVAL_11;
  wire [2:0] dmInner__EVAL_12;
  wire [31:0] dmInner__EVAL_13;
  wire  dmInner__EVAL_14;
  wire  dmInner__EVAL_15;
  wire  dmInner__EVAL_16;
  wire  dmInner__EVAL_17;
  wire  dmInner__EVAL_18;
  wire  dmInner__EVAL_19;
  wire  dmInner__EVAL_20;
  wire [1:0] dmInner__EVAL_21;
  wire  dmInner__EVAL_22;
  wire [7:0] dmInner__EVAL_23;
  wire  dmInner__EVAL_24;
  wire [9:0] dmInner__EVAL_25;
  wire [2:0] dmInner__EVAL_26;
  wire [2:0] dmInner__EVAL_27;
  wire  dmInner__EVAL_28;
  wire [31:0] dmInner__EVAL_29;
  wire  dmInner__EVAL_30;
  wire  dmInner__EVAL_31;
  wire [3:0] dmInner__EVAL_32;
  wire [1:0] dmInner__EVAL_33;
  wire  dmInner__EVAL_34;
  wire  dmInner__EVAL_35;
  wire  dmInner__EVAL_36;
  wire  dmInner__EVAL_37;
  wire  dmInner__EVAL_38;
  wire [31:0] dmInner__EVAL_39;
  wire [31:0] dmInner__EVAL_40;
  wire [1:0] dmInner__EVAL_41;
  wire [8:0] dmInner__EVAL_42;
  wire [3:0] dmInner__EVAL_43;
  wire  dmInner__EVAL_44;
  wire  dmInner__EVAL_45;
  wire  dmInner__EVAL_46;
  wire [2:0] dmInner__EVAL_47;
  wire  dmInner__EVAL_48;
  wire [1:0] dmInner__EVAL_49;
  wire  dmInner__EVAL_50;
  wire  dmInner__EVAL_51;
  wire  dmInner__EVAL_52;
  wire  dmInner__EVAL_53;
  wire [11:0] dmInner__EVAL_54;
  wire  dmactive_synced_dmInner_io_innerCtrl_sink__EVAL;
  wire  dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_0;
  wire  dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_1;
  wire  dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_2;
  wire  dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_3;
  wire  dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_4;
  wire  dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_5;
  wire  dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_6;
  wire  dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_7;
  wire  dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_8;
  wire  dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_9;
  wire [9:0] dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_10;
  _EVAL_181 dmiXing (
    ._EVAL(dmiXing__EVAL),
    ._EVAL_0(dmiXing__EVAL_0),
    ._EVAL_1(dmiXing__EVAL_1),
    ._EVAL_2(dmiXing__EVAL_2),
    ._EVAL_3(dmiXing__EVAL_3),
    ._EVAL_4(dmiXing__EVAL_4),
    ._EVAL_5(dmiXing__EVAL_5),
    ._EVAL_6(dmiXing__EVAL_6),
    ._EVAL_7(dmiXing__EVAL_7),
    ._EVAL_8(dmiXing__EVAL_8),
    ._EVAL_9(dmiXing__EVAL_9),
    ._EVAL_10(dmiXing__EVAL_10),
    ._EVAL_11(dmiXing__EVAL_11),
    ._EVAL_12(dmiXing__EVAL_12),
    ._EVAL_13(dmiXing__EVAL_13),
    ._EVAL_14(dmiXing__EVAL_14),
    ._EVAL_15(dmiXing__EVAL_15),
    ._EVAL_16(dmiXing__EVAL_16),
    ._EVAL_17(dmiXing__EVAL_17),
    ._EVAL_18(dmiXing__EVAL_18),
    ._EVAL_19(dmiXing__EVAL_19),
    ._EVAL_20(dmiXing__EVAL_20),
    ._EVAL_21(dmiXing__EVAL_21),
    ._EVAL_22(dmiXing__EVAL_22),
    ._EVAL_23(dmiXing__EVAL_23),
    ._EVAL_24(dmiXing__EVAL_24),
    ._EVAL_25(dmiXing__EVAL_25),
    ._EVAL_26(dmiXing__EVAL_26),
    ._EVAL_27(dmiXing__EVAL_27)
  );
  _EVAL_176 dmactive_synced_dmactive_synced_dmactiveSync (
    ._EVAL(dmactive_synced_dmactive_synced_dmactiveSync__EVAL),
    ._EVAL_0(dmactive_synced_dmactive_synced_dmactiveSync__EVAL_0),
    ._EVAL_1(dmactive_synced_dmactive_synced_dmactiveSync__EVAL_1),
    ._EVAL_2(dmactive_synced_dmactive_synced_dmactiveSync__EVAL_2)
  );
  _EVAL_177 dmInner (
    ._EVAL(dmInner__EVAL),
    ._EVAL_0(dmInner__EVAL_0),
    ._EVAL_1(dmInner__EVAL_1),
    ._EVAL_2(dmInner__EVAL_2),
    ._EVAL_3(dmInner__EVAL_3),
    ._EVAL_4(dmInner__EVAL_4),
    ._EVAL_5(dmInner__EVAL_5),
    ._EVAL_6(dmInner__EVAL_6),
    ._EVAL_7(dmInner__EVAL_7),
    ._EVAL_8(dmInner__EVAL_8),
    ._EVAL_9(dmInner__EVAL_9),
    ._EVAL_10(dmInner__EVAL_10),
    ._EVAL_11(dmInner__EVAL_11),
    ._EVAL_12(dmInner__EVAL_12),
    ._EVAL_13(dmInner__EVAL_13),
    ._EVAL_14(dmInner__EVAL_14),
    ._EVAL_15(dmInner__EVAL_15),
    ._EVAL_16(dmInner__EVAL_16),
    ._EVAL_17(dmInner__EVAL_17),
    ._EVAL_18(dmInner__EVAL_18),
    ._EVAL_19(dmInner__EVAL_19),
    ._EVAL_20(dmInner__EVAL_20),
    ._EVAL_21(dmInner__EVAL_21),
    ._EVAL_22(dmInner__EVAL_22),
    ._EVAL_23(dmInner__EVAL_23),
    ._EVAL_24(dmInner__EVAL_24),
    ._EVAL_25(dmInner__EVAL_25),
    ._EVAL_26(dmInner__EVAL_26),
    ._EVAL_27(dmInner__EVAL_27),
    ._EVAL_28(dmInner__EVAL_28),
    ._EVAL_29(dmInner__EVAL_29),
    ._EVAL_30(dmInner__EVAL_30),
    ._EVAL_31(dmInner__EVAL_31),
    ._EVAL_32(dmInner__EVAL_32),
    ._EVAL_33(dmInner__EVAL_33),
    ._EVAL_34(dmInner__EVAL_34),
    ._EVAL_35(dmInner__EVAL_35),
    ._EVAL_36(dmInner__EVAL_36),
    ._EVAL_37(dmInner__EVAL_37),
    ._EVAL_38(dmInner__EVAL_38),
    ._EVAL_39(dmInner__EVAL_39),
    ._EVAL_40(dmInner__EVAL_40),
    ._EVAL_41(dmInner__EVAL_41),
    ._EVAL_42(dmInner__EVAL_42),
    ._EVAL_43(dmInner__EVAL_43),
    ._EVAL_44(dmInner__EVAL_44),
    ._EVAL_45(dmInner__EVAL_45),
    ._EVAL_46(dmInner__EVAL_46),
    ._EVAL_47(dmInner__EVAL_47),
    ._EVAL_48(dmInner__EVAL_48),
    ._EVAL_49(dmInner__EVAL_49),
    ._EVAL_50(dmInner__EVAL_50),
    ._EVAL_51(dmInner__EVAL_51),
    ._EVAL_52(dmInner__EVAL_52),
    ._EVAL_53(dmInner__EVAL_53),
    ._EVAL_54(dmInner__EVAL_54)
  );
  _EVAL_183 dmactive_synced_dmInner_io_innerCtrl_sink (
    ._EVAL(dmactive_synced_dmInner_io_innerCtrl_sink__EVAL),
    ._EVAL_0(dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_0),
    ._EVAL_1(dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_1),
    ._EVAL_2(dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_2),
    ._EVAL_3(dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_3),
    ._EVAL_4(dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_4),
    ._EVAL_5(dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_5),
    ._EVAL_6(dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_6),
    ._EVAL_7(dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_7),
    ._EVAL_8(dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_8),
    ._EVAL_9(dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_9),
    ._EVAL_10(dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_10)
  );
  assign _EVAL_1 = dmInner__EVAL_13;
  assign dmiXing__EVAL_11 = dmInner__EVAL_2;
  assign dmInner__EVAL_32 = _EVAL_25;
  assign dmiXing__EVAL_14 = dmInner__EVAL_41;
  assign dmiXing__EVAL_2 = _EVAL_16;
  assign dmiXing__EVAL_22 = _EVAL_28;
  assign dmiXing__EVAL_13 = _EVAL_32;
  assign dmInner__EVAL_3 = dmiXing__EVAL_10;
  assign _EVAL_36 = dmInner__EVAL_0;
  assign _EVAL_48 = dmiXing__EVAL_6;
  assign dmactive_synced_dmactive_synced_dmactiveSync__EVAL_2 = _EVAL_43;
  assign dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_9 = _EVAL_37;
  assign _EVAL_26 = dmInner__EVAL_52;
  assign _EVAL_23 = dmiXing__EVAL_25;
  assign dmiXing__EVAL_15 = dmInner__EVAL_16;
  assign dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_6 = _EVAL_2;
  assign dmInner__EVAL_49 = _EVAL_35;
  assign dmiXing__EVAL_18 = dmInner__EVAL_12;
  assign dmInner__EVAL_30 = _EVAL_10;
  assign dmInner__EVAL_19 = _EVAL_31;
  assign dmiXing__EVAL_4 = _EVAL_10;
  assign dmactive_synced_dmactive_synced_dmactiveSync__EVAL_1 = _EVAL_10;
  assign dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_7 = _EVAL_30;
  assign dmInner__EVAL_15 = _EVAL_41;
  assign _EVAL_18 = dmInner__EVAL_47;
  assign dmInner__EVAL_35 = _EVAL_44;
  assign dmiXing__EVAL_20 = _EVAL_27;
  assign dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_2 = _EVAL_10;
  assign _EVAL_29 = dmiXing__EVAL_24;
  assign dmInner__EVAL_33 = dmiXing__EVAL;
  assign dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_5 = _EVAL_13;
  assign _EVAL_34 = dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_8;
  assign dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_1 = _EVAL_28;
  assign dmInner__EVAL_8 = _EVAL_6;
  assign _EVAL_46 = dmInner__EVAL_24;
  assign _EVAL_45 = dmInner__EVAL_22;
  assign dmInner__EVAL_9 = _EVAL_39;
  assign _EVAL_19 = dmInner__EVAL_7;
  assign dmInner__EVAL_43 = dmiXing__EVAL_19;
  assign dmInner__EVAL_54 = _EVAL_21;
  assign _EVAL = dmiXing__EVAL_7;
  assign dmInner__EVAL_20 = dmactive_synced_dmactive_synced_dmactiveSync__EVAL;
  assign dmInner__EVAL_18 = _EVAL_14;
  assign dmInner__EVAL_45 = dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_4;
  assign dmInner__EVAL_38 = _EVAL_5;
  assign _EVAL_3 = dmInner__EVAL_25;
  assign dmInner__EVAL_6 = _EVAL_0;
  assign _EVAL_15 = dmInner__EVAL_46;
  assign dmInner__EVAL_4 = _EVAL_47;
  assign dmInner__EVAL_50 = _EVAL_4;
  assign dmiXing__EVAL_26 = _EVAL_11;
  assign dmInner__EVAL = dmiXing__EVAL_3;
  assign dmiXing__EVAL_12 = dmInner__EVAL_37;
  assign dmInner__EVAL_14 = _EVAL_28;
  assign dmInner__EVAL_27 = _EVAL_12;
  assign dmiXing__EVAL_8 = dmInner__EVAL_29;
  assign dmInner__EVAL_36 = dmiXing__EVAL_17;
  assign _EVAL_24 = dmiXing__EVAL_27;
  assign dmInner__EVAL_1 = _EVAL_22;
  assign dmInner__EVAL_11 = dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_10;
  assign _EVAL_7 = dmInner__EVAL_5;
  assign dmInner__EVAL_53 = dmactive_synced_dmInner_io_innerCtrl_sink__EVAL;
  assign dmInner__EVAL_42 = dmiXing__EVAL_23;
  assign _EVAL_8 = dmInner__EVAL_21;
  assign dmInner__EVAL_26 = dmiXing__EVAL_21;
  assign _EVAL_17 = dmiXing__EVAL_16;
  assign dmInner__EVAL_39 = dmiXing__EVAL_0;
  assign _EVAL_40 = dmInner__EVAL_10;
  assign dmInner__EVAL_51 = _EVAL_20;
  assign dmiXing__EVAL_5 = _EVAL_42;
  assign dmInner__EVAL_40 = _EVAL_33;
  assign dmInner__EVAL_48 = dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_3;
  assign dmInner__EVAL_31 = dmiXing__EVAL_9;
  assign dmInner__EVAL_17 = dmiXing__EVAL_1;
  assign dmInner__EVAL_44 = dmactive_synced_dmInner_io_innerCtrl_sink__EVAL_0;
  assign _EVAL_9 = dmInner__EVAL_23;
  assign dmactive_synced_dmactive_synced_dmactiveSync__EVAL_0 = _EVAL_28;
  assign dmInner__EVAL_34 = _EVAL_38;
endmodule
