//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_149(
  output [4:0]  _EVAL,
  input  [2:0]  _EVAL_0,
  input         _EVAL_1,
  input  [31:0] _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  output [2:0]  _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  input  [31:0] _EVAL_8,
  input  [31:0] _EVAL_9,
  input  [1:0]  _EVAL_10,
  output [2:0]  _EVAL_11,
  output        _EVAL_12,
  input  [2:0]  _EVAL_13,
  input  [3:0]  _EVAL_14,
  output [2:0]  _EVAL_15,
  output        _EVAL_16,
  output [31:0] _EVAL_17,
  input  [31:0] _EVAL_18,
  output        _EVAL_19,
  output        _EVAL_20,
  input         _EVAL_21,
  output        _EVAL_22,
  input  [4:0]  _EVAL_23,
  input         _EVAL_24,
  input  [1:0]  _EVAL_25,
  output [2:0]  _EVAL_26,
  output [31:0] _EVAL_27,
  output        _EVAL_28,
  input         _EVAL_29,
  input  [2:0]  _EVAL_30,
  output [3:0]  _EVAL_31,
  input         _EVAL_32,
  output [3:0]  _EVAL_33,
  output [31:0] _EVAL_34,
  output        _EVAL_35,
  input         _EVAL_36,
  input         _EVAL_37,
  output [3:0]  _EVAL_38,
  input         _EVAL_39,
  input         _EVAL_40,
  input  [4:0]  _EVAL_41,
  output        _EVAL_42,
  input         _EVAL_43,
  input         _EVAL_44,
  output        _EVAL_45,
  output        _EVAL_46,
  output [3:0]  _EVAL_47,
  input         _EVAL_48,
  input  [1:0]  _EVAL_49,
  output        _EVAL_50,
  output [3:0]  _EVAL_51,
  input         _EVAL_52,
  input         _EVAL_53,
  output [2:0]  _EVAL_54,
  input  [31:0] _EVAL_55,
  output        _EVAL_56,
  input         _EVAL_57,
  input  [2:0]  _EVAL_58,
  input         _EVAL_59,
  output [2:0]  _EVAL_60,
  input         _EVAL_61,
  output [1:0]  _EVAL_62,
  input         _EVAL_63,
  input         _EVAL_64,
  input  [3:0]  _EVAL_65,
  input  [2:0]  _EVAL_66,
  input  [3:0]  _EVAL_67,
  input         _EVAL_68,
  input  [1:0]  _EVAL_69,
  output        _EVAL_70,
  output [2:0]  _EVAL_71,
  input  [3:0]  _EVAL_72,
  input         _EVAL_73,
  input         _EVAL_74,
  input  [1:0]  _EVAL_75,
  output        _EVAL_76,
  input         _EVAL_77,
  input  [3:0]  _EVAL_78,
  output [1:0]  _EVAL_79,
  output        _EVAL_80,
  output [31:0] _EVAL_81,
  output [2:0]  _EVAL_82,
  input  [1:0]  _EVAL_83,
  output        _EVAL_84,
  input         _EVAL_85,
  input  [31:0] _EVAL_86,
  input  [31:0] _EVAL_87,
  output [31:0] _EVAL_88,
  input         _EVAL_89,
  input         _EVAL_90,
  input  [31:0] _EVAL_91,
  output [1:0]  _EVAL_92,
  input         _EVAL_93,
  input         _EVAL_94,
  input         _EVAL_95,
  output        _EVAL_96,
  output [3:0]  _EVAL_97,
  output [1:0]  _EVAL_98,
  output        _EVAL_99,
  input         _EVAL_100,
  input  [31:0] _EVAL_101,
  input  [3:0]  _EVAL_102,
  input  [2:0]  _EVAL_103,
  input         _EVAL_104,
  output [4:0]  _EVAL_105,
  input  [2:0]  _EVAL_106,
  input         _EVAL_107,
  output [31:0] _EVAL_108
);
  wire  _EVAL_109;
  wire [2:0] _EVAL_110;
  wire  rsource__EVAL;
  wire [3:0] rsource__EVAL_0;
  wire  rsource__EVAL_1;
  wire [2:0] rsource__EVAL_2;
  wire [3:0] rsource__EVAL_3;
  wire  rsource__EVAL_4;
  wire [1:0] rsource__EVAL_5;
  wire  rsource__EVAL_6;
  wire [3:0] rsource__EVAL_7;
  wire [1:0] rsource__EVAL_8;
  wire  rsource__EVAL_9;
  wire [31:0] rsource__EVAL_10;
  wire  rsource__EVAL_11;
  wire [3:0] rsource__EVAL_12;
  wire  rsource__EVAL_13;
  wire  rsource__EVAL_14;
  wire [2:0] rsource__EVAL_15;
  wire [2:0] rsource__EVAL_16;
  wire  rsource__EVAL_17;
  wire  rsource__EVAL_18;
  wire [3:0] rsource__EVAL_19;
  wire [31:0] rsource__EVAL_20;
  wire  rsource__EVAL_21;
  wire [3:0] rsource__EVAL_22;
  wire  rsource__EVAL_23;
  wire [1:0] rsource__EVAL_24;
  wire [31:0] rsource__EVAL_25;
  wire  rsource__EVAL_26;
  wire  rsource__EVAL_27;
  wire [3:0] rsource__EVAL_28;
  wire [2:0] rsource__EVAL_29;
  wire  rsource__EVAL_30;
  wire  rsource__EVAL_31;
  wire  rsource__EVAL_32;
  wire  rsource__EVAL_33;
  wire [3:0] rsource__EVAL_34;
  wire [3:0] rsource__EVAL_35;
  wire  rsource__EVAL_36;
  wire [31:0] rsource__EVAL_37;
  wire  rsource__EVAL_38;
  wire [31:0] rsource__EVAL_39;
  wire  rsource__EVAL_40;
  wire [2:0] rsource__EVAL_41;
  wire  rsource__EVAL_42;
  wire  rsource__EVAL_43;
  wire [2:0] rsource__EVAL_44;
  wire [31:0] rsource__EVAL_45;
  wire  rsource__EVAL_46;
  wire  rsource__EVAL_47;
  wire [3:0] rsource__EVAL_48;
  wire  rsource__EVAL_49;
  wire [1:0] rsource__EVAL_50;
  wire [31:0] rsource__EVAL_51;
  wire  rsource__EVAL_52;
  wire [2:0] rsource__EVAL_53;
  wire [2:0] rsource__EVAL_54;
  wire [31:0] rsource__EVAL_55;
  wire [31:0] rsource__EVAL_56;
  wire [1:0] rsource__EVAL_57;
  wire  rsource__EVAL_58;
  wire [1:0] rsource__EVAL_59;
  wire [3:0] rsource__EVAL_60;
  wire  rsource__EVAL_61;
  wire [3:0] rsource__EVAL_62;
  wire [1:0] rsource__EVAL_63;
  wire  rsource__EVAL_64;
  wire  rsource__EVAL_65;
  wire [3:0] rsource__EVAL_66;
  wire [3:0] rsource__EVAL_67;
  wire  rsource__EVAL_68;
  wire  rsource__EVAL_69;
  wire  rsource__EVAL_70;
  wire [2:0] rsource__EVAL_71;
  wire [3:0] rsource__EVAL_72;
  wire  _EVAL_111;
  wire [2:0] _EVAL_112;
  wire  intsource_1__EVAL;
  wire  intsource_1__EVAL_0;
  wire  _EVAL_113;
  wire [3:0] _EVAL_114;
  wire  _EVAL_115;
  wire [1:0] _EVAL_116;
  wire [2:0] _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire [31:0] _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire [31:0] _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire [2:0] _EVAL_131;
  wire  _EVAL_132;
  wire [3:0] _EVAL_133;
  wire  _EVAL_134;
  wire [2:0] _EVAL_135;
  wire [31:0] _EVAL_136;
  wire  _EVAL_137;
  wire [31:0] _EVAL_138;
  wire [3:0] _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire [2:0] _EVAL_142;
  wire [3:0] _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire [4:0] _EVAL_146;
  wire  _EVAL_147;
  wire [31:0] _EVAL_148;
  wire [31:0] _EVAL_149;
  wire  _EVAL_150;
  wire [3:0] _EVAL_151;
  wire [1:0] _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire [2:0] _EVAL_156;
  wire [3:0] _EVAL_157;
  wire [31:0] _EVAL_158;
  wire [2:0] _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire [31:0] _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  intsink__EVAL;
  wire  intsink__EVAL_0;
  wire  intsink__EVAL_1;
  wire  _EVAL_166;
  wire  intsource_3__EVAL;
  wire  intsource_3__EVAL_0;
  wire [31:0] _EVAL_167;
  wire  _EVAL_168;
  wire [3:0] _EVAL_169;
  wire [31:0] _EVAL_170;
  wire  _EVAL_171;
  wire [4:0] rsink__EVAL;
  wire [2:0] rsink__EVAL_0;
  wire [1:0] rsink__EVAL_1;
  wire  rsink__EVAL_2;
  wire [2:0] rsink__EVAL_3;
  wire [31:0] rsink__EVAL_4;
  wire [31:0] rsink__EVAL_5;
  wire [4:0] rsink__EVAL_6;
  wire [1:0] rsink__EVAL_7;
  wire [2:0] rsink__EVAL_8;
  wire [2:0] rsink__EVAL_9;
  wire [3:0] rsink__EVAL_10;
  wire [1:0] rsink__EVAL_11;
  wire [3:0] rsink__EVAL_12;
  wire [2:0] rsink__EVAL_13;
  wire [31:0] rsink__EVAL_14;
  wire  rsink__EVAL_15;
  wire [31:0] rsink__EVAL_16;
  wire [4:0] rsink__EVAL_17;
  wire  rsink__EVAL_18;
  wire [3:0] rsink__EVAL_19;
  wire [31:0] rsink__EVAL_20;
  wire  rsink__EVAL_21;
  wire [2:0] rsink__EVAL_22;
  wire [2:0] rsink__EVAL_23;
  wire [31:0] rsink__EVAL_24;
  wire [4:0] rsink__EVAL_25;
  wire [4:0] rsink__EVAL_26;
  wire [2:0] rsink__EVAL_27;
  wire  rsink__EVAL_28;
  wire [2:0] rsink__EVAL_29;
  wire  rsink__EVAL_30;
  wire [2:0] rsink__EVAL_31;
  wire  rsink__EVAL_32;
  wire [2:0] rsink__EVAL_33;
  wire [2:0] rsink__EVAL_34;
  wire [31:0] rsink__EVAL_35;
  wire [4:0] rsink__EVAL_36;
  wire [2:0] rsink__EVAL_37;
  wire [31:0] rsink__EVAL_38;
  wire  rsink__EVAL_39;
  wire [31:0] rsink__EVAL_40;
  wire  rsink__EVAL_41;
  wire [2:0] rsink__EVAL_42;
  wire [2:0] rsink__EVAL_43;
  wire  rsink__EVAL_44;
  wire [1:0] rsink__EVAL_45;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire [31:0] _EVAL_175;
  wire [3:0] _EVAL_176;
  wire  _EVAL_177;
  wire [2:0] _EVAL_178;
  wire  _EVAL_179;
  wire [4:0] _EVAL_180;
  wire  _EVAL_181;
  wire  intsink_3__EVAL;
  wire  intsink_3__EVAL_0;
  wire  intsink_3__EVAL_1;
  wire  intsink_3__EVAL_2;
  wire  intsink_3__EVAL_3;
  wire  intsink_3__EVAL_4;
  wire  intsink_3__EVAL_5;
  wire  intsink_3__EVAL_6;
  wire  intsink_3__EVAL_7;
  wire  intsink_3__EVAL_8;
  wire  intsink_3__EVAL_9;
  wire  intsink_3__EVAL_10;
  wire  intsink_3__EVAL_11;
  wire  intsink_3__EVAL_12;
  wire  intsink_3__EVAL_13;
  wire  intsink_3__EVAL_14;
  wire  intsink_3__EVAL_15;
  wire  intsink_3__EVAL_16;
  wire  intsink_3__EVAL_17;
  wire  intsink_3__EVAL_18;
  wire  intsink_3__EVAL_19;
  wire  intsink_3__EVAL_20;
  wire  intsink_3__EVAL_21;
  wire  intsink_3__EVAL_22;
  wire  intsink_3__EVAL_23;
  wire  intsink_3__EVAL_24;
  wire  intsink_3__EVAL_25;
  wire  intsink_3__EVAL_26;
  wire  intsink_3__EVAL_27;
  wire  intsink_3__EVAL_28;
  wire  intsink_3__EVAL_29;
  wire  intsink_3__EVAL_30;
  wire [4:0] _EVAL_182;
  wire [31:0] _EVAL_183;
  wire [2:0] _EVAL_184;
  wire  _EVAL_185;
  wire [2:0] _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  intsource_4__EVAL;
  wire  intsource_4__EVAL_0;
  wire  _EVAL_189;
  wire [2:0] _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire [2:0] _EVAL_195;
  wire  _EVAL_196;
  wire [1:0] _EVAL_197;
  wire [3:0] _EVAL_198;
  wire [2:0] _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire [3:0] _EVAL_202;
  wire [2:0] _EVAL_203;
  wire [31:0] _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire [2:0] _EVAL_207;
  wire  _EVAL_208;
  wire [31:0] _EVAL_209;
  wire [2:0] _EVAL_210;
  wire [4:0] _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire [2:0] _EVAL_214;
  wire  _EVAL_215;
  wire [2:0] _EVAL_216;
  wire  _EVAL_217;
  wire [31:0] _EVAL_218;
  wire [31:0] _EVAL_219;
  wire  _EVAL_220;
  wire [3:0] _EVAL_221;
  wire  _EVAL_222;
  wire [3:0] _EVAL_223;
  wire [3:0] _EVAL_224;
  wire [3:0] _EVAL_225;
  wire  _EVAL_226;
  wire [2:0] _EVAL_227;
  wire  tile__EVAL;
  wire  tile__EVAL_0;
  wire [31:0] tile__EVAL_1;
  wire [31:0] tile__EVAL_2;
  wire  tile__EVAL_3;
  wire  tile__EVAL_4;
  wire  tile__EVAL_5;
  wire  tile__EVAL_6;
  wire  tile__EVAL_7;
  wire [3:0] tile__EVAL_8;
  wire  tile__EVAL_9;
  wire [3:0] tile__EVAL_10;
  wire [31:0] tile__EVAL_11;
  wire  tile__EVAL_12;
  wire  tile__EVAL_13;
  wire  tile__EVAL_14;
  wire  tile__EVAL_15;
  wire  tile__EVAL_16;
  wire  tile__EVAL_17;
  wire  tile__EVAL_18;
  wire  tile__EVAL_19;
  wire [2:0] tile__EVAL_20;
  wire  tile__EVAL_21;
  wire  tile__EVAL_22;
  wire  tile__EVAL_23;
  wire  tile__EVAL_24;
  wire  tile__EVAL_25;
  wire  tile__EVAL_26;
  wire  tile__EVAL_27;
  wire  tile__EVAL_28;
  wire  tile__EVAL_29;
  wire [31:0] tile__EVAL_30;
  wire [2:0] tile__EVAL_31;
  wire  tile__EVAL_32;
  wire  tile__EVAL_33;
  wire [31:0] tile__EVAL_34;
  wire [2:0] tile__EVAL_35;
  wire  tile__EVAL_36;
  wire  tile__EVAL_37;
  wire [2:0] tile__EVAL_38;
  wire [4:0] tile__EVAL_39;
  wire  tile__EVAL_40;
  wire  tile__EVAL_41;
  wire  tile__EVAL_42;
  wire  tile__EVAL_43;
  wire [3:0] tile__EVAL_44;
  wire [31:0] tile__EVAL_45;
  wire [31:0] tile__EVAL_46;
  wire [2:0] tile__EVAL_47;
  wire [3:0] tile__EVAL_48;
  wire  tile__EVAL_49;
  wire  tile__EVAL_50;
  wire [3:0] tile__EVAL_51;
  wire  tile__EVAL_52;
  wire [1:0] tile__EVAL_53;
  wire  tile__EVAL_54;
  wire  tile__EVAL_55;
  wire [31:0] tile__EVAL_56;
  wire  tile__EVAL_57;
  wire [2:0] tile__EVAL_58;
  wire  tile__EVAL_59;
  wire [2:0] tile__EVAL_60;
  wire [3:0] tile__EVAL_61;
  wire  tile__EVAL_62;
  wire [2:0] tile__EVAL_63;
  wire  tile__EVAL_64;
  wire [31:0] tile__EVAL_65;
  wire [4:0] tile__EVAL_66;
  wire  tile__EVAL_67;
  wire  tile__EVAL_68;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  intsink_1__EVAL;
  wire  intsink_1__EVAL_0;
  wire  intsink_1__EVAL_1;
  wire  intsink_1__EVAL_2;
  wire  intsink_1__EVAL_3;
  wire  intsink_1__EVAL_4;
  wire [3:0] _EVAL_230;
  wire [31:0] _EVAL_231;
  wire  _EVAL_232;
  wire [31:0] _EVAL_233;
  wire [31:0] _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire [31:0] _EVAL_237;
  wire [4:0] _EVAL_238;
  wire [3:0] _EVAL_239;
  wire [3:0] _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire [2:0] _EVAL_243;
  wire  intsink_2__EVAL;
  wire  intsink_2__EVAL_0;
  wire  intsink_2__EVAL_1;
  wire  intsink_2__EVAL_2;
  wire  _EVAL_244;
  wire [4:0] _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire [3:0] _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire [2:0] _EVAL_253;
  wire [31:0] _EVAL_254;
  wire [2:0] _EVAL_255;
  wire  _EVAL_256;
  wire [2:0] _EVAL_257;
  wire  _EVAL_258;
  wire  intsource_2__EVAL;
  wire  intsource_2__EVAL_0;
  wire  _EVAL_259;
  wire  _EVAL_260;
  _EVAL_138 rsource (
    ._EVAL(rsource__EVAL),
    ._EVAL_0(rsource__EVAL_0),
    ._EVAL_1(rsource__EVAL_1),
    ._EVAL_2(rsource__EVAL_2),
    ._EVAL_3(rsource__EVAL_3),
    ._EVAL_4(rsource__EVAL_4),
    ._EVAL_5(rsource__EVAL_5),
    ._EVAL_6(rsource__EVAL_6),
    ._EVAL_7(rsource__EVAL_7),
    ._EVAL_8(rsource__EVAL_8),
    ._EVAL_9(rsource__EVAL_9),
    ._EVAL_10(rsource__EVAL_10),
    ._EVAL_11(rsource__EVAL_11),
    ._EVAL_12(rsource__EVAL_12),
    ._EVAL_13(rsource__EVAL_13),
    ._EVAL_14(rsource__EVAL_14),
    ._EVAL_15(rsource__EVAL_15),
    ._EVAL_16(rsource__EVAL_16),
    ._EVAL_17(rsource__EVAL_17),
    ._EVAL_18(rsource__EVAL_18),
    ._EVAL_19(rsource__EVAL_19),
    ._EVAL_20(rsource__EVAL_20),
    ._EVAL_21(rsource__EVAL_21),
    ._EVAL_22(rsource__EVAL_22),
    ._EVAL_23(rsource__EVAL_23),
    ._EVAL_24(rsource__EVAL_24),
    ._EVAL_25(rsource__EVAL_25),
    ._EVAL_26(rsource__EVAL_26),
    ._EVAL_27(rsource__EVAL_27),
    ._EVAL_28(rsource__EVAL_28),
    ._EVAL_29(rsource__EVAL_29),
    ._EVAL_30(rsource__EVAL_30),
    ._EVAL_31(rsource__EVAL_31),
    ._EVAL_32(rsource__EVAL_32),
    ._EVAL_33(rsource__EVAL_33),
    ._EVAL_34(rsource__EVAL_34),
    ._EVAL_35(rsource__EVAL_35),
    ._EVAL_36(rsource__EVAL_36),
    ._EVAL_37(rsource__EVAL_37),
    ._EVAL_38(rsource__EVAL_38),
    ._EVAL_39(rsource__EVAL_39),
    ._EVAL_40(rsource__EVAL_40),
    ._EVAL_41(rsource__EVAL_41),
    ._EVAL_42(rsource__EVAL_42),
    ._EVAL_43(rsource__EVAL_43),
    ._EVAL_44(rsource__EVAL_44),
    ._EVAL_45(rsource__EVAL_45),
    ._EVAL_46(rsource__EVAL_46),
    ._EVAL_47(rsource__EVAL_47),
    ._EVAL_48(rsource__EVAL_48),
    ._EVAL_49(rsource__EVAL_49),
    ._EVAL_50(rsource__EVAL_50),
    ._EVAL_51(rsource__EVAL_51),
    ._EVAL_52(rsource__EVAL_52),
    ._EVAL_53(rsource__EVAL_53),
    ._EVAL_54(rsource__EVAL_54),
    ._EVAL_55(rsource__EVAL_55),
    ._EVAL_56(rsource__EVAL_56),
    ._EVAL_57(rsource__EVAL_57),
    ._EVAL_58(rsource__EVAL_58),
    ._EVAL_59(rsource__EVAL_59),
    ._EVAL_60(rsource__EVAL_60),
    ._EVAL_61(rsource__EVAL_61),
    ._EVAL_62(rsource__EVAL_62),
    ._EVAL_63(rsource__EVAL_63),
    ._EVAL_64(rsource__EVAL_64),
    ._EVAL_65(rsource__EVAL_65),
    ._EVAL_66(rsource__EVAL_66),
    ._EVAL_67(rsource__EVAL_67),
    ._EVAL_68(rsource__EVAL_68),
    ._EVAL_69(rsource__EVAL_69),
    ._EVAL_70(rsource__EVAL_70),
    ._EVAL_71(rsource__EVAL_71),
    ._EVAL_72(rsource__EVAL_72)
  );
  _EVAL_148 intsource_1 (
    ._EVAL(intsource_1__EVAL),
    ._EVAL_0(intsource_1__EVAL_0)
  );
  _EVAL_144 intsink (
    ._EVAL(intsink__EVAL),
    ._EVAL_0(intsink__EVAL_0),
    ._EVAL_1(intsink__EVAL_1)
  );
  _EVAL_148 intsource_3 (
    ._EVAL(intsource_3__EVAL),
    ._EVAL_0(intsource_3__EVAL_0)
  );
  _EVAL_141 rsink (
    ._EVAL(rsink__EVAL),
    ._EVAL_0(rsink__EVAL_0),
    ._EVAL_1(rsink__EVAL_1),
    ._EVAL_2(rsink__EVAL_2),
    ._EVAL_3(rsink__EVAL_3),
    ._EVAL_4(rsink__EVAL_4),
    ._EVAL_5(rsink__EVAL_5),
    ._EVAL_6(rsink__EVAL_6),
    ._EVAL_7(rsink__EVAL_7),
    ._EVAL_8(rsink__EVAL_8),
    ._EVAL_9(rsink__EVAL_9),
    ._EVAL_10(rsink__EVAL_10),
    ._EVAL_11(rsink__EVAL_11),
    ._EVAL_12(rsink__EVAL_12),
    ._EVAL_13(rsink__EVAL_13),
    ._EVAL_14(rsink__EVAL_14),
    ._EVAL_15(rsink__EVAL_15),
    ._EVAL_16(rsink__EVAL_16),
    ._EVAL_17(rsink__EVAL_17),
    ._EVAL_18(rsink__EVAL_18),
    ._EVAL_19(rsink__EVAL_19),
    ._EVAL_20(rsink__EVAL_20),
    ._EVAL_21(rsink__EVAL_21),
    ._EVAL_22(rsink__EVAL_22),
    ._EVAL_23(rsink__EVAL_23),
    ._EVAL_24(rsink__EVAL_24),
    ._EVAL_25(rsink__EVAL_25),
    ._EVAL_26(rsink__EVAL_26),
    ._EVAL_27(rsink__EVAL_27),
    ._EVAL_28(rsink__EVAL_28),
    ._EVAL_29(rsink__EVAL_29),
    ._EVAL_30(rsink__EVAL_30),
    ._EVAL_31(rsink__EVAL_31),
    ._EVAL_32(rsink__EVAL_32),
    ._EVAL_33(rsink__EVAL_33),
    ._EVAL_34(rsink__EVAL_34),
    ._EVAL_35(rsink__EVAL_35),
    ._EVAL_36(rsink__EVAL_36),
    ._EVAL_37(rsink__EVAL_37),
    ._EVAL_38(rsink__EVAL_38),
    ._EVAL_39(rsink__EVAL_39),
    ._EVAL_40(rsink__EVAL_40),
    ._EVAL_41(rsink__EVAL_41),
    ._EVAL_42(rsink__EVAL_42),
    ._EVAL_43(rsink__EVAL_43),
    ._EVAL_44(rsink__EVAL_44),
    ._EVAL_45(rsink__EVAL_45)
  );
  _EVAL_147 intsink_3 (
    ._EVAL(intsink_3__EVAL),
    ._EVAL_0(intsink_3__EVAL_0),
    ._EVAL_1(intsink_3__EVAL_1),
    ._EVAL_2(intsink_3__EVAL_2),
    ._EVAL_3(intsink_3__EVAL_3),
    ._EVAL_4(intsink_3__EVAL_4),
    ._EVAL_5(intsink_3__EVAL_5),
    ._EVAL_6(intsink_3__EVAL_6),
    ._EVAL_7(intsink_3__EVAL_7),
    ._EVAL_8(intsink_3__EVAL_8),
    ._EVAL_9(intsink_3__EVAL_9),
    ._EVAL_10(intsink_3__EVAL_10),
    ._EVAL_11(intsink_3__EVAL_11),
    ._EVAL_12(intsink_3__EVAL_12),
    ._EVAL_13(intsink_3__EVAL_13),
    ._EVAL_14(intsink_3__EVAL_14),
    ._EVAL_15(intsink_3__EVAL_15),
    ._EVAL_16(intsink_3__EVAL_16),
    ._EVAL_17(intsink_3__EVAL_17),
    ._EVAL_18(intsink_3__EVAL_18),
    ._EVAL_19(intsink_3__EVAL_19),
    ._EVAL_20(intsink_3__EVAL_20),
    ._EVAL_21(intsink_3__EVAL_21),
    ._EVAL_22(intsink_3__EVAL_22),
    ._EVAL_23(intsink_3__EVAL_23),
    ._EVAL_24(intsink_3__EVAL_24),
    ._EVAL_25(intsink_3__EVAL_25),
    ._EVAL_26(intsink_3__EVAL_26),
    ._EVAL_27(intsink_3__EVAL_27),
    ._EVAL_28(intsink_3__EVAL_28),
    ._EVAL_29(intsink_3__EVAL_29),
    ._EVAL_30(intsink_3__EVAL_30)
  );
  _EVAL_148 intsource_4 (
    ._EVAL(intsource_4__EVAL),
    ._EVAL_0(intsource_4__EVAL_0)
  );
  _EVAL_134 tile (
    ._EVAL(tile__EVAL),
    ._EVAL_0(tile__EVAL_0),
    ._EVAL_1(tile__EVAL_1),
    ._EVAL_2(tile__EVAL_2),
    ._EVAL_3(tile__EVAL_3),
    ._EVAL_4(tile__EVAL_4),
    ._EVAL_5(tile__EVAL_5),
    ._EVAL_6(tile__EVAL_6),
    ._EVAL_7(tile__EVAL_7),
    ._EVAL_8(tile__EVAL_8),
    ._EVAL_9(tile__EVAL_9),
    ._EVAL_10(tile__EVAL_10),
    ._EVAL_11(tile__EVAL_11),
    ._EVAL_12(tile__EVAL_12),
    ._EVAL_13(tile__EVAL_13),
    ._EVAL_14(tile__EVAL_14),
    ._EVAL_15(tile__EVAL_15),
    ._EVAL_16(tile__EVAL_16),
    ._EVAL_17(tile__EVAL_17),
    ._EVAL_18(tile__EVAL_18),
    ._EVAL_19(tile__EVAL_19),
    ._EVAL_20(tile__EVAL_20),
    ._EVAL_21(tile__EVAL_21),
    ._EVAL_22(tile__EVAL_22),
    ._EVAL_23(tile__EVAL_23),
    ._EVAL_24(tile__EVAL_24),
    ._EVAL_25(tile__EVAL_25),
    ._EVAL_26(tile__EVAL_26),
    ._EVAL_27(tile__EVAL_27),
    ._EVAL_28(tile__EVAL_28),
    ._EVAL_29(tile__EVAL_29),
    ._EVAL_30(tile__EVAL_30),
    ._EVAL_31(tile__EVAL_31),
    ._EVAL_32(tile__EVAL_32),
    ._EVAL_33(tile__EVAL_33),
    ._EVAL_34(tile__EVAL_34),
    ._EVAL_35(tile__EVAL_35),
    ._EVAL_36(tile__EVAL_36),
    ._EVAL_37(tile__EVAL_37),
    ._EVAL_38(tile__EVAL_38),
    ._EVAL_39(tile__EVAL_39),
    ._EVAL_40(tile__EVAL_40),
    ._EVAL_41(tile__EVAL_41),
    ._EVAL_42(tile__EVAL_42),
    ._EVAL_43(tile__EVAL_43),
    ._EVAL_44(tile__EVAL_44),
    ._EVAL_45(tile__EVAL_45),
    ._EVAL_46(tile__EVAL_46),
    ._EVAL_47(tile__EVAL_47),
    ._EVAL_48(tile__EVAL_48),
    ._EVAL_49(tile__EVAL_49),
    ._EVAL_50(tile__EVAL_50),
    ._EVAL_51(tile__EVAL_51),
    ._EVAL_52(tile__EVAL_52),
    ._EVAL_53(tile__EVAL_53),
    ._EVAL_54(tile__EVAL_54),
    ._EVAL_55(tile__EVAL_55),
    ._EVAL_56(tile__EVAL_56),
    ._EVAL_57(tile__EVAL_57),
    ._EVAL_58(tile__EVAL_58),
    ._EVAL_59(tile__EVAL_59),
    ._EVAL_60(tile__EVAL_60),
    ._EVAL_61(tile__EVAL_61),
    ._EVAL_62(tile__EVAL_62),
    ._EVAL_63(tile__EVAL_63),
    ._EVAL_64(tile__EVAL_64),
    ._EVAL_65(tile__EVAL_65),
    ._EVAL_66(tile__EVAL_66),
    ._EVAL_67(tile__EVAL_67),
    ._EVAL_68(tile__EVAL_68)
  );
  _EVAL_145 intsink_1 (
    ._EVAL(intsink_1__EVAL),
    ._EVAL_0(intsink_1__EVAL_0),
    ._EVAL_1(intsink_1__EVAL_1),
    ._EVAL_2(intsink_1__EVAL_2),
    ._EVAL_3(intsink_1__EVAL_3),
    ._EVAL_4(intsink_1__EVAL_4)
  );
  _EVAL_146 intsink_2 (
    ._EVAL(intsink_2__EVAL),
    ._EVAL_0(intsink_2__EVAL_0),
    ._EVAL_1(intsink_2__EVAL_1),
    ._EVAL_2(intsink_2__EVAL_2)
  );
  _EVAL_148 intsource_2 (
    ._EVAL(intsource_2__EVAL),
    ._EVAL_0(intsource_2__EVAL_0)
  );
  assign rsink__EVAL_36 = _EVAL_41;
  assign _EVAL_186 = rsink__EVAL_29;
  assign _EVAL_161 = _EVAL_129;
  assign _EVAL_237 = _EVAL_123;
  assign _EVAL = rsink__EVAL_26;
  assign _EVAL_117 = _EVAL_156;
  assign tile__EVAL_13 = _EVAL_260;
  assign rsource__EVAL_1 = _EVAL_252;
  assign _EVAL_20 = rsource__EVAL_38;
  assign _EVAL_70 = rsource__EVAL_43;
  assign rsource__EVAL_70 = _EVAL_90;
  assign tile__EVAL_57 = _EVAL_166;
  assign _EVAL_120 = rsource__EVAL_45;
  assign _EVAL_142 = _EVAL_159;
  assign _EVAL_198 = _EVAL_240;
  assign intsink_2__EVAL_1 = _EVAL_95;
  assign _EVAL_33 = rsource__EVAL_60;
  assign _EVAL_207 = _EVAL_117;
  assign intsink__EVAL_1 = _EVAL_95;
  assign _EVAL_159 = _EVAL_203;
  assign _EVAL_245 = _EVAL_211;
  assign rsource__EVAL_55 = _EVAL_163;
  assign _EVAL_175 = _EVAL_91;
  assign _EVAL_187 = _EVAL_174;
  assign rsource__EVAL_52 = _EVAL_193;
  assign _EVAL_135 = _EVAL_112;
  assign _EVAL_185 = intsink_3__EVAL_9;
  assign _EVAL_22 = rsink__EVAL_30;
  assign _EVAL_50 = rsource__EVAL_13;
  assign _EVAL_143 = rsink__EVAL_10;
  assign _EVAL_130 = rsource__EVAL_18;
  assign _EVAL_97 = rsource__EVAL_67;
  assign tile__EVAL_54 = _EVAL_194;
  assign _EVAL_148 = _EVAL_183;
  assign _EVAL_125 = _EVAL_241;
  assign _EVAL_80 = intsource_2__EVAL;
  assign _EVAL_201 = tile__EVAL;
  assign _EVAL_155 = _EVAL_48;
  assign tile__EVAL_5 = _EVAL_220;
  assign tile__EVAL_58 = _EVAL_110;
  assign _EVAL_19 = rsink__EVAL_32;
  assign intsource_2__EVAL_0 = _EVAL_134;
  assign _EVAL_46 = intsource_1__EVAL;
  assign _EVAL_84 = rsource__EVAL_4;
  assign tile__EVAL_37 = _EVAL_236;
  assign _EVAL_222 = _EVAL_137;
  assign rsink__EVAL_27 = _EVAL_13;
  assign rsource__EVAL_63 = _EVAL_69;
  assign _EVAL_152 = rsource__EVAL_24;
  assign _EVAL_184 = tile__EVAL_63;
  assign _EVAL_205 = tile__EVAL_12;
  assign _EVAL_35 = rsource__EVAL_11;
  assign _EVAL_188 = tile__EVAL_0;
  assign _EVAL_200 = _EVAL_232;
  assign rsource__EVAL_40 = _EVAL_104;
  assign _EVAL_111 = intsink_1__EVAL_4;
  assign _EVAL_172 = intsink_3__EVAL_25;
  assign _EVAL_109 = _EVAL_95;
  assign _EVAL_212 = intsink_3__EVAL_8;
  assign tile__EVAL_30 = _EVAL_138;
  assign _EVAL_141 = intsink_1__EVAL_3;
  assign tile__EVAL_22 = _EVAL_217;
  assign _EVAL_254 = _EVAL_120;
  assign tile__EVAL_7 = _EVAL_172;
  assign _EVAL_257 = _EVAL_184;
  assign _EVAL_112 = _EVAL_195;
  assign _EVAL_158 = _EVAL_254;
  assign _EVAL_38 = rsource__EVAL_48;
  assign rsource__EVAL_23 = _EVAL_249;
  assign intsource_4__EVAL_0 = _EVAL_205;
  assign _EVAL_137 = rsource__EVAL_17;
  assign _EVAL_136 = _EVAL_234;
  assign rsource__EVAL_0 = _EVAL_157;
  assign rsource__EVAL_61 = _EVAL_127;
  assign _EVAL_174 = tile__EVAL_3;
  assign rsink__EVAL_45 = _EVAL_25;
  assign _EVAL_145 = _EVAL_187;
  assign rsource__EVAL_20 = _EVAL_55;
  assign rsink__EVAL_22 = _EVAL_30;
  assign _EVAL_131 = _EVAL_178;
  assign rsource__EVAL_54 = _EVAL_207;
  assign intsink_3__EVAL_10 = _EVAL_37;
  assign tile__EVAL_21 = _EVAL_191;
  assign intsource_3__EVAL_0 = _EVAL_229;
  assign tile__EVAL_42 = _EVAL_185;
  assign _EVAL_166 = _EVAL_100;
  assign _EVAL_194 = _EVAL_160;
  assign _EVAL_147 = _EVAL_226;
  assign _EVAL_121 = _EVAL_130;
  assign rsink__EVAL_13 = _EVAL_7;
  assign _EVAL_79 = rsource__EVAL_50;
  assign rsink__EVAL_28 = _EVAL_113;
  assign tile__EVAL_50 = _EVAL_228;
  assign _EVAL_216 = _EVAL_257;
  assign intsink_3__EVAL_2 = _EVAL_32;
  assign _EVAL_226 = tile__EVAL_24;
  assign rsource__EVAL_46 = _EVAL_57;
  assign rsink__EVAL_31 = _EVAL_58;
  assign _EVAL_182 = _EVAL_238;
  assign _EVAL_81 = rsink__EVAL_5;
  assign _EVAL_255 = _EVAL_210;
  assign _EVAL_119 = _EVAL_196;
  assign _EVAL_160 = _EVAL_155;
  assign intsink_1__EVAL_0 = _EVAL_73;
  assign tile__EVAL_34 = _EVAL_204;
  assign _EVAL_209 = tile__EVAL_11;
  assign rsink__EVAL_1 = _EVAL_49;
  assign _EVAL_76 = rsource__EVAL_49;
  assign _EVAL_27 = rsource__EVAL_25;
  assign rsink__EVAL_20 = _EVAL_87;
  assign _EVAL_124 = _EVAL_188;
  assign tile__EVAL_61 = _EVAL_223;
  assign _EVAL_122 = intsink_3__EVAL_26;
  assign _EVAL_243 = _EVAL_253;
  assign rsource__EVAL_57 = _EVAL_10;
  assign _EVAL_51 = rsource__EVAL_62;
  assign _EVAL_12 = rsource__EVAL_21;
  assign tile__EVAL_68 = _EVAL_173;
  assign _EVAL_225 = rsource__EVAL_22;
  assign _EVAL_241 = tile__EVAL_4;
  assign _EVAL_151 = _EVAL_230;
  assign _EVAL_60 = rsource__EVAL_53;
  assign rsink__EVAL_16 = _EVAL_101;
  assign _EVAL_244 = _EVAL_206;
  assign _EVAL_11 = rsource__EVAL_2;
  assign tile__EVAL_20 = _EVAL_255;
  assign tile__EVAL_23 = _EVAL_213;
  assign _EVAL_133 = _EVAL_169;
  assign tile__EVAL_43 = _EVAL_122;
  assign _EVAL_240 = _EVAL_224;
  assign _EVAL_82 = rsink__EVAL_43;
  assign _EVAL_211 = _EVAL_180;
  assign tile__EVAL_60 = _EVAL_135;
  assign _EVAL_228 = intsink_3__EVAL_6;
  assign _EVAL_26 = rsource__EVAL_29;
  assign _EVAL_154 = _EVAL_121;
  assign _EVAL_206 = tile__EVAL_6;
  assign _EVAL_196 = _EVAL_242;
  assign _EVAL_170 = _EVAL_218;
  assign _EVAL_56 = rsource__EVAL_26;
  assign tile__EVAL_41 = _EVAL_215;
  assign tile__EVAL_66 = _EVAL_245;
  assign _EVAL_183 = rsink__EVAL_14;
  assign tile__EVAL_27 = _EVAL_189;
  assign _EVAL_224 = rsource__EVAL_7;
  assign _EVAL_144 = tile__EVAL_18;
  assign intsink_3__EVAL_16 = _EVAL_64;
  assign _EVAL_219 = _EVAL_167;
  assign tile__EVAL_67 = _EVAL_126;
  assign rsink__EVAL_19 = _EVAL_67;
  assign _EVAL_251 = intsink_3__EVAL_5;
  assign intsink_3__EVAL_24 = _EVAL_3;
  assign _EVAL_156 = tile__EVAL_35;
  assign _EVAL_210 = _EVAL_186;
  assign _EVAL_169 = tile__EVAL_44;
  assign _EVAL_223 = _EVAL_221;
  assign tile__EVAL_51 = _EVAL_202;
  assign _EVAL_238 = _EVAL_146;
  assign _EVAL_239 = tile__EVAL_10;
  assign tile__EVAL_31 = _EVAL_142;
  assign _EVAL_47 = rsource__EVAL_19;
  assign rsource__EVAL_5 = _EVAL_75;
  assign _EVAL_246 = _EVAL_132;
  assign _EVAL_127 = _EVAL_147;
  assign rsource__EVAL_66 = _EVAL_72;
  assign tile__EVAL_14 = _EVAL_154;
  assign _EVAL_34 = rsink__EVAL_40;
  assign rsource__EVAL_31 = _EVAL_95;
  assign intsink_3__EVAL_22 = _EVAL_52;
  assign _EVAL_163 = _EVAL_237;
  assign _EVAL_31 = rsource__EVAL_34;
  assign rsource__EVAL_10 = _EVAL_170;
  assign _EVAL_260 = intsink_3__EVAL_4;
  assign _EVAL_178 = tile__EVAL_47;
  assign _EVAL_215 = intsink_3__EVAL_28;
  assign _EVAL_98 = rsource__EVAL_59;
  assign _EVAL_204 = _EVAL_18;
  assign _EVAL_123 = tile__EVAL_45;
  assign intsink_2__EVAL_0 = _EVAL_48;
  assign rsink__EVAL_34 = _EVAL_243;
  assign _EVAL_139 = tile__EVAL_48;
  assign _EVAL_173 = intsink_3__EVAL_11;
  assign _EVAL_190 = tile__EVAL_38;
  assign intsink_1__EVAL_1 = _EVAL_95;
  assign rsink__EVAL_18 = _EVAL_48;
  assign rsink__EVAL_44 = _EVAL_259;
  assign _EVAL_259 = _EVAL_244;
  assign tile__EVAL_40 = _EVAL_251;
  assign rsource__EVAL_12 = _EVAL_151;
  assign tile__EVAL_32 = _EVAL_212;
  assign _EVAL_150 = intsink_3__EVAL_30;
  assign rsink__EVAL_2 = _EVAL_63;
  assign _EVAL_71 = rsink__EVAL_37;
  assign _EVAL_189 = intsink_3__EVAL_18;
  assign tile__EVAL_29 = _EVAL_153;
  assign tile__EVAL_1 = _EVAL_158;
  assign _EVAL_134 = tile__EVAL_52;
  assign intsink_3__EVAL_14 = _EVAL_93;
  assign rsink__EVAL_4 = _EVAL_136;
  assign _EVAL_191 = intsink_3__EVAL_13;
  assign tile__EVAL_8 = _EVAL_198;
  assign _EVAL_16 = rsource__EVAL_69;
  assign _EVAL_249 = _EVAL_125;
  assign _EVAL_231 = tile__EVAL_46;
  assign intsink_3__EVAL_7 = _EVAL_44;
  assign _EVAL_118 = _EVAL_144;
  assign intsink__EVAL_0 = _EVAL_1;
  assign _EVAL_202 = _EVAL_114;
  assign _EVAL_128 = _EVAL_177;
  assign _EVAL_108 = rsource__EVAL_39;
  assign intsink_1__EVAL = _EVAL_48;
  assign _EVAL_17 = rsource__EVAL_51;
  assign intsink_3__EVAL = _EVAL_53;
  assign rsource__EVAL = _EVAL_145;
  assign rsource__EVAL_42 = _EVAL_68;
  assign intsink_3__EVAL_29 = _EVAL_24;
  assign tile__EVAL_25 = _EVAL_248;
  assign rsource__EVAL_28 = _EVAL_78;
  assign _EVAL_157 = _EVAL_133;
  assign intsource_1__EVAL_0 = 1'h0;
  assign rsink__EVAL_25 = _EVAL_182;
  assign _EVAL_149 = _EVAL_148;
  assign tile__EVAL_56 = _EVAL_219;
  assign _EVAL_180 = rsink__EVAL_17;
  assign tile__EVAL_65 = _EVAL_149;
  assign intsink_1__EVAL_2 = _EVAL_61;
  assign _EVAL_214 = rsink__EVAL_3;
  assign _EVAL_179 = tile__EVAL_62;
  assign _EVAL_132 = _EVAL_201;
  assign rsink__EVAL_38 = _EVAL_86;
  assign _EVAL_54 = rsource__EVAL_44;
  assign _EVAL_140 = _EVAL_164;
  assign _EVAL_28 = intsource_4__EVAL;
  assign _EVAL_88 = rsource__EVAL_56;
  assign _EVAL_113 = _EVAL_161;
  assign _EVAL_230 = _EVAL_139;
  assign _EVAL_250 = _EVAL_176;
  assign _EVAL_126 = intsink_3__EVAL_20;
  assign rsource__EVAL_30 = _EVAL_48;
  assign _EVAL_15 = rsink__EVAL_42;
  assign _EVAL_256 = _EVAL_179;
  assign _EVAL_220 = _EVAL_128;
  assign _EVAL_138 = _EVAL_9;
  assign tile__EVAL_19 = _EVAL_119;
  assign tile__EVAL_17 = _EVAL_165;
  assign tile__EVAL_28 = _EVAL_141;
  assign _EVAL_177 = rsource__EVAL_9;
  assign tile__EVAL_33 = _EVAL_192;
  assign rsource__EVAL_8 = _EVAL_83;
  assign _EVAL_153 = _EVAL_140;
  assign _EVAL_115 = _EVAL_208;
  assign _EVAL_167 = _EVAL_233;
  assign rsource__EVAL_64 = _EVAL_21;
  assign _EVAL_164 = rsource__EVAL_58;
  assign rsource__EVAL_41 = _EVAL_216;
  assign intsink_3__EVAL_3 = _EVAL_43;
  assign _EVAL_235 = _EVAL_124;
  assign _EVAL_195 = rsource__EVAL_71;
  assign _EVAL_110 = _EVAL_199;
  assign rsource__EVAL_16 = _EVAL_0;
  assign _EVAL_192 = intsink_2__EVAL_2;
  assign tile__EVAL_59 = _EVAL_200;
  assign _EVAL_227 = _EVAL_131;
  assign _EVAL_242 = rsource__EVAL_6;
  assign _EVAL_199 = _EVAL_214;
  assign _EVAL_234 = _EVAL_209;
  assign _EVAL_247 = _EVAL_29;
  assign _EVAL_208 = rsink__EVAL_41;
  assign rsource__EVAL_15 = _EVAL_103;
  assign rsource__EVAL_33 = _EVAL_89;
  assign tile__EVAL_26 = _EVAL_111;
  assign _EVAL_213 = _EVAL_115;
  assign rsource__EVAL_47 = _EVAL_94;
  assign _EVAL_217 = _EVAL_36;
  assign rsource__EVAL_27 = _EVAL_59;
  assign _EVAL_252 = _EVAL_256;
  assign rsource__EVAL_68 = _EVAL_235;
  assign _EVAL_105 = rsink__EVAL_6;
  assign _EVAL_258 = _EVAL_109;
  assign tile__EVAL_15 = _EVAL_162;
  assign intsink_3__EVAL_15 = _EVAL_85;
  assign _EVAL_146 = tile__EVAL_39;
  assign rsink__EVAL_35 = _EVAL_2;
  assign _EVAL_193 = _EVAL_118;
  assign _EVAL_96 = intsource_3__EVAL;
  assign rsink__EVAL_0 = _EVAL_227;
  assign intsink_3__EVAL_1 = _EVAL_6;
  assign intsink_2__EVAL = _EVAL_77;
  assign _EVAL_62 = rsink__EVAL_11;
  assign _EVAL_236 = _EVAL_258;
  assign tile__EVAL_36 = _EVAL_247;
  assign _EVAL_42 = rsource__EVAL_65;
  assign _EVAL_221 = _EVAL_225;
  assign _EVAL_176 = _EVAL_239;
  assign tile__EVAL_9 = _EVAL_150;
  assign rsink__EVAL_12 = _EVAL_14;
  assign rsource__EVAL_72 = _EVAL_65;
  assign _EVAL_129 = tile__EVAL_55;
  assign _EVAL_253 = _EVAL_190;
  assign _EVAL_92 = rsink__EVAL_7;
  assign _EVAL_229 = tile__EVAL_16;
  assign rsource__EVAL_3 = _EVAL_102;
  assign rsink__EVAL_23 = _EVAL_106;
  assign _EVAL_162 = _EVAL_222;
  assign _EVAL_168 = intsink_3__EVAL_19;
  assign tile__EVAL_2 = _EVAL_175;
  assign _EVAL_248 = intsink__EVAL;
  assign tile__EVAL_49 = _EVAL_168;
  assign _EVAL_45 = rsource__EVAL_36;
  assign _EVAL_99 = rsource__EVAL_14;
  assign _EVAL_232 = _EVAL_181;
  assign intsink_3__EVAL_12 = _EVAL_39;
  assign rsource__EVAL_35 = _EVAL_250;
  assign intsink_3__EVAL_21 = _EVAL_74;
  assign rsink__EVAL_33 = _EVAL_66;
  assign _EVAL_233 = rsink__EVAL_24;
  assign _EVAL_116 = _EVAL_197;
  assign _EVAL_165 = intsink_3__EVAL_17;
  assign tile__EVAL_64 = _EVAL_171;
  assign _EVAL_5 = rsink__EVAL_9;
  assign intsink_3__EVAL_23 = _EVAL_4;
  assign tile__EVAL_53 = _EVAL_116;
  assign intsink_3__EVAL_27 = _EVAL_107;
  assign rsink__EVAL_39 = _EVAL_40;
  assign _EVAL_218 = _EVAL_231;
  assign rsink__EVAL = _EVAL_23;
  assign _EVAL_197 = _EVAL_152;
  assign rsink__EVAL_15 = _EVAL_95;
  assign _EVAL_114 = _EVAL_143;
  assign _EVAL_203 = rsink__EVAL_8;
  assign rsource__EVAL_37 = _EVAL_8;
  assign _EVAL_171 = intsink_3__EVAL_0;
  assign rsource__EVAL_32 = _EVAL_246;
  assign _EVAL_181 = rsink__EVAL_21;
endmodule
