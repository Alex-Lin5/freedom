//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_177_assert(
  input          _EVAL,
  input          _EVAL_1,
  input  [2:0]   _EVAL_3,
  input  [9:0]   _EVAL_6,
  input  [2:0]   _EVAL_9,
  input          _EVAL_14,
  input          _EVAL_17,
  input          _EVAL_19,
  input  [2:0]   _EVAL_26,
  input  [2:0]   _EVAL_27,
  input          _EVAL_30,
  input          _EVAL_31,
  input  [3:0]   _EVAL_32,
  input  [1:0]   _EVAL_33,
  input          _EVAL_36,
  input  [8:0]   _EVAL_42,
  input  [3:0]   _EVAL_43,
  input  [1:0]   _EVAL_49,
  input          _EVAL_51,
  input  [11:0]  _EVAL_54,
  input          _EVAL_63,
  input          _EVAL_72,
  input          _EVAL_84,
  input          _EVAL_92,
  input          _EVAL_96,
  input          _EVAL_98,
  input          _EVAL_107,
  input          _EVAL_109,
  input          _EVAL_117,
  input          _EVAL_122,
  input          _EVAL_125,
  input          _EVAL_135,
  input          _EVAL_154,
  input          _EVAL_169,
  input          _EVAL_211,
  input          _EVAL_216,
  input          _EVAL_219,
  input          _EVAL_227,
  input          _EVAL_228,
  input          _EVAL_248,
  input          _EVAL_261,
  input          _EVAL_270,
  input          _EVAL_310,
  input          _EVAL_317,
  input          _EVAL_337,
  input          _EVAL_340,
  input          _EVAL_346,
  input          _EVAL_356,
  input          _EVAL_366,
  input          _EVAL_367,
  input          _EVAL_369,
  input          _EVAL_385,
  input          _EVAL_386,
  input          _EVAL_389,
  input          _EVAL_393,
  input          _EVAL_395,
  input          _EVAL_407,
  input          _EVAL_416,
  input          _EVAL_419,
  input          _EVAL_426,
  input          _EVAL_427,
  input          _EVAL_438,
  input          _EVAL_439,
  input          _EVAL_443,
  input          _EVAL_449,
  input          _EVAL_454,
  input          _EVAL_460,
  input          _EVAL_462,
  input          _EVAL_472,
  input  [2:0]   _EVAL_475,
  input          _EVAL_479,
  input          _EVAL_491,
  input          _EVAL_497,
  input          _EVAL_505,
  input          _EVAL_511,
  input          _EVAL_519,
  input          _EVAL_522,
  input          _EVAL_523,
  input          _EVAL_549,
  input          _EVAL_552,
  input  [7:0]   _EVAL_554,
  input          _EVAL_556,
  input          _EVAL_561,
  input          _EVAL_567,
  input          _EVAL_572,
  input          _EVAL_577,
  input  [63:0]  _EVAL_586,
  input          _EVAL_592,
  input          _EVAL_597,
  input          _EVAL_607,
  input          _EVAL_613,
  input          _EVAL_614,
  input          _EVAL_623,
  input          _EVAL_629,
  input          _EVAL_635,
  input          _EVAL_638,
  input          _EVAL_639,
  input          _EVAL_643,
  input          _EVAL_648,
  input          _EVAL_658,
  input          _EVAL_666,
  input          _EVAL_685,
  input          _EVAL_687,
  input          _EVAL_691,
  input          _EVAL_694,
  input          _EVAL_705,
  input          _EVAL_707,
  input  [2:0]   _EVAL_723,
  input          _EVAL_725,
  input          _EVAL_726,
  input          _EVAL_747,
  input          _EVAL_763,
  input  [7:0]   _EVAL_765,
  input          _EVAL_766,
  input          _EVAL_778,
  input          _EVAL_784,
  input          _EVAL_788,
  input          _EVAL_801,
  input          _EVAL_811,
  input          _EVAL_813,
  input          _EVAL_821,
  input          _EVAL_823,
  input          _EVAL_825,
  input          _EVAL_831,
  input          _EVAL_837,
  input          _EVAL_842,
  input          _EVAL_848,
  input          _EVAL_849,
  input          _EVAL_858,
  input          _EVAL_859,
  input          _EVAL_861,
  input          _EVAL_866,
  input          _EVAL_871,
  input          _EVAL_883,
  input          _EVAL_888,
  input          _EVAL_890,
  input          _EVAL_895,
  input          _EVAL_898,
  input          _EVAL_904,
  input          _EVAL_907,
  input          _EVAL_914,
  input          _EVAL_924,
  input          _EVAL_929,
  input  [7:0]   _EVAL_949,
  input          _EVAL_951,
  input          _EVAL_959,
  input          _EVAL_961,
  input          _EVAL_963,
  input          _EVAL_973,
  input          _EVAL_976,
  input          _EVAL_984,
  input          _EVAL_1002,
  input          _EVAL_1022,
  input          _EVAL_1023,
  input          _EVAL_1026,
  input          _EVAL_1028,
  input          _EVAL_1038,
  input          _EVAL_1043,
  input          _EVAL_1047,
  input          _EVAL_1059,
  input          _EVAL_1061,
  input          _EVAL_1070,
  input          _EVAL_1083,
  input          _EVAL_1086,
  input  [1:0]   _EVAL_1096,
  input          _EVAL_1099,
  input          _EVAL_1105,
  input          _EVAL_1109,
  input          _EVAL_1112,
  input          _EVAL_1129,
  input          _EVAL_1138,
  input          _EVAL_1148,
  input          _EVAL_1159,
  input          _EVAL_1160,
  input          _EVAL_1162,
  input          _EVAL_1185,
  input          _EVAL_1203,
  input          _EVAL_1207,
  input          _EVAL_1227,
  input          _EVAL_1236,
  input          _EVAL_1239,
  input          _EVAL_1245,
  input          _EVAL_1247,
  input          _EVAL_1255,
  input          _EVAL_1264,
  input          _EVAL_1267,
  input          _EVAL_1271,
  input          _EVAL_1278,
  input          _EVAL_1280,
  input  [2:0]   _EVAL_1285,
  input          _EVAL_1289,
  input          _EVAL_1290,
  input          _EVAL_1305,
  input          _EVAL_1311,
  input          _EVAL_1317,
  input          _EVAL_1321,
  input          _EVAL_1325,
  input          _EVAL_1326,
  input          _EVAL_1327,
  input          _EVAL_1331,
  input  [511:0] _EVAL_1333,
  input          _EVAL_1338,
  input          _EVAL_1342,
  input          _EVAL_1343,
  input          _EVAL_1348,
  input          _EVAL_1350,
  input          _EVAL_1359,
  input          _EVAL_1364,
  input          _EVAL_1367,
  input          _EVAL_1368,
  input          _EVAL_1375,
  input          _EVAL_1379,
  input          _EVAL_1381,
  input          _EVAL_1396,
  input          _EVAL_1409,
  input          _EVAL_1410,
  input          _EVAL_1411,
  input          _EVAL_1422,
  input          _EVAL_1431,
  input          _EVAL_1445,
  input          _EVAL_1448,
  input          _EVAL_1452,
  input          _EVAL_1463,
  input          _EVAL_1475,
  input          _EVAL_1485,
  input          _EVAL_1498,
  input  [31:0]  _EVAL_1502,
  input          _EVAL_1505,
  input          _EVAL_1516,
  input          _EVAL_1527,
  input          _EVAL_1532,
  input          _EVAL_1534,
  input          _EVAL_1537,
  input          _EVAL_1539,
  input          _EVAL_1545,
  input          _EVAL_1552,
  input          _EVAL_1559,
  input          _EVAL_1568,
  input          _EVAL_1575,
  input          _EVAL_1583,
  input          _EVAL_1596,
  input          _EVAL_1613,
  input          _EVAL_1615,
  input          _EVAL_1640,
  input          _EVAL_1646,
  input          _EVAL_1648,
  input          _EVAL_1658,
  input          _EVAL_1683,
  input  [2:0]   _EVAL_1704,
  input          _EVAL_1707,
  input          _EVAL_1714,
  input  [7:0]   _EVAL_1716,
  input          _EVAL_1726,
  input          _EVAL_1730,
  input          _EVAL_1731,
  input          _EVAL_1744,
  input          _EVAL_1757,
  input          _EVAL_1763,
  input  [15:0]  _EVAL_1775,
  input          _EVAL_1785,
  input          _EVAL_1791,
  input          _EVAL_1792,
  input          _EVAL_1794,
  input          _EVAL_1795,
  input          _EVAL_1805,
  input  [31:0]  _EVAL_1815,
  input          _EVAL_1824,
  input          _EVAL_1834,
  input          _EVAL_1837,
  input          _EVAL_1841,
  input          _EVAL_1850,
  input          _EVAL_1852,
  input          _EVAL_1858,
  input          _EVAL_1859,
  input          _EVAL_1869,
  input          _EVAL_1875,
  input          _EVAL_1876,
  input          _EVAL_1880,
  input          _EVAL_1898,
  input          _EVAL_1904,
  input          _EVAL_1906,
  input          _EVAL_1909,
  input          _EVAL_1925,
  input          _EVAL_1946,
  input          _EVAL_1957,
  input          _EVAL_1958,
  input          _EVAL_1977,
  input          _EVAL_1985,
  input          _EVAL_1987,
  input          _EVAL_1988,
  input          _EVAL_1992,
  input          _EVAL_1996,
  input          _EVAL_2003,
  input          _EVAL_2015,
  input          _EVAL_2017,
  input          _EVAL_2018,
  input          _EVAL_2028,
  input          _EVAL_2031,
  input          _EVAL_2033,
  input          _EVAL_2035,
  input          _EVAL_2037,
  input          _EVAL_2039,
  input          _EVAL_2041,
  input          _EVAL_2043,
  input          _EVAL_2045,
  input          _EVAL_2047,
  input          _EVAL_2052,
  input          sb2tlOpt__EVAL_27,
  input          sb2tlOpt__EVAL_12
);
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_82;
  wire  _EVAL_85;
  wire  _EVAL_88;
  wire  _EVAL_91;
  wire  _EVAL_93;
  wire  _EVAL_95;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_106;
  wire  _EVAL_110;
  wire  _EVAL_113;
  wire  _EVAL_119;
  wire  _EVAL_123;
  wire  _EVAL_136;
  wire  _EVAL_138;
  wire  _EVAL_142;
  wire  _EVAL_149;
  wire  _EVAL_151;
  wire  _EVAL_153;
  wire  _EVAL_157;
  wire  _EVAL_160;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_175;
  wire  _EVAL_179;
  wire  _EVAL_181;
  wire  _EVAL_183;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_197;
  wire  _EVAL_201;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_214;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_224;
  wire  _EVAL_232;
  wire  _EVAL_236;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_260;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_277;
  wire  _EVAL_279;
  wire  _EVAL_292;
  wire  _EVAL_294;
  wire  _EVAL_303;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_318;
  wire  _EVAL_320;
  wire  _EVAL_324;
  wire  _EVAL_329;
  wire  _EVAL_330;
  wire  _EVAL_338;
  wire  _EVAL_365;
  wire  _EVAL_368;
  wire  _EVAL_370;
  wire  _EVAL_371;
  wire  _EVAL_378;
  wire  _EVAL_381;
  wire  _EVAL_387;
  wire  _EVAL_394;
  wire  _EVAL_398;
  wire  _EVAL_401;
  wire  _EVAL_402;
  wire  _EVAL_404;
  wire  _EVAL_405;
  wire  _EVAL_406;
  wire  _EVAL_409;
  wire  _EVAL_414;
  wire  _EVAL_424;
  wire  _EVAL_440;
  wire  _EVAL_442;
  wire  _EVAL_452;
  wire  _EVAL_459;
  wire  _EVAL_461;
  wire  _EVAL_468;
  wire  _EVAL_469;
  wire  _EVAL_477;
  wire  _EVAL_483;
  wire  _EVAL_488;
  wire  _EVAL_489;
  wire  _EVAL_492;
  wire  _EVAL_495;
  wire  _EVAL_509;
  wire  _EVAL_512;
  wire  _EVAL_514;
  wire  _EVAL_518;
  wire  _EVAL_524;
  wire  _EVAL_527;
  wire  _EVAL_533;
  wire  _EVAL_539;
  wire  _EVAL_547;
  wire  _EVAL_551;
  wire  _EVAL_558;
  wire  _EVAL_571;
  wire  _EVAL_573;
  wire  _EVAL_579;
  wire  _EVAL_580;
  wire  _EVAL_581;
  wire  _EVAL_583;
  wire  _EVAL_584;
  wire  _EVAL_588;
  wire  _EVAL_596;
  wire [3:0] _EVAL_599;
  wire  _EVAL_602;
  wire  _EVAL_612;
  wire  _EVAL_615;
  wire  _EVAL_616;
  wire  _EVAL_619;
  wire  _EVAL_622;
  wire  _EVAL_627;
  wire  _EVAL_630;
  wire  _EVAL_633;
  wire  _EVAL_637;
  wire  _EVAL_645;
  wire  _EVAL_646;
  wire  _EVAL_656;
  wire  _EVAL_659;
  wire  _EVAL_662;
  wire [2:0] _EVAL_663;
  wire  _EVAL_672;
  wire  _EVAL_679;
  wire  _EVAL_681;
  wire  _EVAL_682;
  wire  _EVAL_683;
  wire  _EVAL_693;
  wire  _EVAL_695;
  wire  _EVAL_697;
  wire  _EVAL_703;
  wire  _EVAL_706;
  wire  _EVAL_711;
  wire  _EVAL_719;
  wire  _EVAL_720;
  wire  _EVAL_721;
  wire  _EVAL_730;
  wire  _EVAL_731;
  wire  _EVAL_734;
  wire  _EVAL_738;
  wire  _EVAL_746;
  wire  _EVAL_750;
  wire  _EVAL_752;
  wire  _EVAL_759;
  wire  _EVAL_762;
  wire  _EVAL_764;
  wire  _EVAL_770;
  wire  _EVAL_771;
  wire  _EVAL_774;
  wire  _EVAL_780;
  wire  _EVAL_792;
  wire  _EVAL_796;
  wire  _EVAL_798;
  wire  _EVAL_800;
  wire  _EVAL_804;
  wire  _EVAL_806;
  wire  _EVAL_808;
  wire  _EVAL_809;
  wire [2:0] monitor_1__EVAL;
  wire  monitor_1__EVAL_0;
  wire  monitor_1__EVAL_1;
  wire [9:0] monitor_1__EVAL_2;
  wire [1:0] monitor_1__EVAL_3;
  wire [11:0] monitor_1__EVAL_4;
  wire  monitor_1__EVAL_5;
  wire  monitor_1__EVAL_6;
  wire [2:0] monitor_1__EVAL_7;
  wire [1:0] monitor_1__EVAL_8;
  wire [9:0] monitor_1__EVAL_9;
  wire  monitor_1__EVAL_10;
  wire  monitor_1__EVAL_11;
  wire [2:0] monitor_1__EVAL_12;
  wire  monitor_1__EVAL_13;
  wire [3:0] monitor_1__EVAL_14;
  wire [14:0] _EVAL_816;
  wire  _EVAL_824;
  wire  _EVAL_826;
  wire  _EVAL_835;
  wire  _EVAL_843;
  wire  _EVAL_853;
  wire  _EVAL_864;
  wire  _EVAL_872;
  wire  _EVAL_873;
  wire  _EVAL_878;
  wire  _EVAL_879;
  wire  _EVAL_889;
  wire  _EVAL_893;
  wire  _EVAL_909;
  wire  _EVAL_913;
  wire  _EVAL_917;
  wire  _EVAL_918;
  wire  _EVAL_919;
  wire  _EVAL_930;
  wire  _EVAL_932;
  wire  _EVAL_938;
  wire  _EVAL_944;
  wire  _EVAL_947;
  wire  _EVAL_948;
  wire [2:0] monitor__EVAL;
  wire  monitor__EVAL_0;
  wire [1:0] monitor__EVAL_1;
  wire [2:0] monitor__EVAL_2;
  wire [8:0] monitor__EVAL_3;
  wire  monitor__EVAL_4;
  wire  monitor__EVAL_5;
  wire  monitor__EVAL_6;
  wire  monitor__EVAL_7;
  wire  monitor__EVAL_8;
  wire  monitor__EVAL_9;
  wire  monitor__EVAL_10;
  wire [1:0] monitor__EVAL_11;
  wire [2:0] monitor__EVAL_12;
  wire [3:0] monitor__EVAL_13;
  wire  monitor__EVAL_14;
  wire  _EVAL_953;
  wire  _EVAL_955;
  wire  _EVAL_962;
  wire  _EVAL_965;
  wire  _EVAL_970;
  wire  _EVAL_977;
  wire  _EVAL_983;
  wire  _EVAL_985;
  wire  _EVAL_990;
  wire  _EVAL_993;
  wire  _EVAL_997;
  wire  _EVAL_1003;
  wire  _EVAL_1005;
  wire  _EVAL_1006;
  wire  _EVAL_1034;
  wire  _EVAL_1037;
  wire  _EVAL_1039;
  wire  _EVAL_1041;
  wire  _EVAL_1060;
  wire  _EVAL_1064;
  wire  _EVAL_1065;
  wire  _EVAL_1066;
  wire  _EVAL_1076;
  wire  _EVAL_1082;
  wire  _EVAL_1093;
  wire  _EVAL_1095;
  wire  _EVAL_1098;
  wire  _EVAL_1100;
  wire  _EVAL_1103;
  wire  _EVAL_1106;
  wire  _EVAL_1110;
  wire  _EVAL_1115;
  wire  _EVAL_1117;
  wire  _EVAL_1120;
  wire  _EVAL_1121;
  wire  _EVAL_1122;
  wire  _EVAL_1135;
  wire  _EVAL_1137;
  wire  _EVAL_1143;
  wire  _EVAL_1145;
  wire [3:0] _EVAL_1152;
  wire  _EVAL_1157;
  wire  _EVAL_1165;
  wire  _EVAL_1170;
  wire  _EVAL_1172;
  wire  _EVAL_1174;
  wire  _EVAL_1182;
  wire  _EVAL_1190;
  wire  _EVAL_1194;
  wire  _EVAL_1198;
  wire  _EVAL_1205;
  wire  _EVAL_1214;
  wire  _EVAL_1218;
  wire  _EVAL_1221;
  wire  _EVAL_1225;
  wire  _EVAL_1228;
  wire  _EVAL_1235;
  wire  _EVAL_1237;
  wire  _EVAL_1246;
  wire  _EVAL_1250;
  wire  _EVAL_1258;
  wire  _EVAL_1259;
  wire  _EVAL_1266;
  wire  _EVAL_1270;
  wire  _EVAL_1277;
  wire  _EVAL_1287;
  wire  _EVAL_1291;
  wire  _EVAL_1292;
  wire  _EVAL_1293;
  wire  _EVAL_1299;
  wire  _EVAL_1308;
  wire  _EVAL_1319;
  wire  _EVAL_1320;
  wire  _EVAL_1330;
  wire  _EVAL_1332;
  wire  _EVAL_1341;
  wire  _EVAL_1344;
  wire  _EVAL_1351;
  wire  _EVAL_1354;
  wire  _EVAL_1357;
  wire  _EVAL_1360;
  wire  _EVAL_1366;
  wire  _EVAL_1377;
  wire  _EVAL_1382;
  wire  _EVAL_1383;
  wire  _EVAL_1393;
  wire  _EVAL_1395;
  wire  _EVAL_1397;
  wire [1:0] _EVAL_1398;
  wire  _EVAL_1401;
  wire  _EVAL_1402;
  wire  _EVAL_1413;
  wire  _EVAL_1424;
  wire  _EVAL_1429;
  wire  _EVAL_1430;
  wire  _EVAL_1433;
  wire  _EVAL_1434;
  wire  _EVAL_1436;
  wire  _EVAL_1444;
  wire  _EVAL_1456;
  wire  _EVAL_1457;
  wire  _EVAL_1462;
  wire  _EVAL_1469;
  wire  _EVAL_1470;
  wire  _EVAL_1476;
  wire  _EVAL_1478;
  wire  _EVAL_1481;
  wire  _EVAL_1484;
  wire  _EVAL_1487;
  wire  _EVAL_1491;
  wire [4:0] _EVAL_1492;
  wire  _EVAL_1493;
  wire  _EVAL_1494;
  wire  _EVAL_1495;
  wire  _EVAL_1496;
  wire  _EVAL_1499;
  wire [10:0] _EVAL_1500;
  wire  _EVAL_1508;
  wire  _EVAL_1510;
  wire  _EVAL_1511;
  wire  _EVAL_1512;
  wire  _EVAL_1514;
  wire  _EVAL_1517;
  wire  _EVAL_1521;
  wire  _EVAL_1523;
  wire  _EVAL_1528;
  wire  _EVAL_1531;
  wire  _EVAL_1535;
  wire  _EVAL_1538;
  wire  _EVAL_1550;
  wire  _EVAL_1551;
  wire  _EVAL_1554;
  wire  _EVAL_1564;
  wire  _EVAL_1570;
  wire  _EVAL_1573;
  wire  _EVAL_1585;
  wire  _EVAL_1589;
  wire  _EVAL_1597;
  wire [6:0] _EVAL_1598;
  wire  _EVAL_1602;
  wire  _EVAL_1608;
  wire  _EVAL_1609;
  wire  _EVAL_1621;
  wire  _EVAL_1622;
  wire  _EVAL_1624;
  wire  _EVAL_1625;
  wire  _EVAL_1626;
  wire  _EVAL_1628;
  wire  _EVAL_1630;
  wire  _EVAL_1631;
  wire  _EVAL_1645;
  wire  _EVAL_1647;
  wire  _EVAL_1649;
  wire  _EVAL_1651;
  wire  _EVAL_1654;
  wire  _EVAL_1655;
  wire  _EVAL_1656;
  wire  _EVAL_1661;
  wire  _EVAL_1662;
  wire  _EVAL_1665;
  wire  _EVAL_1668;
  wire  _EVAL_1670;
  wire  _EVAL_1671;
  wire [1:0] _EVAL_1673;
  wire  _EVAL_1674;
  wire  _EVAL_1676;
  wire  _EVAL_1680;
  wire  _EVAL_1684;
  wire  _EVAL_1686;
  wire  _EVAL_1695;
  wire  _EVAL_1696;
  wire  _EVAL_1699;
  wire  _EVAL_1709;
  wire  _EVAL_1725;
  wire  _EVAL_1727;
  wire  _EVAL_1734;
  wire  _EVAL_1736;
  wire  _EVAL_1739;
  wire  _EVAL_1741;
  wire  _EVAL_1746;
  wire  _EVAL_1747;
  wire  _EVAL_1750;
  wire  _EVAL_1764;
  wire [5:0] _EVAL_1766;
  wire  _EVAL_1771;
  wire  _EVAL_1777;
  wire  _EVAL_1780;
  wire  _EVAL_1788;
  wire  _EVAL_1797;
  wire  _EVAL_1799;
  wire  _EVAL_1802;
  wire  _EVAL_1806;
  wire  _EVAL_1809;
  wire  _EVAL_1810;
  wire  _EVAL_1818;
  wire  _EVAL_1820;
  wire  _EVAL_1821;
  wire  _EVAL_1822;
  wire  _EVAL_1825;
  wire  _EVAL_1829;
  wire  _EVAL_1831;
  wire  _EVAL_1838;
  wire  _EVAL_1840;
  wire  _EVAL_1842;
  wire  _EVAL_1854;
  wire  _EVAL_1855;
  wire  _EVAL_1856;
  wire  _EVAL_1862;
  wire  _EVAL_1870;
  wire  _EVAL_1871;
  wire  _EVAL_1878;
  wire  _EVAL_1879;
  wire  _EVAL_1883;
  wire  _EVAL_1890;
  wire  _EVAL_1892;
  wire  _EVAL_1893;
  wire  _EVAL_1896;
  wire  _EVAL_1899;
  wire  _EVAL_1902;
  wire  _EVAL_1911;
  wire  _EVAL_1916;
  wire  _EVAL_1924;
  wire  _EVAL_1926;
  wire  _EVAL_1930;
  wire  _EVAL_1938;
  wire  _EVAL_1939;
  wire  _EVAL_1947;
  wire  _EVAL_1952;
  wire  _EVAL_1955;
  wire  _EVAL_1960;
  wire  _EVAL_1963;
  wire  _EVAL_1967;
  wire  _EVAL_1968;
  wire  _EVAL_1981;
  wire  _EVAL_1990;
  wire  _EVAL_2010;
  wire  _EVAL_2012;
  wire  _EVAL_2013;
  wire  _EVAL_2016;
  wire  _EVAL_2021;
  wire  _EVAL_2022;
  wire  _EVAL_2024;
  wire  _EVAL_2026;
  wire  _EVAL_2029;
  wire  _EVAL_2038;
  wire  _EVAL_2048;
  wire  _EVAL_2053;
  _EVAL_175_assert monitor_1 (
    ._EVAL(monitor_1__EVAL),
    ._EVAL_0(monitor_1__EVAL_0),
    ._EVAL_1(monitor_1__EVAL_1),
    ._EVAL_2(monitor_1__EVAL_2),
    ._EVAL_3(monitor_1__EVAL_3),
    ._EVAL_4(monitor_1__EVAL_4),
    ._EVAL_5(monitor_1__EVAL_5),
    ._EVAL_6(monitor_1__EVAL_6),
    ._EVAL_7(monitor_1__EVAL_7),
    ._EVAL_8(monitor_1__EVAL_8),
    ._EVAL_9(monitor_1__EVAL_9),
    ._EVAL_10(monitor_1__EVAL_10),
    ._EVAL_11(monitor_1__EVAL_11),
    ._EVAL_12(monitor_1__EVAL_12),
    ._EVAL_13(monitor_1__EVAL_13),
    ._EVAL_14(monitor_1__EVAL_14)
  );
  _EVAL_174_assert monitor (
    ._EVAL(monitor__EVAL),
    ._EVAL_0(monitor__EVAL_0),
    ._EVAL_1(monitor__EVAL_1),
    ._EVAL_2(monitor__EVAL_2),
    ._EVAL_3(monitor__EVAL_3),
    ._EVAL_4(monitor__EVAL_4),
    ._EVAL_5(monitor__EVAL_5),
    ._EVAL_6(monitor__EVAL_6),
    ._EVAL_7(monitor__EVAL_7),
    ._EVAL_8(monitor__EVAL_8),
    ._EVAL_9(monitor__EVAL_9),
    ._EVAL_10(monitor__EVAL_10),
    ._EVAL_11(monitor__EVAL_11),
    ._EVAL_12(monitor__EVAL_12),
    ._EVAL_13(monitor__EVAL_13),
    ._EVAL_14(monitor__EVAL_14)
  );
  assign _EVAL_1829 = _EVAL_1499 & _EVAL_236;
  assign _EVAL_809 = _EVAL_1330 & _EVAL_268;
  assign _EVAL_746 = _EVAL_100 & _EVAL_959;
  assign _EVAL_1246 = _EVAL_1499 & _EVAL_214;
  assign _EVAL_1528 = _EVAL_1499 & _EVAL_1514;
  assign _EVAL_1341 = |_EVAL_153;
  assign _EVAL_85 = _EVAL_1673 == 2'h3;
  assign _EVAL_990 = _EVAL_1270 & _EVAL_858;
  assign _EVAL_938 = _EVAL_1899 & _EVAL_442;
  assign monitor__EVAL = _EVAL_26;
  assign _EVAL_1492 = _EVAL_1502[28:24];
  assign _EVAL_91 = _EVAL_878 & _EVAL_442;
  assign _EVAL_1137 = _EVAL_1462 & _EVAL_1780;
  assign _EVAL_1398 = _EVAL_1502[21:20];
  assign _EVAL_101 = _EVAL_1484 & _EVAL_367;
  assign _EVAL_1862 = _EVAL_378 & _EVAL_1086;
  assign _EVAL_1060 = _EVAL_878 & _EVAL_1121;
  assign _EVAL_1695 = _EVAL_1499 & _EVAL_356;
  assign _EVAL_1430 = _EVAL_1172 & _EVAL_1121;
  assign _EVAL_800 = _EVAL_1821 & _EVAL_1174;
  assign _EVAL_1402 = |_EVAL_1955;
  assign _EVAL_1291 = _EVAL_1499 & _EVAL_1626;
  assign _EVAL_697 = _EVAL_1436 & _EVAL_442;
  assign monitor_1__EVAL_3 = _EVAL_49;
  assign _EVAL_1855 = _EVAL_1109 | _EVAL_533;
  assign _EVAL_279 = _EVAL_1502[9];
  assign _EVAL_1630 = _EVAL_637 & _EVAL_442;
  assign _EVAL_82 = _EVAL_1499 & _EVAL_924;
  assign _EVAL_633 = _EVAL_1292 & _EVAL_959;
  assign _EVAL_2022 = _EVAL_370 & _EVAL_1741;
  assign _EVAL_1822 = _EVAL_826 & _EVAL_320;
  assign _EVAL_1709 = _EVAL_1429 & _EVAL_1121;
  assign _EVAL_1628 = _EVAL_1165 & _EVAL_442;
  assign _EVAL_269 = _EVAL_1499 & _EVAL_1003;
  assign _EVAL_440 = _EVAL_1436 & _EVAL_1741;
  assign _EVAL_1508 = _EVAL_1333[274];
  assign _EVAL_917 = _EVAL_596 & _EVAL_959;
  assign _EVAL_1680 = |_EVAL_2016;
  assign _EVAL_1809 = _EVAL_164 & _EVAL_1121;
  assign _EVAL_62 = _EVAL_1499 & _EVAL_317;
  assign _EVAL_770 = _EVAL_1305 & _EVAL_385;
  assign _EVAL_759 = ~_EVAL_165;
  assign _EVAL_1512 = _EVAL_1165 & _EVAL_1741;
  assign _EVAL_993 = _EVAL_1333[264];
  assign _EVAL_1538 = _EVAL_1481 & _EVAL_1121;
  assign _EVAL_1899 = _EVAL_1893 & _EVAL_959;
  assign _EVAL_268 = ~_EVAL_2015;
  assign _EVAL_985 = |_EVAL_816;
  assign _EVAL_368 = _EVAL_1952 & _EVAL_117;
  assign _EVAL_948 = |_EVAL_489;
  assign _EVAL_277 = _EVAL_1198 & _EVAL_959;
  assign _EVAL_730 = |_EVAL_813;
  assign _EVAL_970 = _EVAL_1499 & _EVAL_1239;
  assign _EVAL_738 = _EVAL_1499 & _EVAL_1939;
  assign _EVAL_1115 = _EVAL_806 & _EVAL_442;
  assign monitor__EVAL_5 = _EVAL_17;
  assign _EVAL_1696 = _EVAL_277 & _EVAL_1121;
  assign _EVAL_1602 = _EVAL_113 & _EVAL_393;
  assign _EVAL_1496 = _EVAL_1190 & _EVAL_442;
  assign _EVAL_1082 = _EVAL_1902 & _EVAL_959;
  assign _EVAL_99 = _EVAL_1899 & _EVAL_1780;
  assign _EVAL_414 = _EVAL_1746 & _EVAL_1741;
  assign monitor__EVAL_7 = _EVAL_36;
  assign _EVAL_381 = _EVAL_1333[266];
  assign monitor_1__EVAL_11 = _EVAL_1;
  assign _EVAL_1621 = _EVAL_917 & _EVAL_1741;
  assign _EVAL_138 = _EVAL_221 & _EVAL_1780;
  assign _EVAL_853 = _EVAL_1535 & _EVAL_1741;
  assign _EVAL_1676 = _EVAL_1674 & _EVAL_197;
  assign _EVAL_1780 = |_EVAL_765;
  assign _EVAL_1939 = _EVAL_1333[270];
  assign _EVAL_77 = _EVAL_1499 & _EVAL_524;
  assign _EVAL_965 = _EVAL_1564 & _EVAL_442;
  assign _EVAL_1842 = _EVAL_78 & _EVAL_1086;
  assign _EVAL_201 = _EVAL_1797 & _EVAL_519;
  assign _EVAL_1727 = _EVAL_518 & _EVAL_117;
  assign _EVAL_1122 = |_EVAL_1433;
  assign _EVAL_1064 = _EVAL_1499 & _EVAL_1568;
  assign _EVAL_221 = _EVAL_1645 & _EVAL_959;
  assign _EVAL_1006 = _EVAL_1821 & _EVAL_2021;
  assign _EVAL_1777 = |_EVAL_909;
  assign _EVAL_58 = _EVAL_1662 & _EVAL_1741;
  assign _EVAL_1258 = _EVAL_330 & _EVAL_959;
  assign monitor_1__EVAL_9 = _EVAL_6;
  assign _EVAL_1330 = ~_EVAL_1109;
  assign _EVAL_459 = _EVAL_394 & _EVAL_1741;
  assign _EVAL_1622 = _EVAL_1258 & _EVAL_442;
  assign _EVAL_166 = _EVAL_997 & _EVAL_442;
  assign _EVAL_1651 = _EVAL_1838 & _EVAL_405;
  assign _EVAL_602 = _EVAL_1499 & _EVAL_220;
  assign _EVAL_1585 = _EVAL_586[0];
  assign _EVAL_1802 = _EVAL_1871 & _EVAL_442;
  assign _EVAL_1645 = _EVAL_1499 & _EVAL_1250;
  assign _EVAL_1319 = _EVAL_495 & _EVAL_1086;
  assign _EVAL_2016 = _EVAL_1502[7];
  assign _EVAL_1517 = |_EVAL_1987;
  assign _EVAL_2026 = _EVAL_1674 & _EVAL_1517;
  assign _EVAL_119 = _EVAL_1938 & _EVAL_442;
  assign _EVAL_627 = _EVAL_1333[260];
  assign _EVAL_214 = _EVAL_1333[262];
  assign monitor__EVAL_3 = _EVAL_42;
  assign monitor_1__EVAL_6 = _EVAL_51;
  assign _EVAL_1170 = _EVAL_917 & _EVAL_442;
  assign _EVAL_312 = ~_EVAL_14;
  assign _EVAL_1854 = _EVAL_1674 & _EVAL_1511;
  assign _EVAL_193 = _EVAL_149 & _EVAL_442;
  assign _EVAL_110 = _EVAL_1746 & _EVAL_1780;
  assign _EVAL_596 = _EVAL_1499 & _EVAL_895;
  assign _EVAL_580 = _EVAL_1871 & _EVAL_1780;
  assign _EVAL_762 = _EVAL_1510 & _EVAL_442;
  assign _EVAL_1145 = _EVAL_164 & _EVAL_1780;
  assign _EVAL_1631 = _EVAL_637 & _EVAL_1121;
  assign _EVAL_1491 = _EVAL_1821 & _EVAL_1341;
  assign monitor__EVAL_8 = _EVAL_17;
  assign _EVAL_878 = _EVAL_970 & _EVAL_959;
  assign _EVAL_1292 = _EVAL_1499 & _EVAL_993;
  assign _EVAL_1221 = _EVAL_864 & _EVAL_1121;
  assign _EVAL_1686 = _EVAL_1510 & _EVAL_1780;
  assign _EVAL_1684 = _EVAL_1499 & _EVAL_1237;
  assign _EVAL_1066 = _EVAL_997 & _EVAL_1121;
  assign _EVAL_175 = _EVAL_314 & _EVAL_1086;
  assign monitor_1__EVAL_2 = _EVAL_6;
  assign _EVAL_318 = _EVAL_1499 & _EVAL_1924;
  assign _EVAL_1856 = |_EVAL_2053;
  assign _EVAL_1655 = ~_EVAL_1112;
  assign _EVAL_1494 = _EVAL_1499 & _EVAL_627;
  assign _EVAL_477 = _EVAL_1510 & _EVAL_1741;
  assign _EVAL_1968 = _EVAL_1674 & _EVAL_1608;
  assign _EVAL_719 = _EVAL_1429 & _EVAL_442;
  assign _EVAL_303 = _EVAL_1899 & _EVAL_1121;
  assign _EVAL_1625 = _EVAL_1499 & _EVAL_682;
  assign _EVAL_1005 = _EVAL_1333[268];
  assign _EVAL_1135 = _EVAL_175 & _EVAL_452;
  assign _EVAL_320 = |_EVAL_1500;
  assign _EVAL_260 = |_EVAL_1152;
  assign _EVAL_1293 = |_EVAL_475;
  assign _EVAL_2013 = _EVAL_1258 & _EVAL_1741;
  assign _EVAL_2024 = |_EVAL_723;
  assign _EVAL_551 = _EVAL_1333[273];
  assign _EVAL_752 = _EVAL_221 & _EVAL_1121;
  assign _EVAL_452 = |_EVAL_1775;
  assign _EVAL_835 = _EVAL_1325 & _EVAL_1585;
  assign monitor__EVAL_11 = _EVAL_33;
  assign _EVAL_645 = _EVAL_1674 & _EVAL_695;
  assign _EVAL_711 = _EVAL_1499 & _EVAL_1570;
  assign _EVAL_1916 = _EVAL_1258 & _EVAL_1121;
  assign monitor__EVAL_4 = _EVAL_14;
  assign _EVAL_1360 = _EVAL_1258 & _EVAL_1780;
  assign _EVAL_294 = _EVAL_164 & _EVAL_1741;
  assign _EVAL_1383 = _EVAL_1502[4];
  assign _EVAL_1879 = _EVAL_149 & _EVAL_1780;
  assign _EVAL_962 = _EVAL_1674 & _EVAL_953;
  assign _EVAL_1354 = _EVAL_221 & _EVAL_442;
  assign _EVAL_731 = _EVAL_1821 & _EVAL_1825;
  assign _EVAL_1820 = _EVAL_1469 & _EVAL_1780;
  assign _EVAL_1947 = |_EVAL_1840;
  assign _EVAL_1172 = _EVAL_1434 & _EVAL_959;
  assign _EVAL_1911 = _EVAL_633 & _EVAL_1121;
  assign monitor__EVAL_6 = _EVAL_31;
  assign _EVAL_88 = _EVAL_468 & _EVAL_1410;
  assign _EVAL_488 = _EVAL_1938 & _EVAL_1780;
  assign monitor__EVAL_13 = _EVAL_43;
  assign _EVAL_207 = _EVAL_1502[13];
  assign _EVAL_1214 = _EVAL_1082 & _EVAL_1780;
  assign _EVAL_679 = _EVAL_864 & _EVAL_1741;
  assign _EVAL_1457 = _EVAL_893 & _EVAL_1780;
  assign _EVAL_1106 = _EVAL_1821 & _EVAL_224;
  assign _EVAL_1424 = _EVAL_1082 & _EVAL_442;
  assign monitor_1__EVAL_5 = _EVAL_19;
  assign _EVAL_1570 = _EVAL_1333[275];
  assign _EVAL_843 = _EVAL_1095 & _EVAL_179;
  assign _EVAL_1397 = _EVAL_1564 & _EVAL_1780;
  assign _EVAL_1662 = _EVAL_2010 & _EVAL_959;
  assign _EVAL_1332 = _EVAL_1499 & _EVAL_1321;
  assign _EVAL_683 = _EVAL_1521 & _EVAL_1121;
  assign _EVAL_512 = _EVAL_919 & _EVAL_959;
  assign _EVAL_798 = _EVAL_1499 & _EVAL_1005;
  assign _EVAL_1308 = _EVAL_878 & _EVAL_1780;
  assign _EVAL_468 = _EVAL_1499 & _EVAL_792;
  assign _EVAL_313 = _EVAL_893 & _EVAL_442;
  assign _EVAL_637 = _EVAL_1695 & _EVAL_959;
  assign _EVAL_1198 = _EVAL_1499 & _EVAL_369;
  assign _EVAL_1510 = _EVAL_82 & _EVAL_959;
  assign _EVAL_461 = _EVAL_1277 & _EVAL_393;
  assign monitor_1__EVAL_14 = _EVAL_32;
  assign _EVAL_955 = _EVAL_1821 & _EVAL_1608;
  assign _EVAL_1039 = _EVAL_1469 & _EVAL_1741;
  assign _EVAL_527 = _EVAL_864 & _EVAL_442;
  assign _EVAL_581 = _EVAL_721 & _EVAL_1780;
  assign _EVAL_1065 = _EVAL_586[17];
  assign _EVAL_1521 = _EVAL_602 & _EVAL_959;
  assign _EVAL_329 = _EVAL_917 & _EVAL_1780;
  assign _EVAL_930 = _EVAL_1963 & _EVAL_442;
  assign _EVAL_612 = _EVAL_1821 & _EVAL_1517;
  assign _EVAL_1870 = _EVAL_1469 & _EVAL_442;
  assign _EVAL_236 = _EVAL_1333[207];
  assign _EVAL_181 = _EVAL_746 & _EVAL_1780;
  assign _EVAL_1041 = _EVAL_1499 & _EVAL_1138;
  assign _EVAL_1871 = _EVAL_1654 & _EVAL_959;
  assign _EVAL_1436 = _EVAL_1076 & _EVAL_959;
  assign _EVAL_1535 = _EVAL_1235 & _EVAL_959;
  assign _EVAL_1194 = _EVAL_586[19];
  assign _EVAL_1259 = _EVAL_1824 & _EVAL_1649;
  assign _EVAL_873 = _EVAL_1821 & _EVAL_509;
  assign _EVAL_1840 = _EVAL_1502[6];
  assign _EVAL_1597 = _EVAL_1674 & _EVAL_1293;
  assign _EVAL_1741 = |_EVAL_949;
  assign _EVAL_314 = _EVAL_1325 & _EVAL_416;
  assign _EVAL_583 = _EVAL_1333[256];
  assign _EVAL_208 = _EVAL_1871 & _EVAL_1121;
  assign monitor_1__EVAL = _EVAL_27;
  assign _EVAL_483 = _EVAL_809 & _EVAL_96;
  assign monitor__EVAL_2 = _EVAL_3;
  assign _EVAL_61 = _EVAL_878 & _EVAL_1741;
  assign _EVAL_750 = _EVAL_1871 & _EVAL_1741;
  assign _EVAL_977 = _EVAL_1821 & _EVAL_944;
  assign _EVAL_370 = _EVAL_734 & _EVAL_959;
  assign _EVAL_1277 = _EVAL_1270 & _EVAL_366;
  assign monitor_1__EVAL_4 = _EVAL_54;
  assign _EVAL_424 = _EVAL_1502[8];
  assign _EVAL_764 = _EVAL_1821 & _EVAL_730;
  assign _EVAL_682 = _EVAL_1333[259];
  assign _EVAL_1960 = _EVAL_1674 & _EVAL_730;
  assign _EVAL_1344 = _EVAL_826 & _EVAL_1377;
  assign _EVAL_157 = _EVAL_1963 & _EVAL_1780;
  assign _EVAL_1103 = _EVAL_616 & _EVAL_117;
  assign _EVAL_401 = _EVAL_1963 & _EVAL_1121;
  assign _EVAL_622 = |_EVAL_183;
  assign _EVAL_1736 = |_EVAL_1398;
  assign _EVAL_1609 = _EVAL_1172 & _EVAL_1741;
  assign _EVAL_1481 = _EVAL_1656 & _EVAL_959;
  assign _EVAL_165 = _EVAL_2045 | _EVAL_14;
  assign _EVAL_1573 = _EVAL_512 & _EVAL_179;
  assign _EVAL_1608 = |_EVAL_1368;
  assign _EVAL_2021 = |_EVAL_256;
  assign _EVAL_1523 = _EVAL_1190 & _EVAL_1741;
  assign _EVAL_1320 = _EVAL_277 & _EVAL_442;
  assign monitor__EVAL_12 = {{2'd0}, _EVAL_1452};
  assign _EVAL_1157 = _EVAL_1499 & _EVAL_381;
  assign _EVAL_780 = _EVAL_1821 & _EVAL_1402;
  assign _EVAL_547 = ~_EVAL_1699;
  assign _EVAL_662 = _EVAL_826 & _EVAL_1777;
  assign _EVAL_889 = _EVAL_1674 & _EVAL_1856;
  assign _EVAL_1747 = _EVAL_1333[206];
  assign _EVAL_913 = _EVAL_149 & _EVAL_1121;
  assign _EVAL_1739 = _EVAL_711 & _EVAL_959;
  assign _EVAL_1788 = _EVAL_88 & _EVAL_1121;
  assign _EVAL_646 = _EVAL_1674 & _EVAL_706;
  assign _EVAL_734 = _EVAL_1499 & _EVAL_951;
  assign _EVAL_1589 = _EVAL_1564 & _EVAL_1121;
  assign monitor_1__EVAL_7 = _EVAL_9;
  assign _EVAL_1825 = |_EVAL_1382;
  assign _EVAL_599 = _EVAL_1502[3:0];
  assign _EVAL_1799 = _EVAL_1429 & _EVAL_1780;
  assign _EVAL_1237 = _EVAL_1333[267];
  assign _EVAL_1551 = _EVAL_1739 & _EVAL_1780;
  assign _EVAL_1143 = _EVAL_1842 & _EVAL_367;
  assign _EVAL_1484 = _EVAL_835 & _EVAL_2018;
  assign _EVAL_251 = _EVAL_1333[269];
  assign _EVAL_1395 = _EVAL_633 & _EVAL_1741;
  assign _EVAL_1797 = _EVAL_1259 & _EVAL_1112;
  assign _EVAL_371 = _EVAL_370 & _EVAL_442;
  assign _EVAL_1893 = _EVAL_1499 & _EVAL_251;
  assign monitor__EVAL_9 = _EVAL_36;
  assign _EVAL_1174 = |_EVAL_424;
  assign _EVAL_102 = _EVAL_1510 & _EVAL_1121;
  assign _EVAL_774 = _EVAL_318 & _EVAL_959;
  assign _EVAL_1550 = _EVAL_1165 & _EVAL_1780;
  assign _EVAL_1487 = _EVAL_774 & _EVAL_1121;
  assign _EVAL_1699 = _EVAL_1981 | _EVAL_14;
  assign _EVAL_630 = |_EVAL_599;
  assign _EVAL_378 = _EVAL_1325 & _EVAL_778;
  assign _EVAL_153 = _EVAL_1502[12];
  assign _EVAL_1205 = _EVAL_633 & _EVAL_1780;
  assign _EVAL_1668 = _EVAL_164 & _EVAL_442;
  assign _EVAL_255 = ~_EVAL_1305;
  assign _EVAL_1100 = _EVAL_746 & _EVAL_1741;
  assign _EVAL_514 = _EVAL_1521 & _EVAL_1780;
  assign _EVAL_197 = |_EVAL_1422;
  assign _EVAL_932 = _EVAL_774 & _EVAL_442;
  assign _EVAL_1456 = _EVAL_1521 & _EVAL_442;
  assign _EVAL_584 = _EVAL_997 & _EVAL_1741;
  assign _EVAL_1413 = _EVAL_1521 & _EVAL_1741;
  assign _EVAL_792 = _EVAL_1333[0];
  assign _EVAL_365 = _EVAL_1319 & _EVAL_367;
  assign _EVAL_1771 = _EVAL_1285 == 3'h0;
  assign _EVAL_1649 = ~_EVAL_1327;
  assign _EVAL_1382 = _EVAL_1502[10];
  assign _EVAL_1746 = _EVAL_95 & _EVAL_959;
  assign _EVAL_1190 = _EVAL_798 & _EVAL_959;
  assign _EVAL_1095 = _EVAL_1829 & _EVAL_959;
  assign _EVAL_1121 = |_EVAL_554;
  assign _EVAL_123 = |_EVAL_279;
  assign _EVAL_1963 = _EVAL_1041 & _EVAL_959;
  assign _EVAL_1926 = _EVAL_1502[21];
  assign monitor__EVAL_0 = _EVAL;
  assign _EVAL_164 = _EVAL_1670 & _EVAL_959;
  assign _EVAL_2038 = _EVAL_1172 & _EVAL_442;
  assign _EVAL_330 = _EVAL_1499 & _EVAL_449;
  assign _EVAL_1433 = _EVAL_1502[18];
  assign _EVAL_804 = _EVAL_1325 & _EVAL_658;
  assign _EVAL_1037 = _EVAL_746 & _EVAL_1121;
  assign _EVAL_947 = _EVAL_1674 & _EVAL_1764;
  assign monitor__EVAL_10 = _EVAL;
  assign monitor_1__EVAL_8 = _EVAL_49;
  assign _EVAL_1493 = _EVAL_1821 & _EVAL_1777;
  assign _EVAL_672 = _EVAL_893 & _EVAL_1121;
  assign _EVAL_808 = _EVAL_1436 & _EVAL_1121;
  assign _EVAL_1393 = _EVAL_394 & _EVAL_1780;
  assign _EVAL_615 = _EVAL_1746 & _EVAL_442;
  assign _EVAL_1981 = _EVAL_1855 | _EVAL_1112;
  assign _EVAL_1766 = _EVAL_1502[28:23];
  assign _EVAL_113 = _EVAL_1270 & _EVAL_1771;
  assign _EVAL_167 = _EVAL_1963 & _EVAL_1741;
  assign _EVAL_1670 = _EVAL_1499 & _EVAL_1575;
  assign _EVAL_816 = _EVAL_1502[15:1];
  assign _EVAL_1462 = _EVAL_1625 & _EVAL_959;
  assign _EVAL_824 = _EVAL_721 & _EVAL_1121;
  assign _EVAL_1098 = _EVAL_1270 & _EVAL_639;
  assign monitor__EVAL_1 = _EVAL_33;
  assign _EVAL_93 = _EVAL_721 & _EVAL_442;
  assign _EVAL_771 = _EVAL_1502[19];
  assign _EVAL_1656 = _EVAL_1499 & _EVAL_551;
  assign _EVAL_872 = |_EVAL_1598;
  assign _EVAL_1750 = _EVAL_1602 & _EVAL_117;
  assign _EVAL_469 = _EVAL_806 & _EVAL_1121;
  assign _EVAL_1531 = _EVAL_637 & _EVAL_1780;
  assign _EVAL_59 = _EVAL_1481 & _EVAL_1780;
  assign monitor_1__EVAL_10 = _EVAL_14;
  assign _EVAL_796 = _EVAL_1674 & _EVAL_944;
  assign _EVAL_1351 = _EVAL_394 & _EVAL_1121;
  assign _EVAL_1401 = _EVAL_1470 & _EVAL_179;
  assign _EVAL_909 = _EVAL_1502[11];
  assign _EVAL_953 = |_EVAL_1926;
  assign _EVAL_179 = |_EVAL_1815;
  assign _EVAL_1930 = _EVAL_826 & _EVAL_260;
  assign _EVAL_693 = _EVAL_1462 & _EVAL_1741;
  assign _EVAL_1883 = _EVAL_1821 & _EVAL_630;
  assign _EVAL_406 = _EVAL_1270 & _EVAL_1841;
  assign monitor__EVAL_14 = _EVAL_30;
  assign _EVAL_1357 = _EVAL_255 & _EVAL_385;
  assign _EVAL_1225 = _EVAL_1821 & _EVAL_948;
  assign _EVAL_160 = _EVAL_806 & _EVAL_1780;
  assign _EVAL_1725 = _EVAL_1481 & _EVAL_442;
  assign _EVAL_183 = _EVAL_1502[3];
  assign _EVAL_442 = |_EVAL_1716;
  assign _EVAL_997 = _EVAL_269 & _EVAL_959;
  assign _EVAL_918 = _EVAL_1739 & _EVAL_442;
  assign _EVAL_1673 = {{1'd0}, _EVAL_385};
  assign _EVAL_1182 = _EVAL_1739 & _EVAL_1121;
  assign _EVAL_681 = _EVAL_826 & _EVAL_1341;
  assign _EVAL_826 = _EVAL_492 & _EVAL_1086;
  assign _EVAL_1299 = _EVAL_826 & _EVAL_2024;
  assign _EVAL_1093 = _EVAL_1899 & _EVAL_1741;
  assign _EVAL_1120 = _EVAL_1499 & _EVAL_136;
  assign _EVAL_806 = _EVAL_1064 & _EVAL_959;
  assign _EVAL_224 = |_EVAL_207;
  assign _EVAL_1499 = _EVAL_904 & _EVAL_1876;
  assign _EVAL_209 = _EVAL_1429 & _EVAL_1741;
  assign _EVAL_1831 = _EVAL_806 & _EVAL_1741;
  assign _EVAL_404 = _EVAL_633 & _EVAL_442;
  assign _EVAL_879 = _EVAL_864 & _EVAL_1780;
  assign _EVAL_492 = _EVAL_1325 & _EVAL_914;
  assign _EVAL_695 = |_EVAL_1990;
  assign _EVAL_579 = _EVAL_149 & _EVAL_1741;
  assign _EVAL_616 = _EVAL_1098 & _EVAL_393;
  assign monitor_1__EVAL_0 = _EVAL_19;
  assign _EVAL_2010 = _EVAL_1499 & _EVAL_1508;
  assign _EVAL_944 = |_EVAL_1383;
  assign _EVAL_533 = ~_EVAL_519;
  assign _EVAL_983 = _EVAL_1938 & _EVAL_1121;
  assign _EVAL_1554 = _EVAL_1190 & _EVAL_1780;
  assign _EVAL_864 = _EVAL_738 & _EVAL_959;
  assign _EVAL_1896 = _EVAL_1469 & _EVAL_1121;
  assign _EVAL_1470 = _EVAL_77 & _EVAL_959;
  assign _EVAL_1152 = _EVAL_1502[7:4];
  assign _EVAL_338 = |_EVAL_1766;
  assign _EVAL_1654 = _EVAL_1499 & _EVAL_1117;
  assign _EVAL_1034 = _EVAL_175 & _EVAL_985;
  assign _EVAL_509 = |_EVAL_771;
  assign _EVAL_1003 = _EVAL_1333[261];
  assign _EVAL_387 = _EVAL_1662 & _EVAL_442;
  assign _EVAL_524 = _EVAL_1333[192];
  assign _EVAL_151 = _EVAL_1325 & _EVAL_1065;
  assign _EVAL_1117 = _EVAL_1333[265];
  assign _EVAL_78 = _EVAL_1325 & _EVAL_1498;
  assign _EVAL_402 = _EVAL_1662 & _EVAL_1780;
  assign _EVAL_1434 = _EVAL_1499 & _EVAL_890;
  assign _EVAL_1266 = _EVAL_1564 & _EVAL_1741;
  assign _EVAL_136 = _EVAL_1333[257];
  assign _EVAL_1952 = _EVAL_990 & _EVAL_393;
  assign _EVAL_1476 = _EVAL_1436 & _EVAL_1780;
  assign _EVAL_1674 = _EVAL_804 & _EVAL_1086;
  assign _EVAL_2012 = _EVAL_1165 & _EVAL_1121;
  assign _EVAL_142 = _EVAL_1821 & _EVAL_1947;
  assign _EVAL_518 = _EVAL_406 & _EVAL_393;
  assign _EVAL_1366 = _EVAL_277 & _EVAL_1780;
  assign _EVAL_1821 = _EVAL_151 & _EVAL_1086;
  assign _EVAL_1734 = _EVAL_1938 & _EVAL_1741;
  assign _EVAL_1990 = _EVAL_1502[2];
  assign _EVAL_919 = _EVAL_1499 & _EVAL_1747;
  assign _EVAL_703 = _EVAL_221 & _EVAL_1741;
  assign _EVAL_1469 = _EVAL_1684 & _EVAL_959;
  assign _EVAL_1661 = _EVAL_893 & _EVAL_1741;
  assign _EVAL_106 = _EVAL_746 & _EVAL_442;
  assign _EVAL_1892 = _EVAL_1535 & _EVAL_442;
  assign _EVAL_720 = _EVAL_88 & _EVAL_442;
  assign _EVAL_656 = _EVAL_1172 & _EVAL_1780;
  assign _EVAL_1228 = _EVAL_774 & _EVAL_1741;
  assign _EVAL_1235 = _EVAL_1499 & _EVAL_788;
  assign _EVAL_706 = |_EVAL_1002;
  assign _EVAL_1564 = _EVAL_1157 & _EVAL_959;
  assign _EVAL_495 = _EVAL_1325 & _EVAL_1194;
  assign _EVAL_1902 = _EVAL_1499 & _EVAL_552;
  assign _EVAL_1647 = _EVAL_917 & _EVAL_1121;
  assign _EVAL_1624 = _EVAL_370 & _EVAL_1121;
  assign _EVAL_324 = _EVAL_1862 & _EVAL_367;
  assign _EVAL_1806 = _EVAL_1462 & _EVAL_1121;
  assign _EVAL_1626 = _EVAL_1333[263];
  assign monitor_1__EVAL_12 = {{2'd0}, _EVAL_1876};
  assign _EVAL_1287 = _EVAL_1662 & _EVAL_1121;
  assign _EVAL_1511 = |_EVAL_1704;
  assign _EVAL_1165 = _EVAL_1120 & _EVAL_959;
  assign _EVAL_1955 = _EVAL_1502[5];
  assign _EVAL_1890 = _EVAL_277 & _EVAL_1741;
  assign _EVAL_250 = _EVAL_1674 & _EVAL_622;
  assign _EVAL_1938 = _EVAL_1291 & _EVAL_959;
  assign _EVAL_409 = _EVAL_774 & _EVAL_1780;
  assign _EVAL_398 = _EVAL_1821 & _EVAL_1680;
  assign _EVAL_1076 = _EVAL_1499 & _EVAL_1795;
  assign _EVAL_588 = _EVAL_1746 & _EVAL_1121;
  assign _EVAL_220 = _EVAL_1333[271];
  assign _EVAL_1810 = _EVAL_1821 & _EVAL_1122;
  assign _EVAL_194 = _EVAL_826 & _EVAL_630;
  assign _EVAL_893 = _EVAL_1528 & _EVAL_959;
  assign _EVAL_1250 = _EVAL_1333[276];
  assign _EVAL_1665 = _EVAL_1190 & _EVAL_1121;
  assign _EVAL_539 = _EVAL_394 & _EVAL_442;
  assign _EVAL_1500 = _EVAL_1502[23:13];
  assign _EVAL_1270 = sb2tlOpt__EVAL_27 | sb2tlOpt__EVAL_12;
  assign _EVAL_573 = _EVAL_721 & _EVAL_1741;
  assign _EVAL_1429 = _EVAL_1332 & _EVAL_959;
  assign _EVAL_1818 = _EVAL_1535 & _EVAL_1121;
  assign _EVAL_1495 = _EVAL_1535 & _EVAL_1780;
  assign _EVAL_1924 = _EVAL_1333[258];
  assign _EVAL_558 = _EVAL_637 & _EVAL_1741;
  assign _EVAL_1598 = _EVAL_1502[11:5];
  assign _EVAL_2053 = _EVAL_1502[1];
  assign _EVAL_232 = _EVAL_1821 & _EVAL_1736;
  assign monitor_1__EVAL_1 = _EVAL_30;
  assign _EVAL_1478 = _EVAL_461 & _EVAL_117;
  assign _EVAL_663 = _EVAL_1502[31:29];
  assign _EVAL_1764 = |_EVAL_663;
  assign _EVAL_95 = _EVAL_1499 & _EVAL_907;
  assign _EVAL_1514 = _EVAL_1333[272];
  assign _EVAL_2029 = _EVAL_1082 & _EVAL_1121;
  assign _EVAL_256 = _EVAL_1502[17];
  assign _EVAL_571 = _EVAL_1821 & _EVAL_123;
  assign _EVAL_394 = _EVAL_1494 & _EVAL_959;
  assign _EVAL_1444 = _EVAL_1462 & _EVAL_442;
  assign _EVAL_1377 = |_EVAL_1492;
  assign _EVAL_1110 = _EVAL_175 & _EVAL_197;
  assign _EVAL_1878 = _EVAL_997 & _EVAL_1780;
  assign _EVAL_405 = _EVAL_1096 == 2'h3;
  assign _EVAL_292 = _EVAL_1082 & _EVAL_1741;
  assign _EVAL_1838 = _EVAL_1259 & _EVAL_1655;
  assign _EVAL_1218 = _EVAL_1674 & _EVAL_872;
  assign _EVAL_1967 = _EVAL_1270 & _EVAL_1162;
  assign _EVAL_619 = _EVAL_1674 & _EVAL_338;
  assign monitor_1__EVAL_13 = _EVAL_51;
  assign _EVAL_659 = _EVAL_370 & _EVAL_1780;
  assign _EVAL_149 = _EVAL_1246 & _EVAL_959;
  assign _EVAL_721 = _EVAL_62 & _EVAL_959;
  assign _EVAL_489 = _EVAL_1502[14];
  assign _EVAL_100 = _EVAL_1499 & _EVAL_583;
  assign _EVAL_2048 = _EVAL_1481 & _EVAL_1741;
  assign _EVAL_1671 = _EVAL_1739 & _EVAL_1741;
  always @(posedge _EVAL_30) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1393 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6718703)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1038 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3cdaf077)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1267 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1c00d9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1066 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da928c29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1348 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94f4163d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a44b7e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1311 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(610bc934)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1858 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b69a7387)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_666 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8aa02d8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_386 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e08a847)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_913 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91948d74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1424 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a21b3344)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1534 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10a90af8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98ab3488)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d88a029b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1985 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e07903ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1395 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63a72763)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1205 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efa37909)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1367 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe3ac26a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1218 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38b49ac8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_888 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d99bf026)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_395 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60c025ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1364 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc1d7295)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1354 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81833a16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1463 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80b764ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1731 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c784228f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b78abb3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_522 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2413677)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1093 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bed97d6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1148 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3acb473e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1006 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26ad863)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_395 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93acfb47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1726 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(542a8168)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_703 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1763f44e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1622 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4122f57f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2047 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98dd9043)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_389 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d05c6d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_371 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3c9a1f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1100 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0283cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1709 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78d739e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a4f9f69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1850 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2f9c0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1110 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e9ee9c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1898 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68b1b500)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2031 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c9ff8f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1539 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(518c4e14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_573 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bda2c2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1985 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(156ceeb9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_879 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec9d5a39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_645 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b614daf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1290 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3829994e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_849 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99e30811)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1683 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d402c630)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(829701ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1658 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a4d752)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_419 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(555fc0ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2041 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e2f84cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1493 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7dba7b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_571 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(700285a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_801 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5aa4135)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_801 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8614e83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_984 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccfc4eb4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_656 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dbb732a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_898 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f6d10d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_454 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a22155e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3dc6664d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_693 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a20b519)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_766 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b4df4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_694 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30952318)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_346 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34d7666)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_913 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea9c0b77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3cda5f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1624 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58ad73a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2031 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b42b681e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1992 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8fb2953)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_697 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d82759a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2013 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ea4b479)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38f8106d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(170cce1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1734 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47bd99f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_691 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1c0671b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_401 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5bbf705)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1613 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62e471)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1958 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(995682be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_577 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa68ce54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1916 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b6e18388)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_883 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77c6958e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_519 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd8e510a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1357 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2dd25af7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1668 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed39b5a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1791 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(666e590c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_731 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d0a2376)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_505 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98976029)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1731 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9048a374)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1308 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed5ffd99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1496 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b84ce8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1266 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(557c39f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_898 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c88ab927)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76c688c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76f06067)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(967b3f10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24178d15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_409 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb5f29d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2048 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7e2286a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_853 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24ab9a5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1381 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9ef7721)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f3cb64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(667f85f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc784a2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1852 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3d1443f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1105 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b344118e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef31d416)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c83d985e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_961 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c554130)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_861 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd4bd484)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_573 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76080f11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1516 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a40ac00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_983 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9ee3a9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9ecfe55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c3e561f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1640 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b34fa682)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1802 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7649ec7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_623 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34e3009f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92733da8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_497 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(747e90f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_337 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd41a9cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(486b9d98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1958 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de10c600)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1026 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c459e697)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1725 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ae3d026)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_472 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40fc13b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_614 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89675037)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1906 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5c5282a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1916 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1424c6fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_648 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12776ca5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1409 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75da79aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1799 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed79347d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1573 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1dfbbea3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1686 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(246b3b9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_387 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2015a57a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1523 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a80cf8b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1892 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c8af73d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1890 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be25c21a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_703 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d91e324)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_719 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d70e22fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1103 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7b29ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fc1576b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1977 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3fdaa80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1247 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e23895ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1957 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b4c82ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_977 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(542cb533)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(126ecb0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_584 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fa053c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_324 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc904dcc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_643 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(439e9e4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1925 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aed984f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1589 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6a8245c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_780 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b89117a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1875 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb6ac500)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1366 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87161d2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_866 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(960c8931)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1456 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2e3eb86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1527 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48ebbbb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_843 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4b367d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_752 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93350176)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_811 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27bc24f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0dbb88d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1487 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3c58aca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1267 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc48f00c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1255 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8b208ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1892 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53297524)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1628 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2dfcca8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1245 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dff9bf07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1609 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31d38b65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_477 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6434f120)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_580 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46da8340)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_859 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f26300d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_759) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_683 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46cd0be6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1792 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ce852bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_681 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3723620)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1413 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef5f3234)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2013 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6b896fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(243e99d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1331 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f63bcffb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ae84668)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_427 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46bbb18e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_337 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb4f57e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1493 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1457376a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1647 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb790c32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_731 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(751ab156)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_685 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9263210)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1609 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b803e5aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1478 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54868ef6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1878 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71da874)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1034 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8ecb4ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1354 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d09d222)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1106 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8dc89d21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1906 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7e3cc9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1070 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8de8d4c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_581 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96dfdeb6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_763 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d20d5f78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1537 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41b54a68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1476 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bff16c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1822 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(191977f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1837 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab9c0218)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1532 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0dea9cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2017 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b6261f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_824 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ae1603a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1350 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(224ca468)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_842 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c83654d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1366 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4511cd1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1531 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4affb1dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_547) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(628ac917)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1317 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5413e8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1145 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58a5b9e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1487 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e6aa3f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1308 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b82771ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1628 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(883e15f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1805 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bece093d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_821 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c56a53ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1879 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bf3ed81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1559 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d994432)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_85 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b43169f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_666 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f8e8896)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4819da16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1411 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f20cb9fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(232bbab9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1495 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee45801)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1227 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf10e34f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_597 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9887a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_398 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee52154c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_929 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92d54966)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2026 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee7d573)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1348 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8821be1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1802 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db1950a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1858 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(886a05e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1837 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea03ddc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1299 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc9de603)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1831 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(934b5f90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_477 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c1df3a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1338 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf6b1273)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1785 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd779f8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1083 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b658931)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1424 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43a195ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1115 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b87f14c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_638 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed856937)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_579 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22e0c1fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1006 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78a6b627)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1879 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(237505b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_752 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11aafb07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1228 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e93b014)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1203 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(111815df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1145 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1aff897a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_873 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81d9f294)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_407 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb3a8b56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1445 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e68f7e92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_800 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e8cfa25)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(226bc204)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2012 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6b24db3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2026 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(966f5562)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1028 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fcd73b26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1988 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50b4dc80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1022 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca15f147)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_977 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a09191be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_324 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33a0debb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6033fb31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_973 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d3ba9d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1396 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6388b1d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(698d4f2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_687 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c0ccc87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_443 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1b7539c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_329 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36e90ede)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1890 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3e104a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2038 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b947394)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_402 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a410be97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_759) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdc770d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1367 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(850968aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_607 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ed382c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_472 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a057bd1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1545 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b17aa9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_837 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e18e7065)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1714 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4999b0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4359cad7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2043 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7156ac8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1532 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(259aa631)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78801ba5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2022 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1039a174)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(795a66b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_523 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a1b4e3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1683 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76e1f651)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1379 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4494f61a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_976 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fff185c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_571 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(963bfad9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1342 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed76c2da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1135 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a494088)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ea1a8a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37960285)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_612 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a76a3ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_705 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2a04a62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_439 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7e97b2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_371 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dffaa8d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_612 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0fbc547)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1785 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b049f35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1552 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99d04840)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1960 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c40e33cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_469 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f672620)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ecf1d3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1538 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80fd86b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1299 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(306c02ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_346 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fac83098)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1630 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fd25b87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_629 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91804ff1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_685 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b4c7946)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_340 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45fe93d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1326 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe5986c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_825 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f5daad6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1039 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d080c6d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_983 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(765ebbe9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1137 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65291109)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1375 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a03745e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_837 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3367031)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1393 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e79eeac0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_523 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d59b34e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2037 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b9aebb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_619 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(191977f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1203 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97000436)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1182 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e58278eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1135 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43b436cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_808 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95a201a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_580 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc9e2da0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1554 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5174025b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_629 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9707d84b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1448 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c100318)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_588 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(604e6d6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1717a16e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74c5844c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1946 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42a03b4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_549 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b37d8e0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1573 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f97aad06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1100 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2febabf9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b989078d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9d473ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_558 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7db5c2d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1170 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb87ed6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1822 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8ecb4ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1264 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(286259f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2039 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f72cebfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1880 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1626993)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6204f836)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1476 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53abcec7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_549 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc3309cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1624 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dda67dab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_873 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5dd181a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(924ddf77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1381 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdbd4455)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_561 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32dae759)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df3cbfb1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_460 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(903ce25a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1444 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2e0e0b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1850 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff8786b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1727 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a626cf9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1023 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae9e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_440 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b8302d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45aaafe1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1137 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(855c7d0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1531 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e3695ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(277006a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_705 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(605ff5c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_976 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27ec087a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_766 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e774e4ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_248 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62240664)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_831 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(298a42bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_619 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8ecb4ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1996 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a80a866)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1287 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48c342fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_519 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c92ce416)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2033 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4678be71)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8274b7fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1946 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99736d7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9ea351a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1648 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9772b63e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1750 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18355ec3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1266 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59d6b4e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1159 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61d77e07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1661 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81eea502)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1485 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27ddaef0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_681 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e30c9632)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1792 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b2cd183)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1343 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40ff444d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1968 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e4202cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1463 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38db6dfd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1977 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd4d8259)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1485 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1df42e62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_556 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f715309)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fba86cf5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1225 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b5de798)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1344 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c88cfd6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_460 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f57c478a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1129 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d5d3239)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_824 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7edbecd5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_784 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67cf2aa1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fa86e6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1615 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52c49248)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1883 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74e180ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16799fed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_719 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31fd8f15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_808 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7318303d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_687 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6625f8a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1491 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91082b3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_747 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1761e43c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2052 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df6dd3bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1852 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24d0c934)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2029 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e6fa4c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1342 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7889462c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1375 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dea35549)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1457 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb34e47a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_672 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3cc3ab1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1589 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cf2868)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8ecb4ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_763 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73d0d7d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1869 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33bbe629)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_930 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81d624e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2028 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f37d2d52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_825 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d61f7a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_426 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1c712e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1794 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdab4ee8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae5c02e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_683 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6504a70e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1552 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aecef768)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(585643c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_539 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a545cce5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_232 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(191977f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db444bb1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1491 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43ec2944)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_404 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22ffc49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1105 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6e194fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_764 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db7dae42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1028 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca5d454c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2037 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(830f9e69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1350 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3158b9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1665 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9cbdf9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1344 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6acbc23d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70d6a54a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1925 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f9ad5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1148 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a8d28c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de528f26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1289 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d93b164e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1271 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5010d98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1160 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e82322d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_645 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64034a6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1409 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d35f875c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1516 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1513086)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_764 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(913a57cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_462 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc88df77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1043 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(460f8b03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_597 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(408db4da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_861 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c283efd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1431 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16d7699e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_918 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a3b6c1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_780 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8d58f38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1880 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(887214aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1707 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4dc79f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1170 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4c7cbea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39e380ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_961 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46f181b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1671 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8909c0da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_693 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c2f9fee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1360 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf2f5099)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1870 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bba1a05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1255 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91abc0e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_955 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf31e13f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_511 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4a6dc95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_567 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac19f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1099 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29e64578)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1214 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2373d465)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1523 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(389ab718)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_963 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ead326ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1820 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ddcca87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1869 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff952f41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2003 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4203e63f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1527 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad4bfd4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1676 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a3d28c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1326 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86d509fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_750 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5fbd9c73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be7cee42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_866 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69156e3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_511 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ccaaa54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1059 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5c4fc03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1280 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1d4eecb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2048 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(181781e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1475 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(347562a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1401 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54cab99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1445 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35df1fa9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_615 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39628e9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_459 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b81ef0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1788 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f7ceec4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1143 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b599d8e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_539 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11e549d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2028 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(941090e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_962 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0591b9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1631 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b8d3646)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2043 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb102807)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1646 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a905155)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1630 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bfdad4e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1278 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e3048f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_725 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6c97496)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1185 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e98f6b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1505 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df66f6d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1640 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(402e7853)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1359 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21c6f538)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1621 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(271ba828)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1665 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d984994)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64f2376b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_679 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50fb62c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_648 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a627493)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1047 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e677e667)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1338 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b99277af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2017 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a995e1d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1709 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70aa406f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1757 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab7725c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_329 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c12d587c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_726 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c7aad85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b3f31b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_842 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6507261b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46791c43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_707 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6362533)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12fa9eb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1763 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc8d05d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1236 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7eb6c11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1214 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ad8d4d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_694 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58c8e36a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_462 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54b8d7bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1512 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a7fc4b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1247 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a02b4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1909 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3613aad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_747 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3dd28b0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_527 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e963496)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1221 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61080962)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1806 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71f18d9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1225 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99d830b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_871 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d618e33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1896 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21233c80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1185 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75925830)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_796 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7eb9efa2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_387 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c9c9fb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1411 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3f5e669)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_672 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(319abeb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_491 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(527e1dba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1596 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(105338b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1930 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8ecb4ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_488 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bb69273)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1143 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef48d72a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0e47e0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1831 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58f94b09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb197e50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1129 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f49ab032)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1245 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd3aef79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1859 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e1a6ff9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1159 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62d028ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_879 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db36a141)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_592 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(803f9c71)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_662 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(191977f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_883 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1df98018)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_659 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3433772)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_707 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba3905dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1022 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(686ced20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_843 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6300c37a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1622 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(284cbe9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3be3bff4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1115 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f53f6079)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1834 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41505092)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1648 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56348146)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2047 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(459b877)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_643 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7efc25e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1957 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9431e928)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_646 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e36c573)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1744 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be47845d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1038 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6406ffcb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1744 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fa4ed43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1395 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b4c31f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1039 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8da2e85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1280 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cf06edf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1791 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d661fc89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1351 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1198bfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1495 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35bad4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_547) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_389 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbc11529)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1854 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b707b32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_656 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1074052)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1911 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e50ba90a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1554 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(934ee9f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1809 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d1fadbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_720 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2fd4e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_527 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41629e77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_438 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa0cd9b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_859 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9faf14e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1278 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(905875e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1834 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45b37841)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1160 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95b50ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1550 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6716906)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e91aee24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1810 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a9202a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2d14083)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1854 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(169fa2b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_770 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa9a53a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_459 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0e97cf2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1550 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20aa2bfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8f0a27e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8c29fc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1583 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(543d1353)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_635 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2669447b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65229a6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1351 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4816603)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1448 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99508172)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1061 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ffb34f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_614 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd972ba0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1988 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4ac928)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2038 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b34b1dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1534 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b20229)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1583 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8a9ca15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1207 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(861390b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_483 & _EVAL_759) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1878 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b87316a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1551 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65cbcdd8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_613 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee43b8af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1317 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b8ba5cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1359 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f56a0ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_479 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e8e15d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_929 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f7718cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_505 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(849644e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1930 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(191977f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1757 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62d0e47e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1397 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cebe2ab9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_615 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e25c3fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1290 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6bb5419c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_401 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0112e6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1431 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16a2d578)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_96 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4373f7a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_762 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d247a66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_762 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ded99cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1799 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(777c3558)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_426 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3de23f5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1788 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1efd4ffd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bfdc4a2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1457 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c220e8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1875 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(398c901)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1539 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a81bf03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2035 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63b7f9b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1037 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(152bb908)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1207 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df30b250)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_558 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4193f316)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2b1d739)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_938 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc384926)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1413 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ce10ab1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_888 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b3985f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1730 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bb8a6fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d11e50b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1794 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94eceb96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1696 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4005f2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_588 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ab26fb6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1661 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4cf802ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1734 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fba44ae2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_947 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70fadc7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef9eb483)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2012 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9204f5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1227 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ca78b36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1496 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(970daf8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1551 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36bedc85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9029997)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_514 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(141008a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1343 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c6512d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1597 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf709638)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_479 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6519cca2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1070 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46e37578)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1904 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b01c443)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d82a1556)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_848 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(640f1d87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(339d50e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2003 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c4c09b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1034 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(191977f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1023 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fba9ea8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_592 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c14d692e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1725 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0be4b70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_849 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46031fed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1401 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35383319)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2029 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9333c729)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1818 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca2b60a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_930 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1281e545)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1205 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2fc354e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_962 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b73c67d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1444 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c5a188e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_823 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6bf666a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_947 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96071b91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_965 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3be986ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1545 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(695d2faa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1898 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45b55f4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_963 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b651c99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_438 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3699950f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_340 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43e3c9a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1538 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f63e5043)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e89bffd3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_581 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(869e1dc4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56b239a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(feaeb366)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9565a639)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1615 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4330efd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e772ef1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1026 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53acbb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1909 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23fd188)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_386 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c0bcc1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1271 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e91e445)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6329ea47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1809 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5657555)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1264 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a13bbb2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_800 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3598c2ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_607 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94c600e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1099 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ee60045)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1597 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72bd9649)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_556 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b1d3339)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2052 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1efaead)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_469 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7291a160)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_726 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b2570c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1047 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfe738ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1651 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6031993f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_514 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81234877)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_439 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e340042)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_823 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(564be713)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(673e88cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1651 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_398 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(103feb10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88276a1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1061 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0c9c43a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6a27a6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_497 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2d0079c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1658 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad1d77fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1331 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e49ae14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b627b39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1059 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56a42998)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_955 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b346f7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_491 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffb66f77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_635 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1a225ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_414 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(639c5692)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_811 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d26ff4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1805 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6598cd5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1960 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a25a5ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1218 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a975f6d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1613 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4aa6f3db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_483 & _EVAL_759) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(268676bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1060 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b97769b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1676 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76367449)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0e3fb9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_440 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af25d956)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1883 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30fa0293)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87311ce0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_691 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a146d8d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_662 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8ecb4ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1818 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b52573d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efd365a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4ed3bd6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_848 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(862b45ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1221 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c80797be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_984 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d8a303)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1379 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(addc8cd5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_572 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f255c2f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_414 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bda92a47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1475 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3011c77e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_407 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c77ade3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1763 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9963408a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1066 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b1fcf2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_932 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2aacb19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_831 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(574ee0ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77844be4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_889 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1badfda6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_623 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(922f8d34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1320 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d51bee91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2039 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b442c1b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_720 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a200caad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_402 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f25cd5e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1505 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b66c1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_725 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b855b9ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1320 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41dbb2c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1559 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2199a50a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_750 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(195c81de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_409 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68e6e66d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1182 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(634a2dac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1714 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(898cac2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_821 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af73f2fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_572 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8925492)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_419 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5909b74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1647 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba0a70d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_567 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e230e76)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1287 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(185828b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_796 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12847fbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1859 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13f5ca9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1968 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1612a914)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_889 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7eefbbed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1364 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7555a6e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1396 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(569d0806)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_522 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a210434e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_679 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a8e2b28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_938 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aff1b147)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1060 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8657010)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2041 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(561d782d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1730 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3cf7513e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1430 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73e12890)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1093 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4eb8d16c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1236 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfbc2444)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_368 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9dfaa237)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1289 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9887aacb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_646 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46960080)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1537 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(178230c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1512 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4c1f915)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1106 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad52ef29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_638 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(545b76b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2022 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df9d8223)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_784 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f26d461)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_932 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2119c90f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_454 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b3e4c07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1456 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1c91aed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_577 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29548af3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2035 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3ab8232)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1967 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(773cd99d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1668 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(277f99dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afed7ec2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(538ecd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_561 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f29b5c53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_579 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a76a4495)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1397 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cf177d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1043 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21fcf349)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_427 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3cc14a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1110 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40f9fe13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1430 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0beaee5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1896 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85313fd3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3d42133)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1992 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11c765e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf25ac4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1810 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e9aae93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_488 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91770a31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a944b7a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_918 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abe89db9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_871 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b31ba5e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2033 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5eb7fb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(208694ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1707 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b366ab03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1996 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(739ce5ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1646 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b49e3a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1360 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5654a847)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c76b503)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1621 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49bae7a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1311 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59163cdd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1696 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87bae75d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1631 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac34e087)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_613 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68c6aaee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1806 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a80fa655)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1726 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b622a6fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1037 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e6d7407)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1911 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4ede0cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1870 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d75663ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1820 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bb0d84c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1671 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23a0b71)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1686 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5ca0b56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_853 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4839d66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1083 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bdfcd16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_697 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(872c9337)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1596 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c07897e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1228 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f48d7ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_973 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b0ab574)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_965 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f13778d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_659 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e90b60da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
