//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_99(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input  [1:0]  _EVAL_17,
  input         _EVAL_18,
  output        _EVAL_19,
  input         _EVAL_20,
  input         _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  input         _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  input         _EVAL_30,
  input         _EVAL_31,
  output [2:0]  _EVAL_32,
  input         _EVAL_33,
  input         _EVAL_34,
  input         _EVAL_35,
  input         _EVAL_36,
  input         _EVAL_37,
  input         _EVAL_38,
  input         _EVAL_39,
  input         _EVAL_40,
  input         _EVAL_41,
  input         _EVAL_42,
  input         _EVAL_43,
  input         _EVAL_44,
  input         _EVAL_45,
  input         _EVAL_46,
  output        _EVAL_47,
  input         _EVAL_48,
  input         _EVAL_49,
  input         _EVAL_50,
  input         _EVAL_51,
  input         _EVAL_52,
  input         _EVAL_53,
  input         _EVAL_54,
  input         _EVAL_55,
  input         _EVAL_56,
  input         _EVAL_57,
  input         _EVAL_58,
  input         _EVAL_59,
  output        _EVAL_60,
  input         _EVAL_61,
  input         _EVAL_62,
  input         _EVAL_63,
  input         _EVAL_64,
  input         _EVAL_65,
  input         _EVAL_66,
  input         _EVAL_67,
  input         _EVAL_68,
  input         _EVAL_69,
  input  [2:0]  _EVAL_70,
  input         _EVAL_71,
  input         _EVAL_72,
  input  [9:0]  _EVAL_73,
  input         _EVAL_74,
  input         _EVAL_75,
  input         _EVAL_76,
  input         _EVAL_77,
  input         _EVAL_78,
  input         _EVAL_79,
  input         _EVAL_80,
  input         _EVAL_81,
  input         _EVAL_82,
  input         _EVAL_83,
  input  [3:0]  _EVAL_84,
  input         _EVAL_85,
  input         _EVAL_86,
  input         _EVAL_87,
  input         _EVAL_88,
  input         _EVAL_89,
  input         _EVAL_90,
  input         _EVAL_91,
  input         _EVAL_92,
  input         _EVAL_93,
  input         _EVAL_94,
  input         _EVAL_95,
  input         _EVAL_96,
  output [31:0] _EVAL_97,
  input         _EVAL_98,
  input         _EVAL_99,
  input         _EVAL_100,
  input  [31:0] _EVAL_101,
  input         _EVAL_102,
  input         _EVAL_103,
  input         _EVAL_104,
  input         _EVAL_105,
  input         _EVAL_106,
  input         _EVAL_107,
  input         _EVAL_108,
  input         _EVAL_109,
  input         _EVAL_110,
  input         _EVAL_111,
  input         _EVAL_112,
  input         _EVAL_113,
  input         _EVAL_114,
  input         _EVAL_115,
  input         _EVAL_116,
  input         _EVAL_117,
  input         _EVAL_118,
  input         _EVAL_119,
  input         _EVAL_120,
  input         _EVAL_121,
  input         _EVAL_122,
  input         _EVAL_123,
  output [9:0]  _EVAL_124,
  input         _EVAL_125,
  output [1:0]  _EVAL_126,
  input         _EVAL_127,
  input         _EVAL_128,
  input         _EVAL_129,
  input  [27:0] _EVAL_130,
  input         _EVAL_131,
  input         _EVAL_132,
  input         _EVAL_133,
  input         _EVAL_134,
  input         _EVAL_135,
  input         _EVAL_136,
  input         _EVAL_137,
  input         _EVAL_138,
  input         _EVAL_139,
  input         _EVAL_140,
  input         _EVAL_141,
  input         _EVAL_142,
  input         _EVAL_143,
  input         _EVAL_144
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_148;
  wire [31:0] _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_156;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  reg [2:0] _EVAL_167;
  reg  _EVAL_168;
  wire [31:0] _EVAL_170;
  wire  _EVAL_171;
  reg [2:0] _EVAL_172;
  wire  gateways_gateway_45__EVAL;
  wire  gateways_gateway_45__EVAL_0;
  wire  gateways_gateway_45__EVAL_1;
  wire  gateways_gateway_45__EVAL_2;
  wire  gateways_gateway_45__EVAL_3;
  wire  gateways_gateway_45__EVAL_4;
  wire [31:0] _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_184;
  wire  _EVAL_185;
  reg [2:0] _EVAL_189;
  wire [31:0] _EVAL_190;
  reg  _EVAL_193;
  wire  _EVAL_195;
  wire  _EVAL_196;
  reg  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_219;
  reg [2:0] _EVAL_222;
  wire  _EVAL_223;
  wire [9:0] _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_228;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_236;
  wire  _EVAL_238;
  reg [2:0] _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_247;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_265;
  wire [7:0] _EVAL_267;
  wire  _EVAL_270;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  reg  _EVAL_276;
  wire  _EVAL_278;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  reg  _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_288;
  reg [2:0] _EVAL_289;
  wire [31:0] _EVAL_293;
  wire  _EVAL_294;
  wire  _EVAL_295;
  wire  _EVAL_296;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  reg  _EVAL_302;
  wire [126:0] _EVAL_304;
  wire [31:0] _EVAL_309;
  wire [31:0] _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_318;
  wire  _EVAL_320;
  wire [31:0] _EVAL_321;
  wire  _EVAL_322;
  wire  _EVAL_323;
  wire  _EVAL_324;
  reg  _EVAL_325;
  wire  _EVAL_330;
  wire  _EVAL_331;
  wire  _EVAL_333;
  wire  _EVAL_334;
  wire  _EVAL_335;
  wire  _EVAL_337;
  wire  _EVAL_338;
  wire [31:0] _EVAL_339;
  wire  _EVAL_340;
  wire  _EVAL_341;
  wire  _EVAL_342;
  wire  _EVAL_343;
  wire  _EVAL_344;
  reg  _EVAL_350;
  wire  _EVAL_353;
  wire  _EVAL_354;
  reg [2:0] _EVAL_355;
  wire  _EVAL_356;
  wire  _EVAL_362;
  wire  _EVAL_364;
  wire  _EVAL_365;
  wire [31:0] _EVAL_366;
  wire  _EVAL_367;
  wire  _EVAL_368;
  wire  _EVAL_369;
  wire  _EVAL_371;
  wire  gateways_gateway_87__EVAL;
  wire  gateways_gateway_87__EVAL_0;
  wire  gateways_gateway_87__EVAL_1;
  wire  gateways_gateway_87__EVAL_2;
  wire  gateways_gateway_87__EVAL_3;
  wire  gateways_gateway_87__EVAL_4;
  wire  _EVAL_374;
  wire  _EVAL_378;
  wire  _EVAL_379;
  wire  _EVAL_381;
  wire  _EVAL_382;
  wire  _EVAL_383;
  wire  _EVAL_385;
  wire [18:0] _EVAL_386;
  wire  gateways_gateway_58__EVAL;
  wire  gateways_gateway_58__EVAL_0;
  wire  gateways_gateway_58__EVAL_1;
  wire  gateways_gateway_58__EVAL_2;
  wire  gateways_gateway_58__EVAL_3;
  wire  gateways_gateway_58__EVAL_4;
  wire  _EVAL_390;
  reg [7:0] _EVAL_394;
  wire  _EVAL_402;
  wire  _EVAL_403;
  wire  _EVAL_404;
  wire  _EVAL_408;
  wire  _EVAL_410;
  wire  _EVAL_411;
  wire  _EVAL_412;
  reg  _EVAL_414;
  reg  _EVAL_415;
  wire  _EVAL_416;
  wire  _EVAL_421;
  wire  _EVAL_422;
  reg  _EVAL_423;
  wire  _EVAL_425;
  wire [7:0] _EVAL_428;
  wire [31:0] _EVAL_434;
  wire  _EVAL_435;
  wire [31:0] _EVAL_440;
  wire  gateways_gateway_7__EVAL;
  wire  gateways_gateway_7__EVAL_0;
  wire  gateways_gateway_7__EVAL_1;
  wire  gateways_gateway_7__EVAL_2;
  wire  gateways_gateway_7__EVAL_3;
  wire  gateways_gateway_7__EVAL_4;
  reg [7:0] _EVAL_445;
  wire  _EVAL_446;
  wire [31:0] _EVAL_449;
  wire  gateways_gateway_22__EVAL;
  wire  gateways_gateway_22__EVAL_0;
  wire  gateways_gateway_22__EVAL_1;
  wire  gateways_gateway_22__EVAL_2;
  wire  gateways_gateway_22__EVAL_3;
  wire  gateways_gateway_22__EVAL_4;
  wire  gateways_gateway_41__EVAL;
  wire  gateways_gateway_41__EVAL_0;
  wire  gateways_gateway_41__EVAL_1;
  wire  gateways_gateway_41__EVAL_2;
  wire  gateways_gateway_41__EVAL_3;
  wire  gateways_gateway_41__EVAL_4;
  wire  _EVAL_451;
  reg [2:0] _EVAL_456;
  wire  gateways_gateway_111__EVAL;
  wire  gateways_gateway_111__EVAL_0;
  wire  gateways_gateway_111__EVAL_1;
  wire  gateways_gateway_111__EVAL_2;
  wire  gateways_gateway_111__EVAL_3;
  wire  gateways_gateway_111__EVAL_4;
  wire  _EVAL_458;
  reg [2:0] _EVAL_461;
  wire  _EVAL_462;
  wire  _EVAL_463;
  wire  _EVAL_466;
  wire  _EVAL_467;
  wire  _EVAL_468;
  wire [7:0] _EVAL_469;
  wire  _EVAL_471;
  wire  _EVAL_473;
  wire  _EVAL_476;
  wire [31:0] _EVAL_478;
  wire  _EVAL_480;
  wire  gateways_gateway_122__EVAL;
  wire  gateways_gateway_122__EVAL_0;
  wire  gateways_gateway_122__EVAL_1;
  wire  gateways_gateway_122__EVAL_2;
  wire  gateways_gateway_122__EVAL_3;
  wire  gateways_gateway_122__EVAL_4;
  wire  _EVAL_482;
  wire  _EVAL_485;
  wire  _EVAL_487;
  wire  _EVAL_488;
  wire  _EVAL_489;
  wire  _EVAL_490;
  wire [31:0] _EVAL_492;
  wire  _EVAL_495;
  wire  _EVAL_496;
  reg  _EVAL_498;
  wire  _EVAL_499;
  wire [31:0] _EVAL_500;
  wire  _EVAL_504;
  wire  _EVAL_505;
  wire  _EVAL_506;
  wire  _EVAL_509;
  wire  _EVAL_510;
  reg [2:0] _EVAL_513;
  wire  _EVAL_515;
  reg [2:0] _EVAL_517;
  wire  _EVAL_520;
  wire [31:0] _EVAL_524;
  reg  _EVAL_526;
  wire  gateways_gateway_24__EVAL;
  wire  gateways_gateway_24__EVAL_0;
  wire  gateways_gateway_24__EVAL_1;
  wire  gateways_gateway_24__EVAL_2;
  wire  gateways_gateway_24__EVAL_3;
  wire  gateways_gateway_24__EVAL_4;
  wire  gateways_gateway_40__EVAL;
  wire  gateways_gateway_40__EVAL_0;
  wire  gateways_gateway_40__EVAL_1;
  wire  gateways_gateway_40__EVAL_2;
  wire  gateways_gateway_40__EVAL_3;
  wire  gateways_gateway_40__EVAL_4;
  wire  _EVAL_531;
  wire [31:0] _EVAL_532;
  wire  _EVAL_533;
  wire  _EVAL_534;
  wire  _EVAL_536;
  wire  gateways_gateway_102__EVAL;
  wire  gateways_gateway_102__EVAL_0;
  wire  gateways_gateway_102__EVAL_1;
  wire  gateways_gateway_102__EVAL_2;
  wire  gateways_gateway_102__EVAL_3;
  wire  gateways_gateway_102__EVAL_4;
  wire  _EVAL_540;
  wire  gateways_gateway_113__EVAL;
  wire  gateways_gateway_113__EVAL_0;
  wire  gateways_gateway_113__EVAL_1;
  wire  gateways_gateway_113__EVAL_2;
  wire  gateways_gateway_113__EVAL_3;
  wire  gateways_gateway_113__EVAL_4;
  wire  _EVAL_544;
  wire [31:0] _EVAL_547;
  reg  _EVAL_552;
  wire  _EVAL_560;
  wire  gateways_gateway_89__EVAL;
  wire  gateways_gateway_89__EVAL_0;
  wire  gateways_gateway_89__EVAL_1;
  wire  gateways_gateway_89__EVAL_2;
  wire  gateways_gateway_89__EVAL_3;
  wire  gateways_gateway_89__EVAL_4;
  wire  _EVAL_567;
  wire [31:0] _EVAL_569;
  reg [2:0] _EVAL_570;
  wire  _EVAL_571;
  wire  _EVAL_573;
  wire  _EVAL_575;
  wire [9:0] _EVAL_576;
  wire  _EVAL_583;
  wire  _EVAL_584;
  wire  _EVAL_585;
  wire  _EVAL_588;
  wire  _EVAL_590;
  wire  _EVAL_592;
  wire  _EVAL_593;
  reg  _EVAL_594;
  wire  _EVAL_595;
  wire  _EVAL_602;
  wire  _EVAL_603;
  wire  _EVAL_604;
  wire  _EVAL_605;
  wire  _EVAL_607;
  wire  _EVAL_609;
  wire  _EVAL_610;
  reg  _EVAL_612;
  wire  _EVAL_613;
  wire  _EVAL_614;
  wire  _EVAL_615;
  wire  _EVAL_625;
  wire  _EVAL_627;
  wire  gateways_gateway_91__EVAL;
  wire  gateways_gateway_91__EVAL_0;
  wire  gateways_gateway_91__EVAL_1;
  wire  gateways_gateway_91__EVAL_2;
  wire  gateways_gateway_91__EVAL_3;
  wire  gateways_gateway_91__EVAL_4;
  reg [2:0] _EVAL_628;
  wire  _EVAL_630;
  wire  _EVAL_631;
  wire  _EVAL_632;
  wire  gateways_gateway_96__EVAL;
  wire  gateways_gateway_96__EVAL_0;
  wire  gateways_gateway_96__EVAL_1;
  wire  gateways_gateway_96__EVAL_2;
  wire  gateways_gateway_96__EVAL_3;
  wire  gateways_gateway_96__EVAL_4;
  wire  _EVAL_638;
  wire  _EVAL_639;
  wire  _EVAL_640;
  wire  _EVAL_641;
  reg [2:0] _EVAL_642;
  wire  _EVAL_643;
  wire  _EVAL_644;
  wire  gateways_gateway_46__EVAL;
  wire  gateways_gateway_46__EVAL_0;
  wire  gateways_gateway_46__EVAL_1;
  wire  gateways_gateway_46__EVAL_2;
  wire  gateways_gateway_46__EVAL_3;
  wire  gateways_gateway_46__EVAL_4;
  wire  _EVAL_645;
  wire  _EVAL_646;
  wire  gateways_gateway_1__EVAL;
  wire  gateways_gateway_1__EVAL_0;
  wire  gateways_gateway_1__EVAL_1;
  wire  gateways_gateway_1__EVAL_2;
  wire  gateways_gateway_1__EVAL_3;
  wire  gateways_gateway_1__EVAL_4;
  wire  _EVAL_647;
  wire  _EVAL_648;
  wire [1023:0] _EVAL_651;
  wire  _EVAL_652;
  wire  _EVAL_653;
  wire  _EVAL_655;
  wire  gateways_gateway_28__EVAL;
  wire  gateways_gateway_28__EVAL_0;
  wire  gateways_gateway_28__EVAL_1;
  wire  gateways_gateway_28__EVAL_2;
  wire  gateways_gateway_28__EVAL_3;
  wire  gateways_gateway_28__EVAL_4;
  wire  _EVAL_657;
  wire  _EVAL_667;
  reg  _EVAL_668;
  wire [31:0] _EVAL_669;
  wire  _EVAL_670;
  wire  _EVAL_673;
  reg  _EVAL_677;
  wire  _EVAL_678;
  wire  _EVAL_679;
  wire [31:0] _EVAL_683;
  wire  _EVAL_685;
  wire  _EVAL_687;
  wire  _EVAL_688;
  wire [31:0] _EVAL_689;
  wire  _EVAL_691;
  reg [2:0] _EVAL_692;
  wire  _EVAL_693;
  wire  _EVAL_695;
  wire  gateways_gateway_44__EVAL;
  wire  gateways_gateway_44__EVAL_0;
  wire  gateways_gateway_44__EVAL_1;
  wire  gateways_gateway_44__EVAL_2;
  wire  gateways_gateway_44__EVAL_3;
  wire  gateways_gateway_44__EVAL_4;
  wire  _EVAL_696;
  wire  _EVAL_697;
  wire  _EVAL_699;
  reg [2:0] _EVAL_700;
  wire  gateways_gateway_103__EVAL;
  wire  gateways_gateway_103__EVAL_0;
  wire  gateways_gateway_103__EVAL_1;
  wire  gateways_gateway_103__EVAL_2;
  wire  gateways_gateway_103__EVAL_3;
  wire  gateways_gateway_103__EVAL_4;
  wire  gateways_gateway_2__EVAL;
  wire  gateways_gateway_2__EVAL_0;
  wire  gateways_gateway_2__EVAL_1;
  wire  gateways_gateway_2__EVAL_2;
  wire  gateways_gateway_2__EVAL_3;
  wire  gateways_gateway_2__EVAL_4;
  wire  _EVAL_703;
  reg [2:0] _EVAL_707;
  wire  _EVAL_709;
  wire  _EVAL_710;
  wire  _EVAL_712;
  wire  _EVAL_715;
  wire  _EVAL_719;
  wire  _EVAL_721;
  wire  _EVAL_723;
  wire  _EVAL_726;
  reg  _EVAL_727;
  wire  _EVAL_733;
  wire  _EVAL_735;
  wire  _EVAL_736;
  wire  _EVAL_739;
  wire  _EVAL_741;
  wire  gateways_gateway_42__EVAL;
  wire  gateways_gateway_42__EVAL_0;
  wire  gateways_gateway_42__EVAL_1;
  wire  gateways_gateway_42__EVAL_2;
  wire  gateways_gateway_42__EVAL_3;
  wire  gateways_gateway_42__EVAL_4;
  wire [31:0] _EVAL_743;
  reg  _EVAL_744;
  wire  _EVAL_751;
  wire  _EVAL_752;
  wire  _EVAL_753;
  wire  _EVAL_755;
  wire  _EVAL_758;
  wire  _EVAL_759;
  wire  _EVAL_762;
  wire  _EVAL_765;
  reg  _EVAL_770;
  wire  _EVAL_771;
  wire  _EVAL_772;
  wire  _EVAL_775;
  wire  _EVAL_776;
  wire  _EVAL_777;
  reg [2:0] _EVAL_778;
  reg [2:0] _EVAL_779;
  reg  _EVAL_780;
  wire  gateways_gateway_68__EVAL;
  wire  gateways_gateway_68__EVAL_0;
  wire  gateways_gateway_68__EVAL_1;
  wire  gateways_gateway_68__EVAL_2;
  wire  gateways_gateway_68__EVAL_3;
  wire  gateways_gateway_68__EVAL_4;
  wire  _EVAL_783;
  wire  _EVAL_784;
  wire  _EVAL_787;
  wire  gateways_gateway_116__EVAL;
  wire  gateways_gateway_116__EVAL_0;
  wire  gateways_gateway_116__EVAL_1;
  wire  gateways_gateway_116__EVAL_2;
  wire  gateways_gateway_116__EVAL_3;
  wire  gateways_gateway_116__EVAL_4;
  wire  gateways_gateway_84__EVAL;
  wire  gateways_gateway_84__EVAL_0;
  wire  gateways_gateway_84__EVAL_1;
  wire  gateways_gateway_84__EVAL_2;
  wire  gateways_gateway_84__EVAL_3;
  wire  gateways_gateway_84__EVAL_4;
  wire  _EVAL_792;
  wire  _EVAL_793;
  wire  _EVAL_794;
  wire  _EVAL_796;
  reg [2:0] _EVAL_797;
  wire  _EVAL_799;
  wire  _EVAL_801;
  wire  _EVAL_804;
  reg [2:0] _EVAL_809;
  wire [2:0] _EVAL_810;
  reg  _EVAL_811;
  reg  _EVAL_813;
  wire [31:0] _EVAL_815;
  wire  _EVAL_817;
  reg  _EVAL_819;
  wire  _EVAL_820;
  wire  gateways_gateway_17__EVAL;
  wire  gateways_gateway_17__EVAL_0;
  wire  gateways_gateway_17__EVAL_1;
  wire  gateways_gateway_17__EVAL_2;
  wire  gateways_gateway_17__EVAL_3;
  wire  gateways_gateway_17__EVAL_4;
  wire  _EVAL_826;
  wire  _EVAL_827;
  wire  _EVAL_828;
  wire  gateways_gateway_55__EVAL;
  wire  gateways_gateway_55__EVAL_0;
  wire  gateways_gateway_55__EVAL_1;
  wire  gateways_gateway_55__EVAL_2;
  wire  gateways_gateway_55__EVAL_3;
  wire  gateways_gateway_55__EVAL_4;
  wire [31:0] _EVAL_832;
  wire  _EVAL_834;
  wire  _EVAL_837;
  wire  _EVAL_838;
  wire  _EVAL_840;
  wire  _EVAL_841;
  wire  _EVAL_842;
  wire  _EVAL_844;
  wire [31:0] _EVAL_845;
  wire  _EVAL_847;
  wire  gateways_gateway_86__EVAL;
  wire  gateways_gateway_86__EVAL_0;
  wire  gateways_gateway_86__EVAL_1;
  wire  gateways_gateway_86__EVAL_2;
  wire  gateways_gateway_86__EVAL_3;
  wire  gateways_gateway_86__EVAL_4;
  wire  _EVAL_848;
  wire  _EVAL_849;
  wire  _EVAL_850;
  wire  _EVAL_851;
  reg [2:0] _EVAL_853;
  reg [2:0] _EVAL_854;
  wire  _EVAL_855;
  wire  _EVAL_856;
  wire  _EVAL_858;
  wire  _EVAL_860;
  wire  _EVAL_862;
  reg [2:0] _EVAL_865;
  wire  gateways_gateway_30__EVAL;
  wire  gateways_gateway_30__EVAL_0;
  wire  gateways_gateway_30__EVAL_1;
  wire  gateways_gateway_30__EVAL_2;
  wire  gateways_gateway_30__EVAL_3;
  wire  gateways_gateway_30__EVAL_4;
  wire  _EVAL_868;
  wire  _EVAL_869;
  wire  _EVAL_870;
  wire  _EVAL_871;
  reg  _EVAL_872;
  wire  _EVAL_873;
  wire  _EVAL_876;
  wire  _EVAL_886;
  wire  _EVAL_889;
  wire  _EVAL_890;
  wire [31:0] _EVAL_892;
  wire [31:0] _EVAL_894;
  wire  _EVAL_899;
  reg  _EVAL_902;
  wire  _EVAL_903;
  wire  _EVAL_904;
  wire [31:0] _EVAL_905;
  wire  _EVAL_906;
  wire  gateways_gateway_108__EVAL;
  wire  gateways_gateway_108__EVAL_0;
  wire  gateways_gateway_108__EVAL_1;
  wire  gateways_gateway_108__EVAL_2;
  wire  gateways_gateway_108__EVAL_3;
  wire  gateways_gateway_108__EVAL_4;
  wire  _EVAL_907;
  wire  _EVAL_908;
  wire [18:0] _EVAL_909;
  wire  _EVAL_910;
  reg  _EVAL_911;
  wire  _EVAL_913;
  wire  _EVAL_916;
  wire  _EVAL_917;
  wire  _EVAL_918;
  wire  _EVAL_921;
  wire  _EVAL_925;
  reg [7:0] _EVAL_930;
  wire  _EVAL_933;
  reg [2:0] _EVAL_936;
  wire  _EVAL_937;
  wire  _EVAL_939;
  wire  _EVAL_944;
  reg [2:0] _EVAL_953;
  wire  _EVAL_954;
  wire  _EVAL_955;
  wire  _EVAL_956;
  wire [31:0] _EVAL_957;
  wire  _EVAL_959;
  wire  _EVAL_962;
  wire  _EVAL_963;
  wire  _EVAL_964;
  reg  _EVAL_965;
  reg [2:0] _EVAL_966;
  wire  _EVAL_967;
  wire [31:0] _EVAL_970;
  wire  _EVAL_973;
  wire  _EVAL_975;
  wire  gateways_gateway_114__EVAL;
  wire  gateways_gateway_114__EVAL_0;
  wire  gateways_gateway_114__EVAL_1;
  wire  gateways_gateway_114__EVAL_2;
  wire  gateways_gateway_114__EVAL_3;
  wire  gateways_gateway_114__EVAL_4;
  wire [31:0] _EVAL_978;
  wire  _EVAL_979;
  wire  _EVAL_980;
  wire [18:0] _EVAL_982;
  wire  _EVAL_987;
  wire  _EVAL_988;
  wire  _EVAL_989;
  wire  _EVAL_991;
  wire  _EVAL_992;
  wire  _EVAL_994;
  wire  _EVAL_995;
  wire  _EVAL_996;
  wire  _EVAL_997;
  wire [31:0] _EVAL_1000;
  wire  _EVAL_1002;
  reg [2:0] _EVAL_1005;
  wire [31:0] _EVAL_1008;
  wire [31:0] _EVAL_1009;
  wire  _EVAL_1010;
  wire  _EVAL_1011;
  wire  _EVAL_1012;
  wire  _EVAL_1014;
  wire  _EVAL_1015;
  wire [7:0] _EVAL_1016;
  wire  _EVAL_1017;
  wire  _EVAL_1020;
  wire  gateways_gateway_83__EVAL;
  wire  gateways_gateway_83__EVAL_0;
  wire  gateways_gateway_83__EVAL_1;
  wire  gateways_gateway_83__EVAL_2;
  wire  gateways_gateway_83__EVAL_3;
  wire  gateways_gateway_83__EVAL_4;
  wire  _EVAL_1021;
  wire  _EVAL_1022;
  wire  _EVAL_1023;
  wire  _EVAL_1024;
  wire  _EVAL_1026;
  reg [7:0] _EVAL_1030;
  wire  _EVAL_1031;
  wire  _EVAL_1032;
  wire  _EVAL_1033;
  wire  _EVAL_1034;
  wire [31:0] _EVAL_1036;
  wire  _EVAL_1039;
  wire  _EVAL_1040;
  wire  _EVAL_1043;
  wire  _EVAL_1046;
  wire  _EVAL_1051;
  wire  _EVAL_1052;
  wire  _EVAL_1053;
  wire  _EVAL_1056;
  wire  _EVAL_1057;
  wire  _EVAL_1061;
  wire  _EVAL_1065;
  wire  _EVAL_1066;
  wire [31:0] _EVAL_1071;
  wire  _EVAL_1072;
  wire  _EVAL_1074;
  wire [31:0] _EVAL_1076;
  wire  _EVAL_1081;
  reg [2:0] _EVAL_1085;
  wire  _EVAL_1086;
  wire  _EVAL_1087;
  wire [31:0] _EVAL_1088;
  wire  gateways_gateway_34__EVAL;
  wire  gateways_gateway_34__EVAL_0;
  wire  gateways_gateway_34__EVAL_1;
  wire  gateways_gateway_34__EVAL_2;
  wire  gateways_gateway_34__EVAL_3;
  wire  gateways_gateway_34__EVAL_4;
  wire  _EVAL_1089;
  wire  _EVAL_1090;
  wire [31:0] _EVAL_1093;
  wire  _EVAL_1094;
  wire  _EVAL_1096;
  reg [2:0] _EVAL_1099;
  wire  _EVAL_1101;
  wire  _EVAL_1102;
  wire  _EVAL_1103;
  wire  _EVAL_1112;
  reg  _EVAL_1116;
  wire  _EVAL_1118;
  reg  _EVAL_1120;
  wire  _EVAL_1122;
  reg  _EVAL_1127;
  wire [31:0] _EVAL_1130;
  wire  _EVAL_1133;
  reg [2:0] _EVAL_1134;
  wire  _EVAL_1135;
  reg  _EVAL_1138;
  wire  _EVAL_1140;
  wire  _EVAL_1143;
  wire  _EVAL_1144;
  wire  _EVAL_1146;
  reg  _EVAL_1147;
  wire  _EVAL_1148;
  wire  gateways_gateway_37__EVAL;
  wire  gateways_gateway_37__EVAL_0;
  wire  gateways_gateway_37__EVAL_1;
  wire  gateways_gateway_37__EVAL_2;
  wire  gateways_gateway_37__EVAL_3;
  wire  gateways_gateway_37__EVAL_4;
  wire  _EVAL_1151;
  wire  _EVAL_1153;
  wire  _EVAL_1158;
  wire  _EVAL_1164;
  wire [31:0] _EVAL_1167;
  wire  _EVAL_1170;
  wire  _EVAL_1171;
  wire  _EVAL_1172;
  wire  _EVAL_1174;
  reg  _EVAL_1175;
  wire  _EVAL_1178;
  wire  gateways_gateway_6__EVAL;
  wire  gateways_gateway_6__EVAL_0;
  wire  gateways_gateway_6__EVAL_1;
  wire  gateways_gateway_6__EVAL_2;
  wire  gateways_gateway_6__EVAL_3;
  wire  gateways_gateway_6__EVAL_4;
  wire  _EVAL_1180;
  wire  _EVAL_1181;
  wire  _EVAL_1182;
  wire  _EVAL_1183;
  wire  _EVAL_1184;
  wire  _EVAL_1187;
  wire  _EVAL_1190;
  wire  _EVAL_1191;
  wire  _EVAL_1193;
  wire  _EVAL_1195;
  reg [2:0] _EVAL_1199;
  wire  _EVAL_1202;
  wire  _EVAL_1203;
  wire  _EVAL_1209;
  wire  _EVAL_1211;
  wire  gateways_gateway_92__EVAL;
  wire  gateways_gateway_92__EVAL_0;
  wire  gateways_gateway_92__EVAL_1;
  wire  gateways_gateway_92__EVAL_2;
  wire  gateways_gateway_92__EVAL_3;
  wire  gateways_gateway_92__EVAL_4;
  wire  _EVAL_1218;
  wire  _EVAL_1220;
  wire  _EVAL_1222;
  wire  _EVAL_1224;
  wire  _EVAL_1237;
  wire  _EVAL_1238;
  wire  _EVAL_1239;
  wire [31:0] _EVAL_1241;
  wire  _EVAL_1243;
  wire  _EVAL_1248;
  wire  _EVAL_1250;
  wire  _EVAL_1251;
  reg [2:0] _EVAL_1252;
  wire  _EVAL_1254;
  wire  _EVAL_1255;
  wire  _EVAL_1257;
  wire  _EVAL_1263;
  wire  _EVAL_1264;
  wire  _EVAL_1267;
  reg [2:0] _EVAL_1268;
  wire  _EVAL_1269;
  reg  _EVAL_1270;
  wire  _EVAL_1274;
  wire  _EVAL_1278;
  wire  _EVAL_1280;
  wire  _EVAL_1281;
  wire  _EVAL_1282;
  reg [2:0] _EVAL_1283;
  wire  _EVAL_1286;
  wire  _EVAL_1288;
  wire  _EVAL_1292;
  reg [2:0] _EVAL_1293;
  wire [31:0] _EVAL_1299;
  wire  _EVAL_1301;
  wire  _EVAL_1303;
  wire  _EVAL_1304;
  wire  _EVAL_1307;
  wire  _EVAL_1308;
  wire  gateways_gateway_90__EVAL;
  wire  gateways_gateway_90__EVAL_0;
  wire  gateways_gateway_90__EVAL_1;
  wire  gateways_gateway_90__EVAL_2;
  wire  gateways_gateway_90__EVAL_3;
  wire  gateways_gateway_90__EVAL_4;
  wire [31:0] _EVAL_1310;
  wire  _EVAL_1311;
  wire  _EVAL_1314;
  wire [31:0] _EVAL_1315;
  wire  _EVAL_1320;
  wire  _EVAL_1325;
  wire  _EVAL_1328;
  wire  _EVAL_1333;
  wire  _EVAL_1336;
  wire  _EVAL_1338;
  wire  _EVAL_1339;
  reg [7:0] _EVAL_1340;
  reg [2:0] _EVAL_1341;
  wire  _EVAL_1342;
  wire  _EVAL_1343;
  wire  _EVAL_1346;
  reg  _EVAL_1347;
  wire  gateways_gateway_14__EVAL;
  wire  gateways_gateway_14__EVAL_0;
  wire  gateways_gateway_14__EVAL_1;
  wire  gateways_gateway_14__EVAL_2;
  wire  gateways_gateway_14__EVAL_3;
  wire  gateways_gateway_14__EVAL_4;
  wire  _EVAL_1349;
  wire  _EVAL_1354;
  reg [2:0] _EVAL_1358;
  wire  _EVAL_1359;
  wire  _EVAL_1364;
  reg  _EVAL_1365;
  wire  _EVAL_1366;
  wire  _EVAL_1367;
  reg  _EVAL_1368;
  reg  _EVAL_1369;
  wire  _EVAL_1371;
  wire [31:0] _EVAL_1374;
  wire  gateways_gateway_125__EVAL;
  wire  gateways_gateway_125__EVAL_0;
  wire  gateways_gateway_125__EVAL_1;
  wire  gateways_gateway_125__EVAL_2;
  wire  gateways_gateway_125__EVAL_3;
  wire  gateways_gateway_125__EVAL_4;
  reg [7:0] _EVAL_1380;
  wire  gateways_gateway_88__EVAL;
  wire  gateways_gateway_88__EVAL_0;
  wire  gateways_gateway_88__EVAL_1;
  wire  gateways_gateway_88__EVAL_2;
  wire  gateways_gateway_88__EVAL_3;
  wire  gateways_gateway_88__EVAL_4;
  wire  _EVAL_1382;
  wire  _EVAL_1385;
  reg  _EVAL_1392;
  wire [31:0] _EVAL_1395;
  wire  _EVAL_1396;
  wire  _EVAL_1398;
  wire  _EVAL_1401;
  reg [2:0] _EVAL_1407;
  wire [6:0] _EVAL_1408;
  wire [6:0] _EVAL_1411;
  wire  _EVAL_1413;
  wire  gateways_gateway_72__EVAL;
  wire  gateways_gateway_72__EVAL_0;
  wire  gateways_gateway_72__EVAL_1;
  wire  gateways_gateway_72__EVAL_2;
  wire  gateways_gateway_72__EVAL_3;
  wire  gateways_gateway_72__EVAL_4;
  wire [31:0] _EVAL_1415;
  reg  _EVAL_1417;
  wire  _EVAL_1418;
  wire  _EVAL_1419;
  wire  _EVAL_1422;
  wire  _EVAL_1426;
  wire  _EVAL_1428;
  wire  _EVAL_1430;
  wire  _EVAL_1433;
  reg  _EVAL_1434;
  wire  _EVAL_1435;
  wire  _EVAL_1438;
  wire  _EVAL_1439;
  wire  _EVAL_1440;
  wire [31:0] _EVAL_1441;
  wire  _EVAL_1443;
  wire  _EVAL_1444;
  wire  _EVAL_1446;
  wire  _EVAL_1447;
  wire  _EVAL_1451;
  wire  _EVAL_1452;
  reg [2:0] _EVAL_1459;
  wire  _EVAL_1466;
  reg  _EVAL_1467;
  wire  out_back__EVAL;
  wire [19:0] out_back__EVAL_0;
  wire [31:0] out_back__EVAL_1;
  wire  out_back__EVAL_2;
  wire [19:0] out_back__EVAL_3;
  wire  out_back__EVAL_4;
  wire [3:0] out_back__EVAL_5;
  wire [1:0] out_back__EVAL_6;
  wire  out_back__EVAL_7;
  wire  out_back__EVAL_8;
  wire [9:0] out_back__EVAL_9;
  wire [31:0] out_back__EVAL_10;
  wire [9:0] out_back__EVAL_11;
  wire [3:0] out_back__EVAL_12;
  wire  out_back__EVAL_13;
  wire [1:0] out_back__EVAL_14;
  wire  out_back__EVAL_15;
  wire  out_back__EVAL_16;
  reg [7:0] _EVAL_1471;
  wire  _EVAL_1472;
  wire  _EVAL_1473;
  wire  _EVAL_1476;
  wire  gateways_gateway_39__EVAL;
  wire  gateways_gateway_39__EVAL_0;
  wire  gateways_gateway_39__EVAL_1;
  wire  gateways_gateway_39__EVAL_2;
  wire  gateways_gateway_39__EVAL_3;
  wire  gateways_gateway_39__EVAL_4;
  wire  _EVAL_1480;
  wire [31:0] _EVAL_1481;
  wire  _EVAL_1482;
  wire  _EVAL_1483;
  wire  _EVAL_1485;
  wire  _EVAL_1486;
  wire  _EVAL_1488;
  wire  _EVAL_1489;
  wire [31:0] _EVAL_1496;
  wire  _EVAL_1499;
  wire  _EVAL_1500;
  wire  _EVAL_1504;
  wire  _EVAL_1505;
  wire  _EVAL_1506;
  reg  _EVAL_1507;
  wire  _EVAL_1509;
  wire  _EVAL_1510;
  wire  _EVAL_1512;
  wire  _EVAL_1516;
  reg [7:0] _EVAL_1517;
  wire  _EVAL_1518;
  wire  _EVAL_1520;
  wire  _EVAL_1521;
  reg  _EVAL_1524;
  reg [2:0] _EVAL_1527;
  reg [2:0] _EVAL_1528;
  wire  _EVAL_1529;
  wire  _EVAL_1532;
  wire  _EVAL_1534;
  wire  _EVAL_1535;
  wire  _EVAL_1536;
  wire  _EVAL_1537;
  wire  gateways_gateway_10__EVAL;
  wire  gateways_gateway_10__EVAL_0;
  wire  gateways_gateway_10__EVAL_1;
  wire  gateways_gateway_10__EVAL_2;
  wire  gateways_gateway_10__EVAL_3;
  wire  gateways_gateway_10__EVAL_4;
  wire  _EVAL_1539;
  wire  _EVAL_1540;
  wire  gateways_gateway_70__EVAL;
  wire  gateways_gateway_70__EVAL_0;
  wire  gateways_gateway_70__EVAL_1;
  wire  gateways_gateway_70__EVAL_2;
  wire  gateways_gateway_70__EVAL_3;
  wire  gateways_gateway_70__EVAL_4;
  wire  _EVAL_1541;
  wire  _EVAL_1542;
  wire  gateways_gateway_16__EVAL;
  wire  gateways_gateway_16__EVAL_0;
  wire  gateways_gateway_16__EVAL_1;
  wire  gateways_gateway_16__EVAL_2;
  wire  gateways_gateway_16__EVAL_3;
  wire  gateways_gateway_16__EVAL_4;
  wire  _EVAL_1544;
  wire  _EVAL_1547;
  reg [7:0] _EVAL_1548;
  wire  _EVAL_1549;
  wire  _EVAL_1550;
  wire  _EVAL_1554;
  wire  _EVAL_1555;
  wire  _EVAL_1560;
  wire  _EVAL_1564;
  reg  _EVAL_1565;
  wire [31:0] _EVAL_1568;
  reg [2:0] _EVAL_1569;
  reg  _EVAL_1576;
  wire  _EVAL_1578;
  wire  _EVAL_1579;
  wire [7:0] _EVAL_1587;
  wire  _EVAL_1591;
  wire  _EVAL_1592;
  wire  _EVAL_1593;
  wire  _EVAL_1594;
  wire  _EVAL_1595;
  wire  _EVAL_1596;
  wire  _EVAL_1597;
  wire  _EVAL_1601;
  wire [31:0] _EVAL_1605;
  wire [31:0] _EVAL_1608;
  wire  _EVAL_1610;
  wire  _EVAL_1613;
  wire  _EVAL_1618;
  reg [2:0] _EVAL_1621;
  wire  _EVAL_1622;
  wire [31:0] _EVAL_1623;
  wire  _EVAL_1624;
  wire  _EVAL_1627;
  wire  gateways_gateway_38__EVAL;
  wire  gateways_gateway_38__EVAL_0;
  wire  gateways_gateway_38__EVAL_1;
  wire  gateways_gateway_38__EVAL_2;
  wire  gateways_gateway_38__EVAL_3;
  wire  gateways_gateway_38__EVAL_4;
  wire  gateways_gateway_31__EVAL;
  wire  gateways_gateway_31__EVAL_0;
  wire  gateways_gateway_31__EVAL_1;
  wire  gateways_gateway_31__EVAL_2;
  wire  gateways_gateway_31__EVAL_3;
  wire  gateways_gateway_31__EVAL_4;
  wire  _EVAL_1630;
  wire  _EVAL_1631;
  reg [2:0] _EVAL_1634;
  wire  _EVAL_1637;
  reg  _EVAL_1638;
  wire  gateways_gateway_71__EVAL;
  wire  gateways_gateway_71__EVAL_0;
  wire  gateways_gateway_71__EVAL_1;
  wire  gateways_gateway_71__EVAL_2;
  wire  gateways_gateway_71__EVAL_3;
  wire  gateways_gateway_71__EVAL_4;
  wire  _EVAL_1644;
  wire  _EVAL_1645;
  reg [2:0] _EVAL_1647;
  wire  _EVAL_1649;
  reg [2:0] _EVAL_1655;
  wire  _EVAL_1657;
  wire  _EVAL_1658;
  wire [31:0] _EVAL_1659;
  wire [31:0] _EVAL_1661;
  wire  _EVAL_1662;
  wire  _EVAL_1664;
  wire  _EVAL_1666;
  wire  gateways_gateway_77__EVAL;
  wire  gateways_gateway_77__EVAL_0;
  wire  gateways_gateway_77__EVAL_1;
  wire  gateways_gateway_77__EVAL_2;
  wire  gateways_gateway_77__EVAL_3;
  wire  gateways_gateway_77__EVAL_4;
  wire  _EVAL_1670;
  reg  _EVAL_1673;
  wire  _EVAL_1674;
  wire  _EVAL_1677;
  wire [31:0] _EVAL_1678;
  wire  _EVAL_1680;
  wire  _EVAL_1681;
  wire  _EVAL_1683;
  wire  _EVAL_1684;
  reg [2:0] _EVAL_1687;
  wire  _EVAL_1688;
  wire  _EVAL_1689;
  reg [2:0] _EVAL_1692;
  reg [2:0] _EVAL_1695;
  wire [7:0] _EVAL_1696;
  wire  _EVAL_1697;
  wire  _EVAL_1698;
  wire  _EVAL_1700;
  wire  gateways_gateway_61__EVAL;
  wire  gateways_gateway_61__EVAL_0;
  wire  gateways_gateway_61__EVAL_1;
  wire  gateways_gateway_61__EVAL_2;
  wire  gateways_gateway_61__EVAL_3;
  wire  gateways_gateway_61__EVAL_4;
  wire  gateways_gateway_59__EVAL;
  wire  gateways_gateway_59__EVAL_0;
  wire  gateways_gateway_59__EVAL_1;
  wire  gateways_gateway_59__EVAL_2;
  wire  gateways_gateway_59__EVAL_3;
  wire  gateways_gateway_59__EVAL_4;
  wire [31:0] _EVAL_1702;
  wire  _EVAL_1707;
  reg  _EVAL_1710;
  wire  _EVAL_1711;
  wire  _EVAL_1712;
  wire  _EVAL_1715;
  wire  gateways_gateway_15__EVAL;
  wire  gateways_gateway_15__EVAL_0;
  wire  gateways_gateway_15__EVAL_1;
  wire  gateways_gateway_15__EVAL_2;
  wire  gateways_gateway_15__EVAL_3;
  wire  gateways_gateway_15__EVAL_4;
  wire  _EVAL_1718;
  wire  _EVAL_1720;
  wire  _EVAL_1722;
  wire [7:0] _EVAL_1723;
  wire  _EVAL_1729;
  wire  _EVAL_1731;
  wire  _EVAL_1733;
  wire  _EVAL_1738;
  wire  _EVAL_1739;
  wire  _EVAL_1740;
  wire  _EVAL_1741;
  reg [2:0] _EVAL_1745;
  wire  gateways_gateway_105__EVAL;
  wire  gateways_gateway_105__EVAL_0;
  wire  gateways_gateway_105__EVAL_1;
  wire  gateways_gateway_105__EVAL_2;
  wire  gateways_gateway_105__EVAL_3;
  wire  gateways_gateway_105__EVAL_4;
  reg  _EVAL_1749;
  wire  _EVAL_1750;
  wire  _EVAL_1751;
  wire  _EVAL_1752;
  wire  _EVAL_1754;
  wire  _EVAL_1755;
  wire  _EVAL_1757;
  reg [2:0] _EVAL_1758;
  wire  _EVAL_1761;
  wire  _EVAL_1762;
  wire  _EVAL_1763;
  wire  _EVAL_1764;
  wire  _EVAL_1765;
  wire  _EVAL_1768;
  wire  _EVAL_1769;
  reg [2:0] _EVAL_1771;
  wire  _EVAL_1773;
  reg  _EVAL_1774;
  wire [31:0] _EVAL_1779;
  wire  _EVAL_1780;
  wire  _EVAL_1781;
  wire  _EVAL_1783;
  wire  _EVAL_1785;
  wire  _EVAL_1787;
  wire  _EVAL_1788;
  reg [2:0] _EVAL_1789;
  wire  _EVAL_1792;
  wire  _EVAL_1793;
  wire  _EVAL_1794;
  reg [2:0] _EVAL_1796;
  wire  _EVAL_1797;
  wire  _EVAL_1799;
  wire  _EVAL_1801;
  reg [2:0] _EVAL_1805;
  wire  gateways_gateway_115__EVAL;
  wire  gateways_gateway_115__EVAL_0;
  wire  gateways_gateway_115__EVAL_1;
  wire  gateways_gateway_115__EVAL_2;
  wire  gateways_gateway_115__EVAL_3;
  wire  gateways_gateway_115__EVAL_4;
  wire  _EVAL_1809;
  wire  _EVAL_1812;
  wire  _EVAL_1813;
  wire  _EVAL_1815;
  wire  gateways_gateway_98__EVAL;
  wire  gateways_gateway_98__EVAL_0;
  wire  gateways_gateway_98__EVAL_1;
  wire  gateways_gateway_98__EVAL_2;
  wire  gateways_gateway_98__EVAL_3;
  wire  gateways_gateway_98__EVAL_4;
  wire  _EVAL_1822;
  wire  _EVAL_1824;
  wire  gateways_gateway_49__EVAL;
  wire  gateways_gateway_49__EVAL_0;
  wire  gateways_gateway_49__EVAL_1;
  wire  gateways_gateway_49__EVAL_2;
  wire  gateways_gateway_49__EVAL_3;
  wire  gateways_gateway_49__EVAL_4;
  wire  _EVAL_1826;
  wire  _EVAL_1828;
  wire  _EVAL_1830;
  wire  _EVAL_1832;
  wire  _EVAL_1833;
  reg [2:0] _EVAL_1843;
  reg  _EVAL_1847;
  wire  _EVAL_1852;
  wire  _EVAL_1853;
  wire [31:0] _EVAL_1854;
  wire  _EVAL_1855;
  wire  _EVAL_1857;
  wire  gateways_gateway_119__EVAL;
  wire  gateways_gateway_119__EVAL_0;
  wire  gateways_gateway_119__EVAL_1;
  wire  gateways_gateway_119__EVAL_2;
  wire  gateways_gateway_119__EVAL_3;
  wire  gateways_gateway_119__EVAL_4;
  wire  gateways_gateway_112__EVAL;
  wire  gateways_gateway_112__EVAL_0;
  wire  gateways_gateway_112__EVAL_1;
  wire  gateways_gateway_112__EVAL_2;
  wire  gateways_gateway_112__EVAL_3;
  wire  gateways_gateway_112__EVAL_4;
  wire [27:0] _EVAL_1866;
  wire  _EVAL_1867;
  wire  _EVAL_1869;
  wire [31:0] _EVAL_1871;
  reg  _EVAL_1872;
  wire  _EVAL_1875;
  reg [2:0] _EVAL_1876;
  wire  _EVAL_1877;
  wire  _EVAL_1879;
  wire  _EVAL_1880;
  wire [31:0] _EVAL_1882;
  wire  _EVAL_1884;
  wire  _EVAL_1886;
  wire  gateways_gateway_3__EVAL;
  wire  gateways_gateway_3__EVAL_0;
  wire  gateways_gateway_3__EVAL_1;
  wire  gateways_gateway_3__EVAL_2;
  wire  gateways_gateway_3__EVAL_3;
  wire  gateways_gateway_3__EVAL_4;
  wire  _EVAL_1890;
  wire  _EVAL_1892;
  wire  _EVAL_1896;
  wire  gateways_gateway_124__EVAL;
  wire  gateways_gateway_124__EVAL_0;
  wire  gateways_gateway_124__EVAL_1;
  wire  gateways_gateway_124__EVAL_2;
  wire  gateways_gateway_124__EVAL_3;
  wire  gateways_gateway_124__EVAL_4;
  wire  _EVAL_1899;
  wire  _EVAL_1900;
  wire  _EVAL_1902;
  wire  gateways_gateway_21__EVAL;
  wire  gateways_gateway_21__EVAL_0;
  wire  gateways_gateway_21__EVAL_1;
  wire  gateways_gateway_21__EVAL_2;
  wire  gateways_gateway_21__EVAL_3;
  wire  gateways_gateway_21__EVAL_4;
  wire  _EVAL_1903;
  wire  _EVAL_1904;
  wire  _EVAL_1905;
  wire  _EVAL_1907;
  wire  _EVAL_1912;
  wire  gateways_gateway_33__EVAL;
  wire  gateways_gateway_33__EVAL_0;
  wire  gateways_gateway_33__EVAL_1;
  wire  gateways_gateway_33__EVAL_2;
  wire  gateways_gateway_33__EVAL_3;
  wire  gateways_gateway_33__EVAL_4;
  wire  _EVAL_1918;
  wire  _EVAL_1920;
  wire  gateways_gateway_110__EVAL;
  wire  gateways_gateway_110__EVAL_0;
  wire  gateways_gateway_110__EVAL_1;
  wire  gateways_gateway_110__EVAL_2;
  wire  gateways_gateway_110__EVAL_3;
  wire  gateways_gateway_110__EVAL_4;
  wire  _EVAL_1923;
  wire  gateways_gateway_9__EVAL;
  wire  gateways_gateway_9__EVAL_0;
  wire  gateways_gateway_9__EVAL_1;
  wire  gateways_gateway_9__EVAL_2;
  wire  gateways_gateway_9__EVAL_3;
  wire  gateways_gateway_9__EVAL_4;
  reg [6:0] _EVAL_1925;
  reg  _EVAL_1928;
  wire [31:0] _EVAL_1932;
  wire  _EVAL_1935;
  wire  gateways_gateway_51__EVAL;
  wire  gateways_gateway_51__EVAL_0;
  wire  gateways_gateway_51__EVAL_1;
  wire  gateways_gateway_51__EVAL_2;
  wire  gateways_gateway_51__EVAL_3;
  wire  gateways_gateway_51__EVAL_4;
  reg  _EVAL_1937;
  wire  _EVAL_1942;
  reg  _EVAL_1944;
  wire  _EVAL_1946;
  reg  _EVAL_1948;
  wire  _EVAL_1949;
  wire  gateways_gateway_97__EVAL;
  wire  gateways_gateway_97__EVAL_0;
  wire  gateways_gateway_97__EVAL_1;
  wire  gateways_gateway_97__EVAL_2;
  wire  gateways_gateway_97__EVAL_3;
  wire  gateways_gateway_97__EVAL_4;
  wire  _EVAL_1952;
  wire  _EVAL_1953;
  wire  _EVAL_1954;
  wire  _EVAL_1956;
  wire  _EVAL_1957;
  wire  gateways_gateway_123__EVAL;
  wire  gateways_gateway_123__EVAL_0;
  wire  gateways_gateway_123__EVAL_1;
  wire  gateways_gateway_123__EVAL_2;
  wire  gateways_gateway_123__EVAL_3;
  wire  gateways_gateway_123__EVAL_4;
  wire  _EVAL_1960;
  wire  _EVAL_1962;
  reg [2:0] _EVAL_1963;
  reg  _EVAL_1964;
  wire [31:0] _EVAL_1966;
  reg [2:0] _EVAL_1968;
  wire  _EVAL_1969;
  wire  _EVAL_1972;
  wire  _EVAL_1973;
  wire  _EVAL_1976;
  wire  _EVAL_1985;
  wire  _EVAL_1987;
  reg [2:0] _EVAL_1988;
  wire  _EVAL_1990;
  wire [15:0] _EVAL_1994;
  wire [31:0] _EVAL_1997;
  wire  _EVAL_1998;
  reg [2:0] _EVAL_2004;
  wire  _EVAL_2005;
  wire  _EVAL_2008;
  wire  _EVAL_2009;
  wire  _EVAL_2011;
  reg [2:0] _EVAL_2012;
  wire  _EVAL_2015;
  wire  _EVAL_2017;
  wire  _EVAL_2018;
  wire  _EVAL_2019;
  wire [31:0] _EVAL_2020;
  wire  _EVAL_2021;
  wire  _EVAL_2023;
  wire  _EVAL_2027;
  wire  gateways_gateway_104__EVAL;
  wire  gateways_gateway_104__EVAL_0;
  wire  gateways_gateway_104__EVAL_1;
  wire  gateways_gateway_104__EVAL_2;
  wire  gateways_gateway_104__EVAL_3;
  wire  gateways_gateway_104__EVAL_4;
  wire  _EVAL_2028;
  reg [2:0] _EVAL_2030;
  wire  gateways_gateway_81__EVAL;
  wire  gateways_gateway_81__EVAL_0;
  wire  gateways_gateway_81__EVAL_1;
  wire  gateways_gateway_81__EVAL_2;
  wire  gateways_gateway_81__EVAL_3;
  wire  gateways_gateway_81__EVAL_4;
  wire [31:0] _EVAL_2034;
  wire  _EVAL_2035;
  wire  _EVAL_2043;
  wire  gateways_gateway_78__EVAL;
  wire  gateways_gateway_78__EVAL_0;
  wire  gateways_gateway_78__EVAL_1;
  wire  gateways_gateway_78__EVAL_2;
  wire  gateways_gateway_78__EVAL_3;
  wire  gateways_gateway_78__EVAL_4;
  wire  _EVAL_2049;
  wire  _EVAL_2053;
  wire  _EVAL_2054;
  wire  _EVAL_2055;
  wire [31:0] _EVAL_2059;
  wire [31:0] _EVAL_2060;
  wire  _EVAL_2061;
  wire [31:0] _EVAL_2062;
  wire  gateways_gateway_69__EVAL;
  wire  gateways_gateway_69__EVAL_0;
  wire  gateways_gateway_69__EVAL_1;
  wire  gateways_gateway_69__EVAL_2;
  wire  gateways_gateway_69__EVAL_3;
  wire  gateways_gateway_69__EVAL_4;
  wire  gateways_gateway_101__EVAL;
  wire  gateways_gateway_101__EVAL_0;
  wire  gateways_gateway_101__EVAL_1;
  wire  gateways_gateway_101__EVAL_2;
  wire  gateways_gateway_101__EVAL_3;
  wire  gateways_gateway_101__EVAL_4;
  wire  _EVAL_2064;
  wire  gateways_gateway__EVAL;
  wire  gateways_gateway__EVAL_0;
  wire  gateways_gateway__EVAL_1;
  wire  gateways_gateway__EVAL_2;
  wire  gateways_gateway__EVAL_3;
  wire  gateways_gateway__EVAL_4;
  wire [31:0] _EVAL_2069;
  reg [7:0] _EVAL_2070;
  wire  _EVAL_2074;
  wire  _EVAL_2075;
  wire  _EVAL_2077;
  wire [31:0] _EVAL_2078;
  reg [2:0] _EVAL_2079;
  wire  _EVAL_2080;
  wire  _EVAL_2083;
  wire [2:0] _EVAL_2084;
  wire  _EVAL_2087;
  wire  _EVAL_2088;
  wire  _EVAL_2090;
  wire  _EVAL_2094;
  wire [31:0] _EVAL_2095;
  wire  _EVAL_2097;
  wire  _EVAL_2098;
  wire  _EVAL_2099;
  wire [31:0] _EVAL_2102;
  wire  _EVAL_2103;
  wire  _EVAL_2106;
  wire  gateways_gateway_27__EVAL;
  wire  gateways_gateway_27__EVAL_0;
  wire  gateways_gateway_27__EVAL_1;
  wire  gateways_gateway_27__EVAL_2;
  wire  gateways_gateway_27__EVAL_3;
  wire  gateways_gateway_27__EVAL_4;
  wire  _EVAL_2113;
  wire [7:0] _EVAL_2114;
  wire  _EVAL_2119;
  reg [7:0] _EVAL_2121;
  wire  _EVAL_2122;
  wire  _EVAL_2123;
  wire  _EVAL_2130;
  wire  _EVAL_2131;
  wire  _EVAL_2132;
  wire  _EVAL_2133;
  wire  _EVAL_2134;
  wire [31:0] _EVAL_2140;
  wire  _EVAL_2142;
  reg  _EVAL_2143;
  wire  _EVAL_2144;
  wire  _EVAL_2145;
  wire  _EVAL_2147;
  wire  _EVAL_2148;
  wire  _EVAL_2149;
  wire  _EVAL_2150;
  wire  _EVAL_2152;
  reg  _EVAL_2153;
  wire  _EVAL_2155;
  wire  _EVAL_2159;
  reg  _EVAL_2160;
  reg  _EVAL_2165;
  wire  gateways_gateway_76__EVAL;
  wire  gateways_gateway_76__EVAL_0;
  wire  gateways_gateway_76__EVAL_1;
  wire  gateways_gateway_76__EVAL_2;
  wire  gateways_gateway_76__EVAL_3;
  wire  gateways_gateway_76__EVAL_4;
  reg  _EVAL_2167;
  wire  _EVAL_2168;
  wire [31:0] _EVAL_2171;
  reg  _EVAL_2174;
  wire [31:0] _EVAL_2175;
  reg  _EVAL_2178;
  wire  _EVAL_2179;
  reg [2:0] _EVAL_2182;
  reg [2:0] _EVAL_2186;
  wire  _EVAL_2190;
  wire  _EVAL_2191;
  reg  _EVAL_2193;
  wire  _EVAL_2195;
  wire  _EVAL_2196;
  reg  _EVAL_2197;
  wire  _EVAL_2198;
  wire [31:0] _EVAL_2199;
  wire  gateways_gateway_82__EVAL;
  wire  gateways_gateway_82__EVAL_0;
  wire  gateways_gateway_82__EVAL_1;
  wire  gateways_gateway_82__EVAL_2;
  wire  gateways_gateway_82__EVAL_3;
  wire  gateways_gateway_82__EVAL_4;
  wire  _EVAL_2202;
  wire [31:0] _EVAL_2204;
  wire [31:0] _EVAL_2205;
  wire  _EVAL_2206;
  reg [2:0] _EVAL_2211;
  wire  _EVAL_2216;
  wire  _EVAL_2217;
  wire  _EVAL_2218;
  wire  _EVAL_2220;
  reg  _EVAL_2221;
  wire  _EVAL_2222;
  wire  gateways_gateway_94__EVAL;
  wire  gateways_gateway_94__EVAL_0;
  wire  gateways_gateway_94__EVAL_1;
  wire  gateways_gateway_94__EVAL_2;
  wire  gateways_gateway_94__EVAL_3;
  wire  gateways_gateway_94__EVAL_4;
  wire  _EVAL_2224;
  wire [31:0] _EVAL_2226;
  wire  _EVAL_2227;
  wire [31:0] _EVAL_2230;
  wire  _EVAL_2231;
  wire  _EVAL_2233;
  wire  _EVAL_2234;
  wire  _EVAL_2236;
  wire  _EVAL_2249;
  wire  _EVAL_2251;
  wire  _EVAL_2252;
  wire  _EVAL_2253;
  wire  _EVAL_2254;
  wire  _EVAL_2257;
  reg [2:0] _EVAL_2262;
  wire  _EVAL_2263;
  wire  _EVAL_2264;
  reg  _EVAL_2268;
  wire  _EVAL_2270;
  wire  _EVAL_2274;
  wire [31:0] _EVAL_2275;
  wire  _EVAL_2276;
  wire  _EVAL_2279;
  reg [2:0] _EVAL_2281;
  wire  _EVAL_2282;
  wire [31:0] _EVAL_2284;
  wire [31:0] _EVAL_2285;
  wire  gateways_gateway_47__EVAL;
  wire  gateways_gateway_47__EVAL_0;
  wire  gateways_gateway_47__EVAL_1;
  wire  gateways_gateway_47__EVAL_2;
  wire  gateways_gateway_47__EVAL_3;
  wire  gateways_gateway_47__EVAL_4;
  wire  _EVAL_2289;
  wire  _EVAL_2294;
  wire [126:0] _EVAL_2296;
  reg  _EVAL_2297;
  wire  _EVAL_2298;
  wire [31:0] _EVAL_2300;
  wire  _EVAL_2303;
  reg [2:0] _EVAL_2306;
  wire  _EVAL_2308;
  reg [2:0] _EVAL_2309;
  wire  _EVAL_2312;
  wire  _EVAL_2313;
  wire [31:0] _EVAL_2314;
  wire  _EVAL_2315;
  wire  _EVAL_2316;
  wire  _EVAL_2318;
  wire  _EVAL_2320;
  wire  _EVAL_2321;
  wire  _EVAL_2322;
  wire  _EVAL_2327;
  wire  _EVAL_2328;
  wire  _EVAL_2329;
  wire  _EVAL_2337;
  wire  _EVAL_2341;
  wire  _EVAL_2342;
  reg  _EVAL_2344;
  wire  _EVAL_2345;
  wire  _EVAL_2346;
  wire  _EVAL_2347;
  wire  _EVAL_2348;
  wire  _EVAL_2349;
  wire  _EVAL_2350;
  wire [3:0] _EVAL_2352;
  wire  _EVAL_2354;
  wire [31:0] _EVAL_2361;
  wire  _EVAL_2362;
  wire  _EVAL_2366;
  wire  _EVAL_2369;
  reg  _EVAL_2370;
  wire  _EVAL_2375;
  wire [127:0] _EVAL_2377;
  wire  _EVAL_2378;
  wire [7:0] _EVAL_2379;
  wire  _EVAL_2380;
  reg [2:0] _EVAL_2384;
  wire [31:0] _EVAL_2385;
  wire [31:0] _EVAL_2386;
  wire  _EVAL_2389;
  wire [31:0] _EVAL_2391;
  wire  gateways_gateway_54__EVAL;
  wire  gateways_gateway_54__EVAL_0;
  wire  gateways_gateway_54__EVAL_1;
  wire  gateways_gateway_54__EVAL_2;
  wire  gateways_gateway_54__EVAL_3;
  wire  gateways_gateway_54__EVAL_4;
  wire  _EVAL_2392;
  reg  _EVAL_2396;
  wire  _EVAL_2397;
  wire  _EVAL_2399;
  wire  _EVAL_2403;
  wire  _EVAL_2406;
  wire  _EVAL_2408;
  wire  _EVAL_2410;
  wire  gateways_gateway_118__EVAL;
  wire  gateways_gateway_118__EVAL_0;
  wire  gateways_gateway_118__EVAL_1;
  wire  gateways_gateway_118__EVAL_2;
  wire  gateways_gateway_118__EVAL_3;
  wire  gateways_gateway_118__EVAL_4;
  wire  _EVAL_2415;
  wire  _EVAL_2417;
  reg [7:0] _EVAL_2418;
  wire  _EVAL_2425;
  reg  _EVAL_2427;
  wire  _EVAL_2428;
  wire  _EVAL_2431;
  wire  gateways_gateway_120__EVAL;
  wire  gateways_gateway_120__EVAL_0;
  wire  gateways_gateway_120__EVAL_1;
  wire  gateways_gateway_120__EVAL_2;
  wire  gateways_gateway_120__EVAL_3;
  wire  gateways_gateway_120__EVAL_4;
  wire  gateways_gateway_99__EVAL;
  wire  gateways_gateway_99__EVAL_0;
  wire  gateways_gateway_99__EVAL_1;
  wire  gateways_gateway_99__EVAL_2;
  wire  gateways_gateway_99__EVAL_3;
  wire  gateways_gateway_99__EVAL_4;
  wire  _EVAL_2438;
  wire  _EVAL_2439;
  wire [19:0] _EVAL_2440;
  wire  _EVAL_2441;
  wire  _EVAL_2444;
  wire  gateways_gateway_75__EVAL;
  wire  gateways_gateway_75__EVAL_0;
  wire  gateways_gateway_75__EVAL_1;
  wire  gateways_gateway_75__EVAL_2;
  wire  gateways_gateway_75__EVAL_3;
  wire  gateways_gateway_75__EVAL_4;
  wire  gateways_gateway_73__EVAL;
  wire  gateways_gateway_73__EVAL_0;
  wire  gateways_gateway_73__EVAL_1;
  wire  gateways_gateway_73__EVAL_2;
  wire  gateways_gateway_73__EVAL_3;
  wire  gateways_gateway_73__EVAL_4;
  wire [30:0] _EVAL_2450;
  wire [31:0] _EVAL_2451;
  wire  _EVAL_2453;
  wire  _EVAL_2454;
  wire  _EVAL_2455;
  wire  _EVAL_2460;
  wire  _EVAL_2462;
  wire  _EVAL_2465;
  reg [2:0] _EVAL_2466;
  wire [31:0] _EVAL_2469;
  wire [18:0] _EVAL_2472;
  wire  gateways_gateway_53__EVAL;
  wire  gateways_gateway_53__EVAL_0;
  wire  gateways_gateway_53__EVAL_1;
  wire  gateways_gateway_53__EVAL_2;
  wire  gateways_gateway_53__EVAL_3;
  wire  gateways_gateway_53__EVAL_4;
  wire  _EVAL_2473;
  wire  _EVAL_2474;
  wire  _EVAL_2476;
  reg [2:0] _EVAL_2477;
  wire [25:0] _EVAL_2478;
  wire  _EVAL_2479;
  wire  _EVAL_2482;
  wire  _EVAL_2483;
  wire  _EVAL_2484;
  wire [31:0] _EVAL_2486;
  reg  _EVAL_2488;
  wire  _EVAL_2490;
  wire  _EVAL_2492;
  wire  _EVAL_2494;
  wire  _EVAL_2498;
  wire  _EVAL_2499;
  reg  _EVAL_2502;
  wire  _EVAL_2503;
  reg  _EVAL_2509;
  wire  _EVAL_2511;
  wire  _EVAL_2515;
  wire  _EVAL_2517;
  reg [2:0] _EVAL_2518;
  wire [7:0] _EVAL_2520;
  wire  _EVAL_2521;
  wire  _EVAL_2525;
  wire  _EVAL_2527;
  wire  _EVAL_2530;
  reg [2:0] _EVAL_2531;
  wire  _EVAL_2533;
  wire  _EVAL_2534;
  wire  _EVAL_2537;
  wire  gateways_gateway_23__EVAL;
  wire  gateways_gateway_23__EVAL_0;
  wire  gateways_gateway_23__EVAL_1;
  wire  gateways_gateway_23__EVAL_2;
  wire  gateways_gateway_23__EVAL_3;
  wire  gateways_gateway_23__EVAL_4;
  wire  _EVAL_2542;
  wire [31:0] _EVAL_2549;
  wire  _EVAL_2554;
  wire  _EVAL_2555;
  wire  _EVAL_2556;
  wire  _EVAL_2557;
  wire  _EVAL_2558;
  wire  _EVAL_2559;
  wire  _EVAL_2561;
  wire  _EVAL_2565;
  wire  _EVAL_2568;
  wire  gateways_gateway_100__EVAL;
  wire  gateways_gateway_100__EVAL_0;
  wire  gateways_gateway_100__EVAL_1;
  wire  gateways_gateway_100__EVAL_2;
  wire  gateways_gateway_100__EVAL_3;
  wire  gateways_gateway_100__EVAL_4;
  reg [2:0] _EVAL_2575;
  wire [31:0] _EVAL_2576;
  wire  _EVAL_2577;
  reg [2:0] _EVAL_2580;
  wire  _EVAL_2586;
  wire  _EVAL_2589;
  wire  _EVAL_2593;
  wire  gateways_gateway_126__EVAL;
  wire  gateways_gateway_126__EVAL_0;
  wire  gateways_gateway_126__EVAL_1;
  wire  gateways_gateway_126__EVAL_2;
  wire  gateways_gateway_126__EVAL_3;
  wire  gateways_gateway_126__EVAL_4;
  wire  _EVAL_2601;
  wire  _EVAL_2604;
  wire  _EVAL_2607;
  wire  _EVAL_2612;
  wire  _EVAL_2615;
  wire  _EVAL_2616;
  wire  _EVAL_2617;
  reg  _EVAL_2618;
  wire  _EVAL_2619;
  reg [2:0] _EVAL_2621;
  wire  _EVAL_2622;
  wire  _EVAL_2623;
  wire  _EVAL_2624;
  wire  _EVAL_2626;
  reg  _EVAL_2627;
  wire [31:0] _EVAL_2628;
  wire  _EVAL_2629;
  wire  gateways_gateway_117__EVAL;
  wire  gateways_gateway_117__EVAL_0;
  wire  gateways_gateway_117__EVAL_1;
  wire  gateways_gateway_117__EVAL_2;
  wire  gateways_gateway_117__EVAL_3;
  wire  gateways_gateway_117__EVAL_4;
  wire  _EVAL_2632;
  wire  _EVAL_2633;
  reg [2:0] _EVAL_2637;
  wire [31:0] _EVAL_2639;
  wire  _EVAL_2649;
  wire [31:0] _EVAL_2650;
  wire  _EVAL_2651;
  wire  _EVAL_2653;
  wire [31:0] _EVAL_2654;
  reg  _EVAL_2655;
  wire  _EVAL_2658;
  wire  _EVAL_2659;
  wire  _EVAL_2660;
  wire  _EVAL_2661;
  wire [31:0] _EVAL_2663;
  wire  gateways_gateway_63__EVAL;
  wire  gateways_gateway_63__EVAL_0;
  wire  gateways_gateway_63__EVAL_1;
  wire  gateways_gateway_63__EVAL_2;
  wire  gateways_gateway_63__EVAL_3;
  wire  gateways_gateway_63__EVAL_4;
  wire  _EVAL_2667;
  reg  _EVAL_2668;
  wire  _EVAL_2671;
  wire  _EVAL_2672;
  wire  _EVAL_2676;
  wire [2:0] fanin__EVAL;
  wire [2:0] fanin__EVAL_0;
  wire [2:0] fanin__EVAL_1;
  wire [2:0] fanin__EVAL_2;
  wire [2:0] fanin__EVAL_3;
  wire [2:0] fanin__EVAL_4;
  wire [2:0] fanin__EVAL_5;
  wire [2:0] fanin__EVAL_6;
  wire [2:0] fanin__EVAL_7;
  wire [2:0] fanin__EVAL_8;
  wire [2:0] fanin__EVAL_9;
  wire [2:0] fanin__EVAL_10;
  wire [2:0] fanin__EVAL_11;
  wire [2:0] fanin__EVAL_12;
  wire [2:0] fanin__EVAL_13;
  wire [2:0] fanin__EVAL_14;
  wire [2:0] fanin__EVAL_15;
  wire [2:0] fanin__EVAL_16;
  wire [2:0] fanin__EVAL_17;
  wire [2:0] fanin__EVAL_18;
  wire [2:0] fanin__EVAL_19;
  wire [2:0] fanin__EVAL_20;
  wire [2:0] fanin__EVAL_21;
  wire [2:0] fanin__EVAL_22;
  wire [2:0] fanin__EVAL_23;
  wire [2:0] fanin__EVAL_24;
  wire [2:0] fanin__EVAL_25;
  wire [2:0] fanin__EVAL_26;
  wire [2:0] fanin__EVAL_27;
  wire [2:0] fanin__EVAL_28;
  wire [2:0] fanin__EVAL_29;
  wire [2:0] fanin__EVAL_30;
  wire [2:0] fanin__EVAL_31;
  wire [2:0] fanin__EVAL_32;
  wire [2:0] fanin__EVAL_33;
  wire [2:0] fanin__EVAL_34;
  wire [2:0] fanin__EVAL_35;
  wire [2:0] fanin__EVAL_36;
  wire [2:0] fanin__EVAL_37;
  wire [2:0] fanin__EVAL_38;
  wire [2:0] fanin__EVAL_39;
  wire [2:0] fanin__EVAL_40;
  wire [2:0] fanin__EVAL_41;
  wire [2:0] fanin__EVAL_42;
  wire [2:0] fanin__EVAL_43;
  wire [2:0] fanin__EVAL_44;
  wire [2:0] fanin__EVAL_45;
  wire [2:0] fanin__EVAL_46;
  wire [2:0] fanin__EVAL_47;
  wire [126:0] fanin__EVAL_48;
  wire [2:0] fanin__EVAL_49;
  wire [2:0] fanin__EVAL_50;
  wire [2:0] fanin__EVAL_51;
  wire [2:0] fanin__EVAL_52;
  wire [2:0] fanin__EVAL_53;
  wire [2:0] fanin__EVAL_54;
  wire [2:0] fanin__EVAL_55;
  wire [2:0] fanin__EVAL_56;
  wire [2:0] fanin__EVAL_57;
  wire [2:0] fanin__EVAL_58;
  wire [2:0] fanin__EVAL_59;
  wire [2:0] fanin__EVAL_60;
  wire [2:0] fanin__EVAL_61;
  wire [2:0] fanin__EVAL_62;
  wire [2:0] fanin__EVAL_63;
  wire [2:0] fanin__EVAL_64;
  wire [2:0] fanin__EVAL_65;
  wire [2:0] fanin__EVAL_66;
  wire [2:0] fanin__EVAL_67;
  wire [2:0] fanin__EVAL_68;
  wire [2:0] fanin__EVAL_69;
  wire [2:0] fanin__EVAL_70;
  wire [2:0] fanin__EVAL_71;
  wire [2:0] fanin__EVAL_72;
  wire [2:0] fanin__EVAL_73;
  wire [2:0] fanin__EVAL_74;
  wire [2:0] fanin__EVAL_75;
  wire [2:0] fanin__EVAL_76;
  wire [2:0] fanin__EVAL_77;
  wire [2:0] fanin__EVAL_78;
  wire [2:0] fanin__EVAL_79;
  wire [2:0] fanin__EVAL_80;
  wire [2:0] fanin__EVAL_81;
  wire [2:0] fanin__EVAL_82;
  wire [2:0] fanin__EVAL_83;
  wire [2:0] fanin__EVAL_84;
  wire [2:0] fanin__EVAL_85;
  wire [6:0] fanin__EVAL_86;
  wire [2:0] fanin__EVAL_87;
  wire [2:0] fanin__EVAL_88;
  wire [2:0] fanin__EVAL_89;
  wire [2:0] fanin__EVAL_90;
  wire [2:0] fanin__EVAL_91;
  wire [2:0] fanin__EVAL_92;
  wire [2:0] fanin__EVAL_93;
  wire [2:0] fanin__EVAL_94;
  wire [2:0] fanin__EVAL_95;
  wire [2:0] fanin__EVAL_96;
  wire [2:0] fanin__EVAL_97;
  wire [2:0] fanin__EVAL_98;
  wire [2:0] fanin__EVAL_99;
  wire [2:0] fanin__EVAL_100;
  wire [2:0] fanin__EVAL_101;
  wire [2:0] fanin__EVAL_102;
  wire [2:0] fanin__EVAL_103;
  wire [2:0] fanin__EVAL_104;
  wire [2:0] fanin__EVAL_105;
  wire [2:0] fanin__EVAL_106;
  wire [2:0] fanin__EVAL_107;
  wire [2:0] fanin__EVAL_108;
  wire [2:0] fanin__EVAL_109;
  wire [2:0] fanin__EVAL_110;
  wire [2:0] fanin__EVAL_111;
  wire [2:0] fanin__EVAL_112;
  wire [2:0] fanin__EVAL_113;
  wire [2:0] fanin__EVAL_114;
  wire [2:0] fanin__EVAL_115;
  wire [2:0] fanin__EVAL_116;
  wire [2:0] fanin__EVAL_117;
  wire [2:0] fanin__EVAL_118;
  wire [2:0] fanin__EVAL_119;
  wire [2:0] fanin__EVAL_120;
  wire [2:0] fanin__EVAL_121;
  wire [2:0] fanin__EVAL_122;
  wire [2:0] fanin__EVAL_123;
  wire [2:0] fanin__EVAL_124;
  wire [2:0] fanin__EVAL_125;
  wire [2:0] fanin__EVAL_126;
  wire [2:0] fanin__EVAL_127;
  wire [2:0] fanin__EVAL_128;
  reg  _EVAL_2682;
  reg  _EVAL_2685;
  wire  _EVAL_2686;
  wire  _EVAL_2689;
  wire  _EVAL_2692;
  wire  _EVAL_2693;
  wire  gateways_gateway_29__EVAL;
  wire  gateways_gateway_29__EVAL_0;
  wire  gateways_gateway_29__EVAL_1;
  wire  gateways_gateway_29__EVAL_2;
  wire  gateways_gateway_29__EVAL_3;
  wire  gateways_gateway_29__EVAL_4;
  wire [15:0] _EVAL_2694;
  wire  _EVAL_2696;
  wire [6:0] _EVAL_2697;
  reg  _EVAL_2698;
  wire  _EVAL_2700;
  wire  _EVAL_2701;
  wire  gateways_gateway_79__EVAL;
  wire  gateways_gateway_79__EVAL_0;
  wire  gateways_gateway_79__EVAL_1;
  wire  gateways_gateway_79__EVAL_2;
  wire  gateways_gateway_79__EVAL_3;
  wire  gateways_gateway_79__EVAL_4;
  wire  _EVAL_2702;
  wire  _EVAL_2710;
  reg [2:0] _EVAL_2711;
  wire  _EVAL_2712;
  reg  _EVAL_2719;
  wire  _EVAL_2720;
  wire [31:0] _EVAL_2722;
  wire  _EVAL_2724;
  wire  _EVAL_2727;
  wire  _EVAL_2728;
  wire  _EVAL_2730;
  wire  _EVAL_2732;
  wire  _EVAL_2733;
  wire  _EVAL_2734;
  reg  _EVAL_2737;
  wire  _EVAL_2738;
  wire  _EVAL_2739;
  wire  _EVAL_2742;
  wire [7:0] _EVAL_2745;
  wire  _EVAL_2747;
  reg [2:0] _EVAL_2753;
  wire  gateways_gateway_106__EVAL;
  wire  gateways_gateway_106__EVAL_0;
  wire  gateways_gateway_106__EVAL_1;
  wire  gateways_gateway_106__EVAL_2;
  wire  gateways_gateway_106__EVAL_3;
  wire  gateways_gateway_106__EVAL_4;
  wire  _EVAL_2756;
  reg [6:0] _EVAL_2757;
  wire  gateways_gateway_121__EVAL;
  wire  gateways_gateway_121__EVAL_0;
  wire  gateways_gateway_121__EVAL_1;
  wire  gateways_gateway_121__EVAL_2;
  wire  gateways_gateway_121__EVAL_3;
  wire  gateways_gateway_121__EVAL_4;
  wire [127:0] _EVAL_2758;
  wire  _EVAL_2759;
  wire  _EVAL_2763;
  wire  _EVAL_2770;
  wire  _EVAL_2772;
  wire  _EVAL_2773;
  wire  _EVAL_2774;
  wire  _EVAL_2777;
  wire  _EVAL_2779;
  wire  _EVAL_2784;
  wire  _EVAL_2787;
  wire  _EVAL_2788;
  wire [31:0] _EVAL_2789;
  wire [31:0] _EVAL_2791;
  reg  _EVAL_2793;
  wire  _EVAL_2795;
  wire  _EVAL_2798;
  reg  _EVAL_2799;
  wire [31:0] _EVAL_2800;
  wire  _EVAL_2801;
  wire  _EVAL_2803;
  wire  _EVAL_2805;
  wire  _EVAL_2810;
  wire  _EVAL_2811;
  wire  _EVAL_2812;
  wire  _EVAL_2814;
  wire  _EVAL_2817;
  wire  _EVAL_2822;
  reg [2:0] _EVAL_2828;
  wire  _EVAL_2832;
  wire  _EVAL_2833;
  wire [31:0] _EVAL_2838;
  wire  _EVAL_2841;
  wire  _EVAL_2842;
  wire  _EVAL_2844;
  reg [2:0] _EVAL_2845;
  wire  _EVAL_2846;
  wire [31:0] _EVAL_2850;
  wire  _EVAL_2852;
  reg [2:0] _EVAL_2853;
  wire  _EVAL_2855;
  wire  _EVAL_2856;
  wire  _EVAL_2860;
  wire  _EVAL_2861;
  wire  _EVAL_2862;
  wire  _EVAL_2865;
  wire  _EVAL_2868;
  wire [31:0] _EVAL_2871;
  wire [31:0] _EVAL_2872;
  reg [2:0] _EVAL_2873;
  wire  _EVAL_2874;
  reg [7:0] _EVAL_2877;
  reg [2:0] _EVAL_2878;
  wire  _EVAL_2879;
  wire  _EVAL_2880;
  wire  _EVAL_2881;
  wire  _EVAL_2885;
  wire  _EVAL_2888;
  wire [14:0] _EVAL_2889;
  wire  _EVAL_2892;
  wire  _EVAL_2896;
  reg  _EVAL_2900;
  wire [62:0] _EVAL_2902;
  wire [27:0] _EVAL_2903;
  wire  _EVAL_2904;
  wire  _EVAL_2906;
  wire  _EVAL_2907;
  wire  _EVAL_2910;
  wire  gateways_gateway_35__EVAL;
  wire  gateways_gateway_35__EVAL_0;
  wire  gateways_gateway_35__EVAL_1;
  wire  gateways_gateway_35__EVAL_2;
  wire  gateways_gateway_35__EVAL_3;
  wire  gateways_gateway_35__EVAL_4;
  wire  _EVAL_2911;
  wire  _EVAL_2913;
  wire [7:0] _EVAL_2914;
  wire  _EVAL_2915;
  wire [127:0] _EVAL_2917;
  wire [31:0] _EVAL_2918;
  wire  gateways_gateway_74__EVAL;
  wire  gateways_gateway_74__EVAL_0;
  wire  gateways_gateway_74__EVAL_1;
  wire  gateways_gateway_74__EVAL_2;
  wire  gateways_gateway_74__EVAL_3;
  wire  gateways_gateway_74__EVAL_4;
  wire  _EVAL_2919;
  reg [2:0] _EVAL_2921;
  wire  _EVAL_2922;
  wire  gateways_gateway_66__EVAL;
  wire  gateways_gateway_66__EVAL_0;
  wire  gateways_gateway_66__EVAL_1;
  wire  gateways_gateway_66__EVAL_2;
  wire  gateways_gateway_66__EVAL_3;
  wire  gateways_gateway_66__EVAL_4;
  wire  _EVAL_2926;
  wire  _EVAL_2927;
  wire  _EVAL_2928;
  wire  _EVAL_2929;
  wire  _EVAL_2934;
  wire  gateways_gateway_56__EVAL;
  wire  gateways_gateway_56__EVAL_0;
  wire  gateways_gateway_56__EVAL_1;
  wire  gateways_gateway_56__EVAL_2;
  wire  gateways_gateway_56__EVAL_3;
  wire  gateways_gateway_56__EVAL_4;
  wire  _EVAL_2936;
  wire [31:0] _EVAL_2938;
  wire  _EVAL_2942;
  reg  _EVAL_2944;
  wire  _EVAL_2945;
  wire [31:0] _EVAL_2946;
  reg  _EVAL_2951;
  wire  _EVAL_2952;
  wire  _EVAL_2956;
  wire  _EVAL_2957;
  wire  gateways_gateway_107__EVAL;
  wire  gateways_gateway_107__EVAL_0;
  wire  gateways_gateway_107__EVAL_1;
  wire  gateways_gateway_107__EVAL_2;
  wire  gateways_gateway_107__EVAL_3;
  wire  gateways_gateway_107__EVAL_4;
  reg  _EVAL_2961;
  wire  gateways_gateway_8__EVAL;
  wire  gateways_gateway_8__EVAL_0;
  wire  gateways_gateway_8__EVAL_1;
  wire  gateways_gateway_8__EVAL_2;
  wire  gateways_gateway_8__EVAL_3;
  wire  gateways_gateway_8__EVAL_4;
  wire  _EVAL_2963;
  wire  _EVAL_2965;
  wire  _EVAL_2966;
  wire [31:0] _EVAL_2969;
  wire  _EVAL_2970;
  wire  _EVAL_2974;
  wire  _EVAL_2977;
  wire  _EVAL_2978;
  wire [31:0] _EVAL_2979;
  wire  _EVAL_2980;
  reg [2:0] _EVAL_2981;
  reg [2:0] _EVAL_2982;
  wire  _EVAL_2983;
  wire  _EVAL_2985;
  reg [2:0] _EVAL_2986;
  wire  _EVAL_2987;
  reg [2:0] _EVAL_2988;
  wire  _EVAL_2989;
  wire  _EVAL_2990;
  wire  _EVAL_2992;
  reg [2:0] _EVAL_2996;
  wire  gateways_gateway_11__EVAL;
  wire  gateways_gateway_11__EVAL_0;
  wire  gateways_gateway_11__EVAL_1;
  wire  gateways_gateway_11__EVAL_2;
  wire  gateways_gateway_11__EVAL_3;
  wire  gateways_gateway_11__EVAL_4;
  wire [9:0] _EVAL_2998;
  wire  _EVAL_2999;
  wire  _EVAL_3000;
  wire  _EVAL_3001;
  wire  _EVAL_3002;
  reg [2:0] _EVAL_3005;
  wire  _EVAL_3007;
  wire  gateways_gateway_12__EVAL;
  wire  gateways_gateway_12__EVAL_0;
  wire  gateways_gateway_12__EVAL_1;
  wire  gateways_gateway_12__EVAL_2;
  wire  gateways_gateway_12__EVAL_3;
  wire  gateways_gateway_12__EVAL_4;
  wire  _EVAL_3008;
  reg  _EVAL_3011;
  reg [2:0] _EVAL_3013;
  reg  _EVAL_3014;
  wire [127:0] _EVAL_3015;
  wire [31:0] _EVAL_3017;
  wire  _EVAL_3027;
  wire  _EVAL_3029;
  wire  _EVAL_3030;
  wire [31:0] _EVAL_3033;
  wire  _EVAL_3034;
  wire  _EVAL_3035;
  wire  _EVAL_3036;
  wire  _EVAL_3037;
  wire [7:0] _EVAL_3038;
  wire  _EVAL_3039;
  wire  _EVAL_3040;
  reg  _EVAL_3043;
  wire  _EVAL_3047;
  reg [2:0] _EVAL_3055;
  wire  _EVAL_3056;
  reg  _EVAL_3059;
  wire  _EVAL_3061;
  reg [2:0] _EVAL_3063;
  wire  _EVAL_3064;
  wire  _EVAL_3067;
  wire  _EVAL_3068;
  wire  _EVAL_3069;
  wire  _EVAL_3071;
  reg [2:0] _EVAL_3072;
  wire  _EVAL_3074;
  wire [31:0] _EVAL_3075;
  wire [31:0] _EVAL_3076;
  wire [31:0] _EVAL_3077;
  wire  gateways_gateway_57__EVAL;
  wire  gateways_gateway_57__EVAL_0;
  wire  gateways_gateway_57__EVAL_1;
  wire  gateways_gateway_57__EVAL_2;
  wire  gateways_gateway_57__EVAL_3;
  wire  gateways_gateway_57__EVAL_4;
  reg [2:0] _EVAL_3080;
  wire  _EVAL_3081;
  wire [31:0] _EVAL_3082;
  wire [31:0] _EVAL_3084;
  wire  _EVAL_3086;
  wire  _EVAL_3089;
  wire  _EVAL_3094;
  reg [2:0] _EVAL_3096;
  wire  _EVAL_3097;
  wire  _EVAL_3099;
  wire  _EVAL_3101;
  wire [31:0] _EVAL_3102;
  wire  _EVAL_3104;
  wire  _EVAL_3105;
  wire  _EVAL_3106;
  reg  _EVAL_3107;
  wire  _EVAL_3108;
  wire  gateways_gateway_43__EVAL;
  wire  gateways_gateway_43__EVAL_0;
  wire  gateways_gateway_43__EVAL_1;
  wire  gateways_gateway_43__EVAL_2;
  wire  gateways_gateway_43__EVAL_3;
  wire  gateways_gateway_43__EVAL_4;
  wire  gateways_gateway_4__EVAL;
  wire  gateways_gateway_4__EVAL_0;
  wire  gateways_gateway_4__EVAL_1;
  wire  gateways_gateway_4__EVAL_2;
  wire  gateways_gateway_4__EVAL_3;
  wire  gateways_gateway_4__EVAL_4;
  wire  _EVAL_3111;
  reg  _EVAL_3112;
  wire  _EVAL_3114;
  wire  _EVAL_3115;
  wire  _EVAL_3122;
  wire  _EVAL_3123;
  wire [31:0] _EVAL_3124;
  wire  gateways_gateway_36__EVAL;
  wire  gateways_gateway_36__EVAL_0;
  wire  gateways_gateway_36__EVAL_1;
  wire  gateways_gateway_36__EVAL_2;
  wire  gateways_gateway_36__EVAL_3;
  wire  gateways_gateway_36__EVAL_4;
  wire  _EVAL_3127;
  reg  _EVAL_3129;
  wire  _EVAL_3130;
  wire  _EVAL_3133;
  wire [31:0] _EVAL_3134;
  wire  _EVAL_3138;
  reg  _EVAL_3140;
  wire  _EVAL_3142;
  reg  _EVAL_3145;
  wire  _EVAL_3147;
  wire  _EVAL_3148;
  reg  _EVAL_3150;
  reg  _EVAL_3151;
  wire  _EVAL_3152;
  wire  _EVAL_3153;
  wire  _EVAL_3155;
  reg [2:0] _EVAL_3156;
  wire  _EVAL_3157;
  wire  _EVAL_3161;
  wire  _EVAL_3162;
  wire  _EVAL_3165;
  wire [31:0] _EVAL_3166;
  wire  _EVAL_3167;
  wire  _EVAL_3171;
  wire  _EVAL_3172;
  wire  gateways_gateway_5__EVAL;
  wire  gateways_gateway_5__EVAL_0;
  wire  gateways_gateway_5__EVAL_1;
  wire  gateways_gateway_5__EVAL_2;
  wire  gateways_gateway_5__EVAL_3;
  wire  gateways_gateway_5__EVAL_4;
  wire  _EVAL_3174;
  wire  _EVAL_3179;
  wire  gateways_gateway_18__EVAL;
  wire  gateways_gateway_18__EVAL_0;
  wire  gateways_gateway_18__EVAL_1;
  wire  gateways_gateway_18__EVAL_2;
  wire  gateways_gateway_18__EVAL_3;
  wire  gateways_gateway_18__EVAL_4;
  wire  _EVAL_3182;
  wire  _EVAL_3183;
  wire  _EVAL_3185;
  wire  _EVAL_3186;
  wire  _EVAL_3189;
  reg [2:0] _EVAL_3191;
  wire  _EVAL_3193;
  wire [31:0] _EVAL_3198;
  reg  _EVAL_3199;
  reg  _EVAL_3200;
  wire  _EVAL_3201;
  wire  _EVAL_3204;
  wire  _EVAL_3205;
  wire  _EVAL_3206;
  wire  _EVAL_3209;
  wire  _EVAL_3210;
  wire  _EVAL_3211;
  reg  _EVAL_3213;
  wire [9:0] _EVAL_3214;
  reg [2:0] _EVAL_3216;
  wire  _EVAL_3217;
  reg [2:0] _EVAL_3218;
  wire  _EVAL_3219;
  wire  _EVAL_3220;
  wire  _EVAL_3221;
  wire [7:0] _EVAL_3222;
  wire  _EVAL_3223;
  wire [31:0] _EVAL_3225;
  wire  gateways_gateway_50__EVAL;
  wire  gateways_gateway_50__EVAL_0;
  wire  gateways_gateway_50__EVAL_1;
  wire  gateways_gateway_50__EVAL_2;
  wire  gateways_gateway_50__EVAL_3;
  wire  gateways_gateway_50__EVAL_4;
  wire  _EVAL_3236;
  wire  _EVAL_3237;
  wire [15:0] _EVAL_3240;
  wire [7:0] _EVAL_3241;
  reg  _EVAL_3242;
  wire  _EVAL_3243;
  wire  _EVAL_3244;
  wire [7:0] _EVAL_3245;
  wire  _EVAL_3246;
  wire  _EVAL_3249;
  wire  _EVAL_3251;
  wire  _EVAL_3255;
  wire  _EVAL_3256;
  wire  _EVAL_3259;
  wire  _EVAL_3260;
  wire  _EVAL_3261;
  wire [31:0] _EVAL_3262;
  wire [27:0] _EVAL_3263;
  wire  gateways_gateway_60__EVAL;
  wire  gateways_gateway_60__EVAL_0;
  wire  gateways_gateway_60__EVAL_1;
  wire  gateways_gateway_60__EVAL_2;
  wire  gateways_gateway_60__EVAL_3;
  wire  gateways_gateway_60__EVAL_4;
  wire  _EVAL_3264;
  wire [7:0] _EVAL_3265;
  wire  _EVAL_3266;
  reg  _EVAL_3268;
  wire  _EVAL_3270;
  wire  _EVAL_3271;
  wire  _EVAL_3275;
  wire  _EVAL_3278;
  reg [2:0] _EVAL_3284;
  wire  _EVAL_3285;
  wire  _EVAL_3286;
  wire  _EVAL_3287;
  wire  _EVAL_3288;
  reg [2:0] _EVAL_3290;
  wire  _EVAL_3291;
  wire  _EVAL_3299;
  wire  _EVAL_3303;
  wire  gateways_gateway_95__EVAL;
  wire  gateways_gateway_95__EVAL_0;
  wire  gateways_gateway_95__EVAL_1;
  wire  gateways_gateway_95__EVAL_2;
  wire  gateways_gateway_95__EVAL_3;
  wire  gateways_gateway_95__EVAL_4;
  wire  _EVAL_3304;
  reg  _EVAL_3305;
  wire  _EVAL_3307;
  wire  _EVAL_3311;
  wire  _EVAL_3312;
  reg [2:0] _EVAL_3315;
  wire  _EVAL_3316;
  wire  _EVAL_3317;
  wire  _EVAL_3318;
  wire  _EVAL_3319;
  wire  _EVAL_3321;
  wire  _EVAL_3322;
  wire  gateways_gateway_13__EVAL;
  wire  gateways_gateway_13__EVAL_0;
  wire  gateways_gateway_13__EVAL_1;
  wire  gateways_gateway_13__EVAL_2;
  wire  gateways_gateway_13__EVAL_3;
  wire  gateways_gateway_13__EVAL_4;
  wire  _EVAL_3324;
  wire  _EVAL_3326;
  wire  _EVAL_3328;
  wire  _EVAL_3329;
  reg  _EVAL_3331;
  wire [31:0] _EVAL_3335;
  wire [31:0] _EVAL_3336;
  wire  _EVAL_3337;
  wire  _EVAL_3339;
  wire  _EVAL_3340;
  wire  _EVAL_3341;
  reg [2:0] _EVAL_3342;
  wire  _EVAL_3343;
  reg  _EVAL_3346;
  wire  _EVAL_3347;
  wire [127:0] _EVAL_3349;
  wire  _EVAL_3353;
  wire  _EVAL_3354;
  wire [7:0] _EVAL_3355;
  reg [2:0] _EVAL_3357;
  wire  _EVAL_3358;
  wire  _EVAL_3359;
  wire  _EVAL_3361;
  wire  _EVAL_3363;
  reg  _EVAL_3366;
  wire  _EVAL_3367;
  wire  _EVAL_3368;
  wire  gateways_gateway_20__EVAL;
  wire  gateways_gateway_20__EVAL_0;
  wire  gateways_gateway_20__EVAL_1;
  wire  gateways_gateway_20__EVAL_2;
  wire  gateways_gateway_20__EVAL_3;
  wire  gateways_gateway_20__EVAL_4;
  wire [31:0] _EVAL_3370;
  wire  _EVAL_3374;
  wire  _EVAL_3375;
  wire  _EVAL_3376;
  wire  _EVAL_3378;
  wire  _EVAL_3381;
  wire  _EVAL_3384;
  wire [31:0] _EVAL_3386;
  reg  _EVAL_3387;
  wire  _EVAL_3388;
  wire  _EVAL_3390;
  wire  _EVAL_3391;
  wire  _EVAL_3392;
  wire  _EVAL_3393;
  wire [31:0] _EVAL_3394;
  reg  _EVAL_3395;
  wire [31:0] _EVAL_3397;
  wire  _EVAL_3399;
  wire  _EVAL_3401;
  wire  _EVAL_3402;
  wire [31:0] _EVAL_3404;
  wire  _EVAL_3408;
  wire  _EVAL_3409;
  wire  _EVAL_3410;
  wire [7:0] _EVAL_3412;
  wire  _EVAL_3414;
  wire  _EVAL_3416;
  wire  _EVAL_3417;
  wire  _EVAL_3418;
  reg  _EVAL_3420;
  wire  _EVAL_3422;
  wire  _EVAL_3426;
  wire  gateways_gateway_25__EVAL;
  wire  gateways_gateway_25__EVAL_0;
  wire  gateways_gateway_25__EVAL_1;
  wire  gateways_gateway_25__EVAL_2;
  wire  gateways_gateway_25__EVAL_3;
  wire  gateways_gateway_25__EVAL_4;
  wire  _EVAL_3427;
  wire [31:0] _EVAL_3430;
  wire  _EVAL_3433;
  wire  _EVAL_3434;
  wire  _EVAL_3435;
  wire  _EVAL_3436;
  reg [2:0] _EVAL_3437;
  wire  _EVAL_3438;
  reg  _EVAL_3440;
  wire [31:0] _EVAL_3442;
  wire  _EVAL_3443;
  wire  _EVAL_3444;
  reg [2:0] _EVAL_3446;
  wire  _EVAL_3449;
  wire  _EVAL_3450;
  wire [31:0] _EVAL_3454;
  wire [31:0] _EVAL_3455;
  wire  _EVAL_3456;
  wire  _EVAL_3457;
  wire [31:0] _EVAL_3461;
  wire  _EVAL_3462;
  wire  _EVAL_3463;
  wire  _EVAL_3465;
  wire  _EVAL_3467;
  wire  gateways_gateway_19__EVAL;
  wire  gateways_gateway_19__EVAL_0;
  wire  gateways_gateway_19__EVAL_1;
  wire  gateways_gateway_19__EVAL_2;
  wire  gateways_gateway_19__EVAL_3;
  wire  gateways_gateway_19__EVAL_4;
  wire  _EVAL_3468;
  reg [2:0] _EVAL_3469;
  wire [31:0] _EVAL_3471;
  wire  _EVAL_3474;
  wire [6:0] _EVAL_3475;
  wire  _EVAL_3476;
  wire  _EVAL_3480;
  wire  _EVAL_3481;
  wire  _EVAL_3483;
  wire  _EVAL_3485;
  wire  _EVAL_3486;
  wire  _EVAL_3488;
  wire  _EVAL_3489;
  wire  _EVAL_3490;
  wire  _EVAL_3494;
  wire  _EVAL_3504;
  reg [2:0] _EVAL_3505;
  wire  gateways_gateway_32__EVAL;
  wire  gateways_gateway_32__EVAL_0;
  wire  gateways_gateway_32__EVAL_1;
  wire  gateways_gateway_32__EVAL_2;
  wire  gateways_gateway_32__EVAL_3;
  wire  gateways_gateway_32__EVAL_4;
  reg  _EVAL_3508;
  wire  _EVAL_3510;
  reg [2:0] _EVAL_3513;
  reg [2:0] _EVAL_3516;
  wire  _EVAL_3519;
  wire  _EVAL_3521;
  wire  _EVAL_3523;
  wire  _EVAL_3524;
  wire  _EVAL_3526;
  reg  _EVAL_3527;
  wire  _EVAL_3528;
  wire  _EVAL_3529;
  wire  _EVAL_3530;
  wire  _EVAL_3531;
  wire  _EVAL_3533;
  wire  _EVAL_3534;
  wire  _EVAL_3537;
  wire  _EVAL_3538;
  wire  _EVAL_3545;
  wire  _EVAL_3548;
  wire  _EVAL_3555;
  wire  _EVAL_3557;
  reg [2:0] _EVAL_3559;
  wire  _EVAL_3560;
  wire  _EVAL_3564;
  wire  _EVAL_3566;
  wire  _EVAL_3567;
  wire [31:0] _EVAL_3568;
  wire  _EVAL_3569;
  wire  _EVAL_3571;
  wire  _EVAL_3572;
  wire  _EVAL_3575;
  wire  _EVAL_3576;
  wire  _EVAL_3577;
  wire  _EVAL_3579;
  wire  _EVAL_3587;
  wire  _EVAL_3588;
  wire  gateways_gateway_67__EVAL;
  wire  gateways_gateway_67__EVAL_0;
  wire  gateways_gateway_67__EVAL_1;
  wire  gateways_gateway_67__EVAL_2;
  wire  gateways_gateway_67__EVAL_3;
  wire  gateways_gateway_67__EVAL_4;
  reg  _EVAL_3589;
  reg [2:0] _EVAL_3590;
  wire [31:0] _EVAL_3591;
  wire  _EVAL_3593;
  wire  _EVAL_3595;
  wire  _EVAL_3596;
  wire  _EVAL_3597;
  wire  _EVAL_3599;
  wire  _EVAL_3600;
  wire  _EVAL_3603;
  wire  gateways_gateway_93__EVAL;
  wire  gateways_gateway_93__EVAL_0;
  wire  gateways_gateway_93__EVAL_1;
  wire  gateways_gateway_93__EVAL_2;
  wire  gateways_gateway_93__EVAL_3;
  wire  gateways_gateway_93__EVAL_4;
  wire  _EVAL_3610;
  wire  _EVAL_3612;
  wire [27:0] _EVAL_3615;
  wire  _EVAL_3616;
  wire  _EVAL_3618;
  wire  _EVAL_3619;
  wire  _EVAL_3620;
  wire  gateways_gateway_52__EVAL;
  wire  gateways_gateway_52__EVAL_0;
  wire  gateways_gateway_52__EVAL_1;
  wire  gateways_gateway_52__EVAL_2;
  wire  gateways_gateway_52__EVAL_3;
  wire  gateways_gateway_52__EVAL_4;
  wire  _EVAL_3622;
  reg [2:0] _EVAL_3624;
  wire  _EVAL_3626;
  reg  _EVAL_3627;
  wire  _EVAL_3632;
  wire  _EVAL_3633;
  reg [2:0] _EVAL_3635;
  wire  _EVAL_3637;
  wire  _EVAL_3639;
  wire  _EVAL_3642;
  reg  _EVAL_3643;
  wire [9:0] _EVAL_3644;
  wire  _EVAL_3646;
  wire  _EVAL_3651;
  wire  _EVAL_3652;
  reg [2:0] _EVAL_3653;
  reg [7:0] _EVAL_3654;
  reg  _EVAL_3656;
  reg [2:0] _EVAL_3657;
  wire  _EVAL_3662;
  wire  _EVAL_3663;
  wire  gateways_gateway_109__EVAL;
  wire  gateways_gateway_109__EVAL_0;
  wire  gateways_gateway_109__EVAL_1;
  wire  gateways_gateway_109__EVAL_2;
  wire  gateways_gateway_109__EVAL_3;
  wire  gateways_gateway_109__EVAL_4;
  wire  _EVAL_3667;
  wire  _EVAL_3672;
  wire [31:0] _EVAL_3680;
  wire  _EVAL_3681;
  wire  _EVAL_3683;
  wire  _EVAL_3684;
  wire  _EVAL_3685;
  wire  _EVAL_3686;
  wire  gateways_gateway_64__EVAL;
  wire  gateways_gateway_64__EVAL_0;
  wire  gateways_gateway_64__EVAL_1;
  wire  gateways_gateway_64__EVAL_2;
  wire  gateways_gateway_64__EVAL_3;
  wire  gateways_gateway_64__EVAL_4;
  wire [31:0] _EVAL_3692;
  wire  _EVAL_3695;
  wire  _EVAL_3696;
  wire  _EVAL_3700;
  wire  _EVAL_3701;
  wire [6:0] _EVAL_3702;
  wire  _EVAL_3704;
  wire [31:0] _EVAL_3706;
  wire  _EVAL_3708;
  wire  gateways_gateway_80__EVAL;
  wire  gateways_gateway_80__EVAL_0;
  wire  gateways_gateway_80__EVAL_1;
  wire  gateways_gateway_80__EVAL_2;
  wire  gateways_gateway_80__EVAL_3;
  wire  gateways_gateway_80__EVAL_4;
  reg [2:0] _EVAL_3711;
  wire  gateways_gateway_85__EVAL;
  wire  gateways_gateway_85__EVAL_0;
  wire  gateways_gateway_85__EVAL_1;
  wire  gateways_gateway_85__EVAL_2;
  wire  gateways_gateway_85__EVAL_3;
  wire  gateways_gateway_85__EVAL_4;
  wire [31:0] _EVAL_3714;
  wire  _EVAL_3715;
  wire  _EVAL_3716;
  wire  _EVAL_3717;
  wire  _EVAL_3718;
  wire  _EVAL_3719;
  wire  _EVAL_3720;
  wire  _EVAL_3722;
  wire  _EVAL_3723;
  wire  _EVAL_3725;
  wire  _EVAL_3729;
  wire  _EVAL_3732;
  reg [2:0] _EVAL_3734;
  wire  _EVAL_3735;
  reg [2:0] _EVAL_3737;
  wire  _EVAL_3742;
  wire [31:0] _EVAL_3743;
  reg [2:0] _EVAL_3744;
  wire  _EVAL_3745;
  wire  _EVAL_3747;
  wire  _EVAL_3756;
  wire  _EVAL_3757;
  wire  gateways_gateway_48__EVAL;
  wire  gateways_gateway_48__EVAL_0;
  wire  gateways_gateway_48__EVAL_1;
  wire  gateways_gateway_48__EVAL_2;
  wire  gateways_gateway_48__EVAL_3;
  wire  gateways_gateway_48__EVAL_4;
  wire  _EVAL_3760;
  wire  _EVAL_3762;
  reg  _EVAL_3770;
  wire  _EVAL_3772;
  wire  _EVAL_3775;
  wire  _EVAL_3777;
  wire  _EVAL_3782;
  wire  _EVAL_3786;
  wire  _EVAL_3787;
  wire  _EVAL_3791;
  wire  _EVAL_3793;
  wire  _EVAL_3794;
  wire  _EVAL_3797;
  reg [2:0] _EVAL_3798;
  wire  _EVAL_3800;
  wire  _EVAL_3801;
  wire  _EVAL_3802;
  reg  _EVAL_3803;
  wire  _EVAL_3804;
  wire  _EVAL_3806;
  wire  _EVAL_3807;
  wire  _EVAL_3809;
  wire  _EVAL_3811;
  wire  gateways_gateway_26__EVAL;
  wire  gateways_gateway_26__EVAL_0;
  wire  gateways_gateway_26__EVAL_1;
  wire  gateways_gateway_26__EVAL_2;
  wire  gateways_gateway_26__EVAL_3;
  wire  gateways_gateway_26__EVAL_4;
  wire  _EVAL_3815;
  wire  _EVAL_3819;
  reg  _EVAL_3824;
  reg [2:0] _EVAL_3825;
  wire  _EVAL_3828;
  wire  _EVAL_3834;
  reg [2:0] _EVAL_3835;
  wire  _EVAL_3840;
  wire  gateways_gateway_65__EVAL;
  wire  gateways_gateway_65__EVAL_0;
  wire  gateways_gateway_65__EVAL_1;
  wire  gateways_gateway_65__EVAL_2;
  wire  gateways_gateway_65__EVAL_3;
  wire  gateways_gateway_65__EVAL_4;
  wire  gateways_gateway_62__EVAL;
  wire  gateways_gateway_62__EVAL_0;
  wire  gateways_gateway_62__EVAL_1;
  wire  gateways_gateway_62__EVAL_2;
  wire  gateways_gateway_62__EVAL_3;
  wire  gateways_gateway_62__EVAL_4;
  wire  _EVAL_3844;
  wire  _EVAL_3845;
  wire  _EVAL_3847;
  wire [31:0] _EVAL_3848;
  wire  _EVAL_3849;
  reg [7:0] _EVAL_3850;
  wire  _EVAL_3851;
  wire  _EVAL_3852;
  _EVAL_96 gateways_gateway_45 (
    ._EVAL(gateways_gateway_45__EVAL),
    ._EVAL_0(gateways_gateway_45__EVAL_0),
    ._EVAL_1(gateways_gateway_45__EVAL_1),
    ._EVAL_2(gateways_gateway_45__EVAL_2),
    ._EVAL_3(gateways_gateway_45__EVAL_3),
    ._EVAL_4(gateways_gateway_45__EVAL_4)
  );
  _EVAL_96 gateways_gateway_87 (
    ._EVAL(gateways_gateway_87__EVAL),
    ._EVAL_0(gateways_gateway_87__EVAL_0),
    ._EVAL_1(gateways_gateway_87__EVAL_1),
    ._EVAL_2(gateways_gateway_87__EVAL_2),
    ._EVAL_3(gateways_gateway_87__EVAL_3),
    ._EVAL_4(gateways_gateway_87__EVAL_4)
  );
  _EVAL_96 gateways_gateway_58 (
    ._EVAL(gateways_gateway_58__EVAL),
    ._EVAL_0(gateways_gateway_58__EVAL_0),
    ._EVAL_1(gateways_gateway_58__EVAL_1),
    ._EVAL_2(gateways_gateway_58__EVAL_2),
    ._EVAL_3(gateways_gateway_58__EVAL_3),
    ._EVAL_4(gateways_gateway_58__EVAL_4)
  );
  _EVAL_96 gateways_gateway_7 (
    ._EVAL(gateways_gateway_7__EVAL),
    ._EVAL_0(gateways_gateway_7__EVAL_0),
    ._EVAL_1(gateways_gateway_7__EVAL_1),
    ._EVAL_2(gateways_gateway_7__EVAL_2),
    ._EVAL_3(gateways_gateway_7__EVAL_3),
    ._EVAL_4(gateways_gateway_7__EVAL_4)
  );
  _EVAL_96 gateways_gateway_22 (
    ._EVAL(gateways_gateway_22__EVAL),
    ._EVAL_0(gateways_gateway_22__EVAL_0),
    ._EVAL_1(gateways_gateway_22__EVAL_1),
    ._EVAL_2(gateways_gateway_22__EVAL_2),
    ._EVAL_3(gateways_gateway_22__EVAL_3),
    ._EVAL_4(gateways_gateway_22__EVAL_4)
  );
  _EVAL_96 gateways_gateway_41 (
    ._EVAL(gateways_gateway_41__EVAL),
    ._EVAL_0(gateways_gateway_41__EVAL_0),
    ._EVAL_1(gateways_gateway_41__EVAL_1),
    ._EVAL_2(gateways_gateway_41__EVAL_2),
    ._EVAL_3(gateways_gateway_41__EVAL_3),
    ._EVAL_4(gateways_gateway_41__EVAL_4)
  );
  _EVAL_96 gateways_gateway_111 (
    ._EVAL(gateways_gateway_111__EVAL),
    ._EVAL_0(gateways_gateway_111__EVAL_0),
    ._EVAL_1(gateways_gateway_111__EVAL_1),
    ._EVAL_2(gateways_gateway_111__EVAL_2),
    ._EVAL_3(gateways_gateway_111__EVAL_3),
    ._EVAL_4(gateways_gateway_111__EVAL_4)
  );
  _EVAL_96 gateways_gateway_122 (
    ._EVAL(gateways_gateway_122__EVAL),
    ._EVAL_0(gateways_gateway_122__EVAL_0),
    ._EVAL_1(gateways_gateway_122__EVAL_1),
    ._EVAL_2(gateways_gateway_122__EVAL_2),
    ._EVAL_3(gateways_gateway_122__EVAL_3),
    ._EVAL_4(gateways_gateway_122__EVAL_4)
  );
  _EVAL_96 gateways_gateway_24 (
    ._EVAL(gateways_gateway_24__EVAL),
    ._EVAL_0(gateways_gateway_24__EVAL_0),
    ._EVAL_1(gateways_gateway_24__EVAL_1),
    ._EVAL_2(gateways_gateway_24__EVAL_2),
    ._EVAL_3(gateways_gateway_24__EVAL_3),
    ._EVAL_4(gateways_gateway_24__EVAL_4)
  );
  _EVAL_96 gateways_gateway_40 (
    ._EVAL(gateways_gateway_40__EVAL),
    ._EVAL_0(gateways_gateway_40__EVAL_0),
    ._EVAL_1(gateways_gateway_40__EVAL_1),
    ._EVAL_2(gateways_gateway_40__EVAL_2),
    ._EVAL_3(gateways_gateway_40__EVAL_3),
    ._EVAL_4(gateways_gateway_40__EVAL_4)
  );
  _EVAL_96 gateways_gateway_102 (
    ._EVAL(gateways_gateway_102__EVAL),
    ._EVAL_0(gateways_gateway_102__EVAL_0),
    ._EVAL_1(gateways_gateway_102__EVAL_1),
    ._EVAL_2(gateways_gateway_102__EVAL_2),
    ._EVAL_3(gateways_gateway_102__EVAL_3),
    ._EVAL_4(gateways_gateway_102__EVAL_4)
  );
  _EVAL_96 gateways_gateway_113 (
    ._EVAL(gateways_gateway_113__EVAL),
    ._EVAL_0(gateways_gateway_113__EVAL_0),
    ._EVAL_1(gateways_gateway_113__EVAL_1),
    ._EVAL_2(gateways_gateway_113__EVAL_2),
    ._EVAL_3(gateways_gateway_113__EVAL_3),
    ._EVAL_4(gateways_gateway_113__EVAL_4)
  );
  _EVAL_96 gateways_gateway_89 (
    ._EVAL(gateways_gateway_89__EVAL),
    ._EVAL_0(gateways_gateway_89__EVAL_0),
    ._EVAL_1(gateways_gateway_89__EVAL_1),
    ._EVAL_2(gateways_gateway_89__EVAL_2),
    ._EVAL_3(gateways_gateway_89__EVAL_3),
    ._EVAL_4(gateways_gateway_89__EVAL_4)
  );
  _EVAL_96 gateways_gateway_91 (
    ._EVAL(gateways_gateway_91__EVAL),
    ._EVAL_0(gateways_gateway_91__EVAL_0),
    ._EVAL_1(gateways_gateway_91__EVAL_1),
    ._EVAL_2(gateways_gateway_91__EVAL_2),
    ._EVAL_3(gateways_gateway_91__EVAL_3),
    ._EVAL_4(gateways_gateway_91__EVAL_4)
  );
  _EVAL_96 gateways_gateway_96 (
    ._EVAL(gateways_gateway_96__EVAL),
    ._EVAL_0(gateways_gateway_96__EVAL_0),
    ._EVAL_1(gateways_gateway_96__EVAL_1),
    ._EVAL_2(gateways_gateway_96__EVAL_2),
    ._EVAL_3(gateways_gateway_96__EVAL_3),
    ._EVAL_4(gateways_gateway_96__EVAL_4)
  );
  _EVAL_96 gateways_gateway_46 (
    ._EVAL(gateways_gateway_46__EVAL),
    ._EVAL_0(gateways_gateway_46__EVAL_0),
    ._EVAL_1(gateways_gateway_46__EVAL_1),
    ._EVAL_2(gateways_gateway_46__EVAL_2),
    ._EVAL_3(gateways_gateway_46__EVAL_3),
    ._EVAL_4(gateways_gateway_46__EVAL_4)
  );
  _EVAL_96 gateways_gateway_1 (
    ._EVAL(gateways_gateway_1__EVAL),
    ._EVAL_0(gateways_gateway_1__EVAL_0),
    ._EVAL_1(gateways_gateway_1__EVAL_1),
    ._EVAL_2(gateways_gateway_1__EVAL_2),
    ._EVAL_3(gateways_gateway_1__EVAL_3),
    ._EVAL_4(gateways_gateway_1__EVAL_4)
  );
  _EVAL_96 gateways_gateway_28 (
    ._EVAL(gateways_gateway_28__EVAL),
    ._EVAL_0(gateways_gateway_28__EVAL_0),
    ._EVAL_1(gateways_gateway_28__EVAL_1),
    ._EVAL_2(gateways_gateway_28__EVAL_2),
    ._EVAL_3(gateways_gateway_28__EVAL_3),
    ._EVAL_4(gateways_gateway_28__EVAL_4)
  );
  _EVAL_96 gateways_gateway_44 (
    ._EVAL(gateways_gateway_44__EVAL),
    ._EVAL_0(gateways_gateway_44__EVAL_0),
    ._EVAL_1(gateways_gateway_44__EVAL_1),
    ._EVAL_2(gateways_gateway_44__EVAL_2),
    ._EVAL_3(gateways_gateway_44__EVAL_3),
    ._EVAL_4(gateways_gateway_44__EVAL_4)
  );
  _EVAL_96 gateways_gateway_103 (
    ._EVAL(gateways_gateway_103__EVAL),
    ._EVAL_0(gateways_gateway_103__EVAL_0),
    ._EVAL_1(gateways_gateway_103__EVAL_1),
    ._EVAL_2(gateways_gateway_103__EVAL_2),
    ._EVAL_3(gateways_gateway_103__EVAL_3),
    ._EVAL_4(gateways_gateway_103__EVAL_4)
  );
  _EVAL_96 gateways_gateway_2 (
    ._EVAL(gateways_gateway_2__EVAL),
    ._EVAL_0(gateways_gateway_2__EVAL_0),
    ._EVAL_1(gateways_gateway_2__EVAL_1),
    ._EVAL_2(gateways_gateway_2__EVAL_2),
    ._EVAL_3(gateways_gateway_2__EVAL_3),
    ._EVAL_4(gateways_gateway_2__EVAL_4)
  );
  _EVAL_96 gateways_gateway_42 (
    ._EVAL(gateways_gateway_42__EVAL),
    ._EVAL_0(gateways_gateway_42__EVAL_0),
    ._EVAL_1(gateways_gateway_42__EVAL_1),
    ._EVAL_2(gateways_gateway_42__EVAL_2),
    ._EVAL_3(gateways_gateway_42__EVAL_3),
    ._EVAL_4(gateways_gateway_42__EVAL_4)
  );
  _EVAL_96 gateways_gateway_68 (
    ._EVAL(gateways_gateway_68__EVAL),
    ._EVAL_0(gateways_gateway_68__EVAL_0),
    ._EVAL_1(gateways_gateway_68__EVAL_1),
    ._EVAL_2(gateways_gateway_68__EVAL_2),
    ._EVAL_3(gateways_gateway_68__EVAL_3),
    ._EVAL_4(gateways_gateway_68__EVAL_4)
  );
  _EVAL_96 gateways_gateway_116 (
    ._EVAL(gateways_gateway_116__EVAL),
    ._EVAL_0(gateways_gateway_116__EVAL_0),
    ._EVAL_1(gateways_gateway_116__EVAL_1),
    ._EVAL_2(gateways_gateway_116__EVAL_2),
    ._EVAL_3(gateways_gateway_116__EVAL_3),
    ._EVAL_4(gateways_gateway_116__EVAL_4)
  );
  _EVAL_96 gateways_gateway_84 (
    ._EVAL(gateways_gateway_84__EVAL),
    ._EVAL_0(gateways_gateway_84__EVAL_0),
    ._EVAL_1(gateways_gateway_84__EVAL_1),
    ._EVAL_2(gateways_gateway_84__EVAL_2),
    ._EVAL_3(gateways_gateway_84__EVAL_3),
    ._EVAL_4(gateways_gateway_84__EVAL_4)
  );
  _EVAL_96 gateways_gateway_17 (
    ._EVAL(gateways_gateway_17__EVAL),
    ._EVAL_0(gateways_gateway_17__EVAL_0),
    ._EVAL_1(gateways_gateway_17__EVAL_1),
    ._EVAL_2(gateways_gateway_17__EVAL_2),
    ._EVAL_3(gateways_gateway_17__EVAL_3),
    ._EVAL_4(gateways_gateway_17__EVAL_4)
  );
  _EVAL_96 gateways_gateway_55 (
    ._EVAL(gateways_gateway_55__EVAL),
    ._EVAL_0(gateways_gateway_55__EVAL_0),
    ._EVAL_1(gateways_gateway_55__EVAL_1),
    ._EVAL_2(gateways_gateway_55__EVAL_2),
    ._EVAL_3(gateways_gateway_55__EVAL_3),
    ._EVAL_4(gateways_gateway_55__EVAL_4)
  );
  _EVAL_96 gateways_gateway_86 (
    ._EVAL(gateways_gateway_86__EVAL),
    ._EVAL_0(gateways_gateway_86__EVAL_0),
    ._EVAL_1(gateways_gateway_86__EVAL_1),
    ._EVAL_2(gateways_gateway_86__EVAL_2),
    ._EVAL_3(gateways_gateway_86__EVAL_3),
    ._EVAL_4(gateways_gateway_86__EVAL_4)
  );
  _EVAL_96 gateways_gateway_30 (
    ._EVAL(gateways_gateway_30__EVAL),
    ._EVAL_0(gateways_gateway_30__EVAL_0),
    ._EVAL_1(gateways_gateway_30__EVAL_1),
    ._EVAL_2(gateways_gateway_30__EVAL_2),
    ._EVAL_3(gateways_gateway_30__EVAL_3),
    ._EVAL_4(gateways_gateway_30__EVAL_4)
  );
  _EVAL_96 gateways_gateway_108 (
    ._EVAL(gateways_gateway_108__EVAL),
    ._EVAL_0(gateways_gateway_108__EVAL_0),
    ._EVAL_1(gateways_gateway_108__EVAL_1),
    ._EVAL_2(gateways_gateway_108__EVAL_2),
    ._EVAL_3(gateways_gateway_108__EVAL_3),
    ._EVAL_4(gateways_gateway_108__EVAL_4)
  );
  _EVAL_96 gateways_gateway_114 (
    ._EVAL(gateways_gateway_114__EVAL),
    ._EVAL_0(gateways_gateway_114__EVAL_0),
    ._EVAL_1(gateways_gateway_114__EVAL_1),
    ._EVAL_2(gateways_gateway_114__EVAL_2),
    ._EVAL_3(gateways_gateway_114__EVAL_3),
    ._EVAL_4(gateways_gateway_114__EVAL_4)
  );
  _EVAL_96 gateways_gateway_83 (
    ._EVAL(gateways_gateway_83__EVAL),
    ._EVAL_0(gateways_gateway_83__EVAL_0),
    ._EVAL_1(gateways_gateway_83__EVAL_1),
    ._EVAL_2(gateways_gateway_83__EVAL_2),
    ._EVAL_3(gateways_gateway_83__EVAL_3),
    ._EVAL_4(gateways_gateway_83__EVAL_4)
  );
  _EVAL_96 gateways_gateway_34 (
    ._EVAL(gateways_gateway_34__EVAL),
    ._EVAL_0(gateways_gateway_34__EVAL_0),
    ._EVAL_1(gateways_gateway_34__EVAL_1),
    ._EVAL_2(gateways_gateway_34__EVAL_2),
    ._EVAL_3(gateways_gateway_34__EVAL_3),
    ._EVAL_4(gateways_gateway_34__EVAL_4)
  );
  _EVAL_96 gateways_gateway_37 (
    ._EVAL(gateways_gateway_37__EVAL),
    ._EVAL_0(gateways_gateway_37__EVAL_0),
    ._EVAL_1(gateways_gateway_37__EVAL_1),
    ._EVAL_2(gateways_gateway_37__EVAL_2),
    ._EVAL_3(gateways_gateway_37__EVAL_3),
    ._EVAL_4(gateways_gateway_37__EVAL_4)
  );
  _EVAL_96 gateways_gateway_6 (
    ._EVAL(gateways_gateway_6__EVAL),
    ._EVAL_0(gateways_gateway_6__EVAL_0),
    ._EVAL_1(gateways_gateway_6__EVAL_1),
    ._EVAL_2(gateways_gateway_6__EVAL_2),
    ._EVAL_3(gateways_gateway_6__EVAL_3),
    ._EVAL_4(gateways_gateway_6__EVAL_4)
  );
  _EVAL_96 gateways_gateway_92 (
    ._EVAL(gateways_gateway_92__EVAL),
    ._EVAL_0(gateways_gateway_92__EVAL_0),
    ._EVAL_1(gateways_gateway_92__EVAL_1),
    ._EVAL_2(gateways_gateway_92__EVAL_2),
    ._EVAL_3(gateways_gateway_92__EVAL_3),
    ._EVAL_4(gateways_gateway_92__EVAL_4)
  );
  _EVAL_96 gateways_gateway_90 (
    ._EVAL(gateways_gateway_90__EVAL),
    ._EVAL_0(gateways_gateway_90__EVAL_0),
    ._EVAL_1(gateways_gateway_90__EVAL_1),
    ._EVAL_2(gateways_gateway_90__EVAL_2),
    ._EVAL_3(gateways_gateway_90__EVAL_3),
    ._EVAL_4(gateways_gateway_90__EVAL_4)
  );
  _EVAL_96 gateways_gateway_14 (
    ._EVAL(gateways_gateway_14__EVAL),
    ._EVAL_0(gateways_gateway_14__EVAL_0),
    ._EVAL_1(gateways_gateway_14__EVAL_1),
    ._EVAL_2(gateways_gateway_14__EVAL_2),
    ._EVAL_3(gateways_gateway_14__EVAL_3),
    ._EVAL_4(gateways_gateway_14__EVAL_4)
  );
  _EVAL_96 gateways_gateway_125 (
    ._EVAL(gateways_gateway_125__EVAL),
    ._EVAL_0(gateways_gateway_125__EVAL_0),
    ._EVAL_1(gateways_gateway_125__EVAL_1),
    ._EVAL_2(gateways_gateway_125__EVAL_2),
    ._EVAL_3(gateways_gateway_125__EVAL_3),
    ._EVAL_4(gateways_gateway_125__EVAL_4)
  );
  _EVAL_96 gateways_gateway_88 (
    ._EVAL(gateways_gateway_88__EVAL),
    ._EVAL_0(gateways_gateway_88__EVAL_0),
    ._EVAL_1(gateways_gateway_88__EVAL_1),
    ._EVAL_2(gateways_gateway_88__EVAL_2),
    ._EVAL_3(gateways_gateway_88__EVAL_3),
    ._EVAL_4(gateways_gateway_88__EVAL_4)
  );
  _EVAL_96 gateways_gateway_72 (
    ._EVAL(gateways_gateway_72__EVAL),
    ._EVAL_0(gateways_gateway_72__EVAL_0),
    ._EVAL_1(gateways_gateway_72__EVAL_1),
    ._EVAL_2(gateways_gateway_72__EVAL_2),
    ._EVAL_3(gateways_gateway_72__EVAL_3),
    ._EVAL_4(gateways_gateway_72__EVAL_4)
  );
  _EVAL_98 out_back (
    ._EVAL(out_back__EVAL),
    ._EVAL_0(out_back__EVAL_0),
    ._EVAL_1(out_back__EVAL_1),
    ._EVAL_2(out_back__EVAL_2),
    ._EVAL_3(out_back__EVAL_3),
    ._EVAL_4(out_back__EVAL_4),
    ._EVAL_5(out_back__EVAL_5),
    ._EVAL_6(out_back__EVAL_6),
    ._EVAL_7(out_back__EVAL_7),
    ._EVAL_8(out_back__EVAL_8),
    ._EVAL_9(out_back__EVAL_9),
    ._EVAL_10(out_back__EVAL_10),
    ._EVAL_11(out_back__EVAL_11),
    ._EVAL_12(out_back__EVAL_12),
    ._EVAL_13(out_back__EVAL_13),
    ._EVAL_14(out_back__EVAL_14),
    ._EVAL_15(out_back__EVAL_15),
    ._EVAL_16(out_back__EVAL_16)
  );
  _EVAL_96 gateways_gateway_39 (
    ._EVAL(gateways_gateway_39__EVAL),
    ._EVAL_0(gateways_gateway_39__EVAL_0),
    ._EVAL_1(gateways_gateway_39__EVAL_1),
    ._EVAL_2(gateways_gateway_39__EVAL_2),
    ._EVAL_3(gateways_gateway_39__EVAL_3),
    ._EVAL_4(gateways_gateway_39__EVAL_4)
  );
  _EVAL_96 gateways_gateway_10 (
    ._EVAL(gateways_gateway_10__EVAL),
    ._EVAL_0(gateways_gateway_10__EVAL_0),
    ._EVAL_1(gateways_gateway_10__EVAL_1),
    ._EVAL_2(gateways_gateway_10__EVAL_2),
    ._EVAL_3(gateways_gateway_10__EVAL_3),
    ._EVAL_4(gateways_gateway_10__EVAL_4)
  );
  _EVAL_96 gateways_gateway_70 (
    ._EVAL(gateways_gateway_70__EVAL),
    ._EVAL_0(gateways_gateway_70__EVAL_0),
    ._EVAL_1(gateways_gateway_70__EVAL_1),
    ._EVAL_2(gateways_gateway_70__EVAL_2),
    ._EVAL_3(gateways_gateway_70__EVAL_3),
    ._EVAL_4(gateways_gateway_70__EVAL_4)
  );
  _EVAL_96 gateways_gateway_16 (
    ._EVAL(gateways_gateway_16__EVAL),
    ._EVAL_0(gateways_gateway_16__EVAL_0),
    ._EVAL_1(gateways_gateway_16__EVAL_1),
    ._EVAL_2(gateways_gateway_16__EVAL_2),
    ._EVAL_3(gateways_gateway_16__EVAL_3),
    ._EVAL_4(gateways_gateway_16__EVAL_4)
  );
  _EVAL_96 gateways_gateway_38 (
    ._EVAL(gateways_gateway_38__EVAL),
    ._EVAL_0(gateways_gateway_38__EVAL_0),
    ._EVAL_1(gateways_gateway_38__EVAL_1),
    ._EVAL_2(gateways_gateway_38__EVAL_2),
    ._EVAL_3(gateways_gateway_38__EVAL_3),
    ._EVAL_4(gateways_gateway_38__EVAL_4)
  );
  _EVAL_96 gateways_gateway_31 (
    ._EVAL(gateways_gateway_31__EVAL),
    ._EVAL_0(gateways_gateway_31__EVAL_0),
    ._EVAL_1(gateways_gateway_31__EVAL_1),
    ._EVAL_2(gateways_gateway_31__EVAL_2),
    ._EVAL_3(gateways_gateway_31__EVAL_3),
    ._EVAL_4(gateways_gateway_31__EVAL_4)
  );
  _EVAL_96 gateways_gateway_71 (
    ._EVAL(gateways_gateway_71__EVAL),
    ._EVAL_0(gateways_gateway_71__EVAL_0),
    ._EVAL_1(gateways_gateway_71__EVAL_1),
    ._EVAL_2(gateways_gateway_71__EVAL_2),
    ._EVAL_3(gateways_gateway_71__EVAL_3),
    ._EVAL_4(gateways_gateway_71__EVAL_4)
  );
  _EVAL_96 gateways_gateway_77 (
    ._EVAL(gateways_gateway_77__EVAL),
    ._EVAL_0(gateways_gateway_77__EVAL_0),
    ._EVAL_1(gateways_gateway_77__EVAL_1),
    ._EVAL_2(gateways_gateway_77__EVAL_2),
    ._EVAL_3(gateways_gateway_77__EVAL_3),
    ._EVAL_4(gateways_gateway_77__EVAL_4)
  );
  _EVAL_96 gateways_gateway_61 (
    ._EVAL(gateways_gateway_61__EVAL),
    ._EVAL_0(gateways_gateway_61__EVAL_0),
    ._EVAL_1(gateways_gateway_61__EVAL_1),
    ._EVAL_2(gateways_gateway_61__EVAL_2),
    ._EVAL_3(gateways_gateway_61__EVAL_3),
    ._EVAL_4(gateways_gateway_61__EVAL_4)
  );
  _EVAL_96 gateways_gateway_59 (
    ._EVAL(gateways_gateway_59__EVAL),
    ._EVAL_0(gateways_gateway_59__EVAL_0),
    ._EVAL_1(gateways_gateway_59__EVAL_1),
    ._EVAL_2(gateways_gateway_59__EVAL_2),
    ._EVAL_3(gateways_gateway_59__EVAL_3),
    ._EVAL_4(gateways_gateway_59__EVAL_4)
  );
  _EVAL_96 gateways_gateway_15 (
    ._EVAL(gateways_gateway_15__EVAL),
    ._EVAL_0(gateways_gateway_15__EVAL_0),
    ._EVAL_1(gateways_gateway_15__EVAL_1),
    ._EVAL_2(gateways_gateway_15__EVAL_2),
    ._EVAL_3(gateways_gateway_15__EVAL_3),
    ._EVAL_4(gateways_gateway_15__EVAL_4)
  );
  _EVAL_96 gateways_gateway_105 (
    ._EVAL(gateways_gateway_105__EVAL),
    ._EVAL_0(gateways_gateway_105__EVAL_0),
    ._EVAL_1(gateways_gateway_105__EVAL_1),
    ._EVAL_2(gateways_gateway_105__EVAL_2),
    ._EVAL_3(gateways_gateway_105__EVAL_3),
    ._EVAL_4(gateways_gateway_105__EVAL_4)
  );
  _EVAL_96 gateways_gateway_115 (
    ._EVAL(gateways_gateway_115__EVAL),
    ._EVAL_0(gateways_gateway_115__EVAL_0),
    ._EVAL_1(gateways_gateway_115__EVAL_1),
    ._EVAL_2(gateways_gateway_115__EVAL_2),
    ._EVAL_3(gateways_gateway_115__EVAL_3),
    ._EVAL_4(gateways_gateway_115__EVAL_4)
  );
  _EVAL_96 gateways_gateway_98 (
    ._EVAL(gateways_gateway_98__EVAL),
    ._EVAL_0(gateways_gateway_98__EVAL_0),
    ._EVAL_1(gateways_gateway_98__EVAL_1),
    ._EVAL_2(gateways_gateway_98__EVAL_2),
    ._EVAL_3(gateways_gateway_98__EVAL_3),
    ._EVAL_4(gateways_gateway_98__EVAL_4)
  );
  _EVAL_96 gateways_gateway_49 (
    ._EVAL(gateways_gateway_49__EVAL),
    ._EVAL_0(gateways_gateway_49__EVAL_0),
    ._EVAL_1(gateways_gateway_49__EVAL_1),
    ._EVAL_2(gateways_gateway_49__EVAL_2),
    ._EVAL_3(gateways_gateway_49__EVAL_3),
    ._EVAL_4(gateways_gateway_49__EVAL_4)
  );
  _EVAL_96 gateways_gateway_119 (
    ._EVAL(gateways_gateway_119__EVAL),
    ._EVAL_0(gateways_gateway_119__EVAL_0),
    ._EVAL_1(gateways_gateway_119__EVAL_1),
    ._EVAL_2(gateways_gateway_119__EVAL_2),
    ._EVAL_3(gateways_gateway_119__EVAL_3),
    ._EVAL_4(gateways_gateway_119__EVAL_4)
  );
  _EVAL_96 gateways_gateway_112 (
    ._EVAL(gateways_gateway_112__EVAL),
    ._EVAL_0(gateways_gateway_112__EVAL_0),
    ._EVAL_1(gateways_gateway_112__EVAL_1),
    ._EVAL_2(gateways_gateway_112__EVAL_2),
    ._EVAL_3(gateways_gateway_112__EVAL_3),
    ._EVAL_4(gateways_gateway_112__EVAL_4)
  );
  _EVAL_96 gateways_gateway_3 (
    ._EVAL(gateways_gateway_3__EVAL),
    ._EVAL_0(gateways_gateway_3__EVAL_0),
    ._EVAL_1(gateways_gateway_3__EVAL_1),
    ._EVAL_2(gateways_gateway_3__EVAL_2),
    ._EVAL_3(gateways_gateway_3__EVAL_3),
    ._EVAL_4(gateways_gateway_3__EVAL_4)
  );
  _EVAL_96 gateways_gateway_124 (
    ._EVAL(gateways_gateway_124__EVAL),
    ._EVAL_0(gateways_gateway_124__EVAL_0),
    ._EVAL_1(gateways_gateway_124__EVAL_1),
    ._EVAL_2(gateways_gateway_124__EVAL_2),
    ._EVAL_3(gateways_gateway_124__EVAL_3),
    ._EVAL_4(gateways_gateway_124__EVAL_4)
  );
  _EVAL_96 gateways_gateway_21 (
    ._EVAL(gateways_gateway_21__EVAL),
    ._EVAL_0(gateways_gateway_21__EVAL_0),
    ._EVAL_1(gateways_gateway_21__EVAL_1),
    ._EVAL_2(gateways_gateway_21__EVAL_2),
    ._EVAL_3(gateways_gateway_21__EVAL_3),
    ._EVAL_4(gateways_gateway_21__EVAL_4)
  );
  _EVAL_96 gateways_gateway_33 (
    ._EVAL(gateways_gateway_33__EVAL),
    ._EVAL_0(gateways_gateway_33__EVAL_0),
    ._EVAL_1(gateways_gateway_33__EVAL_1),
    ._EVAL_2(gateways_gateway_33__EVAL_2),
    ._EVAL_3(gateways_gateway_33__EVAL_3),
    ._EVAL_4(gateways_gateway_33__EVAL_4)
  );
  _EVAL_96 gateways_gateway_110 (
    ._EVAL(gateways_gateway_110__EVAL),
    ._EVAL_0(gateways_gateway_110__EVAL_0),
    ._EVAL_1(gateways_gateway_110__EVAL_1),
    ._EVAL_2(gateways_gateway_110__EVAL_2),
    ._EVAL_3(gateways_gateway_110__EVAL_3),
    ._EVAL_4(gateways_gateway_110__EVAL_4)
  );
  _EVAL_96 gateways_gateway_9 (
    ._EVAL(gateways_gateway_9__EVAL),
    ._EVAL_0(gateways_gateway_9__EVAL_0),
    ._EVAL_1(gateways_gateway_9__EVAL_1),
    ._EVAL_2(gateways_gateway_9__EVAL_2),
    ._EVAL_3(gateways_gateway_9__EVAL_3),
    ._EVAL_4(gateways_gateway_9__EVAL_4)
  );
  _EVAL_96 gateways_gateway_51 (
    ._EVAL(gateways_gateway_51__EVAL),
    ._EVAL_0(gateways_gateway_51__EVAL_0),
    ._EVAL_1(gateways_gateway_51__EVAL_1),
    ._EVAL_2(gateways_gateway_51__EVAL_2),
    ._EVAL_3(gateways_gateway_51__EVAL_3),
    ._EVAL_4(gateways_gateway_51__EVAL_4)
  );
  _EVAL_96 gateways_gateway_97 (
    ._EVAL(gateways_gateway_97__EVAL),
    ._EVAL_0(gateways_gateway_97__EVAL_0),
    ._EVAL_1(gateways_gateway_97__EVAL_1),
    ._EVAL_2(gateways_gateway_97__EVAL_2),
    ._EVAL_3(gateways_gateway_97__EVAL_3),
    ._EVAL_4(gateways_gateway_97__EVAL_4)
  );
  _EVAL_96 gateways_gateway_123 (
    ._EVAL(gateways_gateway_123__EVAL),
    ._EVAL_0(gateways_gateway_123__EVAL_0),
    ._EVAL_1(gateways_gateway_123__EVAL_1),
    ._EVAL_2(gateways_gateway_123__EVAL_2),
    ._EVAL_3(gateways_gateway_123__EVAL_3),
    ._EVAL_4(gateways_gateway_123__EVAL_4)
  );
  _EVAL_96 gateways_gateway_104 (
    ._EVAL(gateways_gateway_104__EVAL),
    ._EVAL_0(gateways_gateway_104__EVAL_0),
    ._EVAL_1(gateways_gateway_104__EVAL_1),
    ._EVAL_2(gateways_gateway_104__EVAL_2),
    ._EVAL_3(gateways_gateway_104__EVAL_3),
    ._EVAL_4(gateways_gateway_104__EVAL_4)
  );
  _EVAL_96 gateways_gateway_81 (
    ._EVAL(gateways_gateway_81__EVAL),
    ._EVAL_0(gateways_gateway_81__EVAL_0),
    ._EVAL_1(gateways_gateway_81__EVAL_1),
    ._EVAL_2(gateways_gateway_81__EVAL_2),
    ._EVAL_3(gateways_gateway_81__EVAL_3),
    ._EVAL_4(gateways_gateway_81__EVAL_4)
  );
  _EVAL_96 gateways_gateway_78 (
    ._EVAL(gateways_gateway_78__EVAL),
    ._EVAL_0(gateways_gateway_78__EVAL_0),
    ._EVAL_1(gateways_gateway_78__EVAL_1),
    ._EVAL_2(gateways_gateway_78__EVAL_2),
    ._EVAL_3(gateways_gateway_78__EVAL_3),
    ._EVAL_4(gateways_gateway_78__EVAL_4)
  );
  _EVAL_96 gateways_gateway_69 (
    ._EVAL(gateways_gateway_69__EVAL),
    ._EVAL_0(gateways_gateway_69__EVAL_0),
    ._EVAL_1(gateways_gateway_69__EVAL_1),
    ._EVAL_2(gateways_gateway_69__EVAL_2),
    ._EVAL_3(gateways_gateway_69__EVAL_3),
    ._EVAL_4(gateways_gateway_69__EVAL_4)
  );
  _EVAL_96 gateways_gateway_101 (
    ._EVAL(gateways_gateway_101__EVAL),
    ._EVAL_0(gateways_gateway_101__EVAL_0),
    ._EVAL_1(gateways_gateway_101__EVAL_1),
    ._EVAL_2(gateways_gateway_101__EVAL_2),
    ._EVAL_3(gateways_gateway_101__EVAL_3),
    ._EVAL_4(gateways_gateway_101__EVAL_4)
  );
  _EVAL_96 gateways_gateway (
    ._EVAL(gateways_gateway__EVAL),
    ._EVAL_0(gateways_gateway__EVAL_0),
    ._EVAL_1(gateways_gateway__EVAL_1),
    ._EVAL_2(gateways_gateway__EVAL_2),
    ._EVAL_3(gateways_gateway__EVAL_3),
    ._EVAL_4(gateways_gateway__EVAL_4)
  );
  _EVAL_96 gateways_gateway_27 (
    ._EVAL(gateways_gateway_27__EVAL),
    ._EVAL_0(gateways_gateway_27__EVAL_0),
    ._EVAL_1(gateways_gateway_27__EVAL_1),
    ._EVAL_2(gateways_gateway_27__EVAL_2),
    ._EVAL_3(gateways_gateway_27__EVAL_3),
    ._EVAL_4(gateways_gateway_27__EVAL_4)
  );
  _EVAL_96 gateways_gateway_76 (
    ._EVAL(gateways_gateway_76__EVAL),
    ._EVAL_0(gateways_gateway_76__EVAL_0),
    ._EVAL_1(gateways_gateway_76__EVAL_1),
    ._EVAL_2(gateways_gateway_76__EVAL_2),
    ._EVAL_3(gateways_gateway_76__EVAL_3),
    ._EVAL_4(gateways_gateway_76__EVAL_4)
  );
  _EVAL_96 gateways_gateway_82 (
    ._EVAL(gateways_gateway_82__EVAL),
    ._EVAL_0(gateways_gateway_82__EVAL_0),
    ._EVAL_1(gateways_gateway_82__EVAL_1),
    ._EVAL_2(gateways_gateway_82__EVAL_2),
    ._EVAL_3(gateways_gateway_82__EVAL_3),
    ._EVAL_4(gateways_gateway_82__EVAL_4)
  );
  _EVAL_96 gateways_gateway_94 (
    ._EVAL(gateways_gateway_94__EVAL),
    ._EVAL_0(gateways_gateway_94__EVAL_0),
    ._EVAL_1(gateways_gateway_94__EVAL_1),
    ._EVAL_2(gateways_gateway_94__EVAL_2),
    ._EVAL_3(gateways_gateway_94__EVAL_3),
    ._EVAL_4(gateways_gateway_94__EVAL_4)
  );
  _EVAL_96 gateways_gateway_47 (
    ._EVAL(gateways_gateway_47__EVAL),
    ._EVAL_0(gateways_gateway_47__EVAL_0),
    ._EVAL_1(gateways_gateway_47__EVAL_1),
    ._EVAL_2(gateways_gateway_47__EVAL_2),
    ._EVAL_3(gateways_gateway_47__EVAL_3),
    ._EVAL_4(gateways_gateway_47__EVAL_4)
  );
  _EVAL_96 gateways_gateway_54 (
    ._EVAL(gateways_gateway_54__EVAL),
    ._EVAL_0(gateways_gateway_54__EVAL_0),
    ._EVAL_1(gateways_gateway_54__EVAL_1),
    ._EVAL_2(gateways_gateway_54__EVAL_2),
    ._EVAL_3(gateways_gateway_54__EVAL_3),
    ._EVAL_4(gateways_gateway_54__EVAL_4)
  );
  _EVAL_96 gateways_gateway_118 (
    ._EVAL(gateways_gateway_118__EVAL),
    ._EVAL_0(gateways_gateway_118__EVAL_0),
    ._EVAL_1(gateways_gateway_118__EVAL_1),
    ._EVAL_2(gateways_gateway_118__EVAL_2),
    ._EVAL_3(gateways_gateway_118__EVAL_3),
    ._EVAL_4(gateways_gateway_118__EVAL_4)
  );
  _EVAL_96 gateways_gateway_120 (
    ._EVAL(gateways_gateway_120__EVAL),
    ._EVAL_0(gateways_gateway_120__EVAL_0),
    ._EVAL_1(gateways_gateway_120__EVAL_1),
    ._EVAL_2(gateways_gateway_120__EVAL_2),
    ._EVAL_3(gateways_gateway_120__EVAL_3),
    ._EVAL_4(gateways_gateway_120__EVAL_4)
  );
  _EVAL_96 gateways_gateway_99 (
    ._EVAL(gateways_gateway_99__EVAL),
    ._EVAL_0(gateways_gateway_99__EVAL_0),
    ._EVAL_1(gateways_gateway_99__EVAL_1),
    ._EVAL_2(gateways_gateway_99__EVAL_2),
    ._EVAL_3(gateways_gateway_99__EVAL_3),
    ._EVAL_4(gateways_gateway_99__EVAL_4)
  );
  _EVAL_96 gateways_gateway_75 (
    ._EVAL(gateways_gateway_75__EVAL),
    ._EVAL_0(gateways_gateway_75__EVAL_0),
    ._EVAL_1(gateways_gateway_75__EVAL_1),
    ._EVAL_2(gateways_gateway_75__EVAL_2),
    ._EVAL_3(gateways_gateway_75__EVAL_3),
    ._EVAL_4(gateways_gateway_75__EVAL_4)
  );
  _EVAL_96 gateways_gateway_73 (
    ._EVAL(gateways_gateway_73__EVAL),
    ._EVAL_0(gateways_gateway_73__EVAL_0),
    ._EVAL_1(gateways_gateway_73__EVAL_1),
    ._EVAL_2(gateways_gateway_73__EVAL_2),
    ._EVAL_3(gateways_gateway_73__EVAL_3),
    ._EVAL_4(gateways_gateway_73__EVAL_4)
  );
  _EVAL_96 gateways_gateway_53 (
    ._EVAL(gateways_gateway_53__EVAL),
    ._EVAL_0(gateways_gateway_53__EVAL_0),
    ._EVAL_1(gateways_gateway_53__EVAL_1),
    ._EVAL_2(gateways_gateway_53__EVAL_2),
    ._EVAL_3(gateways_gateway_53__EVAL_3),
    ._EVAL_4(gateways_gateway_53__EVAL_4)
  );
  _EVAL_96 gateways_gateway_23 (
    ._EVAL(gateways_gateway_23__EVAL),
    ._EVAL_0(gateways_gateway_23__EVAL_0),
    ._EVAL_1(gateways_gateway_23__EVAL_1),
    ._EVAL_2(gateways_gateway_23__EVAL_2),
    ._EVAL_3(gateways_gateway_23__EVAL_3),
    ._EVAL_4(gateways_gateway_23__EVAL_4)
  );
  _EVAL_96 gateways_gateway_100 (
    ._EVAL(gateways_gateway_100__EVAL),
    ._EVAL_0(gateways_gateway_100__EVAL_0),
    ._EVAL_1(gateways_gateway_100__EVAL_1),
    ._EVAL_2(gateways_gateway_100__EVAL_2),
    ._EVAL_3(gateways_gateway_100__EVAL_3),
    ._EVAL_4(gateways_gateway_100__EVAL_4)
  );
  _EVAL_96 gateways_gateway_126 (
    ._EVAL(gateways_gateway_126__EVAL),
    ._EVAL_0(gateways_gateway_126__EVAL_0),
    ._EVAL_1(gateways_gateway_126__EVAL_1),
    ._EVAL_2(gateways_gateway_126__EVAL_2),
    ._EVAL_3(gateways_gateway_126__EVAL_3),
    ._EVAL_4(gateways_gateway_126__EVAL_4)
  );
  _EVAL_96 gateways_gateway_117 (
    ._EVAL(gateways_gateway_117__EVAL),
    ._EVAL_0(gateways_gateway_117__EVAL_0),
    ._EVAL_1(gateways_gateway_117__EVAL_1),
    ._EVAL_2(gateways_gateway_117__EVAL_2),
    ._EVAL_3(gateways_gateway_117__EVAL_3),
    ._EVAL_4(gateways_gateway_117__EVAL_4)
  );
  _EVAL_96 gateways_gateway_63 (
    ._EVAL(gateways_gateway_63__EVAL),
    ._EVAL_0(gateways_gateway_63__EVAL_0),
    ._EVAL_1(gateways_gateway_63__EVAL_1),
    ._EVAL_2(gateways_gateway_63__EVAL_2),
    ._EVAL_3(gateways_gateway_63__EVAL_3),
    ._EVAL_4(gateways_gateway_63__EVAL_4)
  );
  _EVAL_97 fanin (
    ._EVAL(fanin__EVAL),
    ._EVAL_0(fanin__EVAL_0),
    ._EVAL_1(fanin__EVAL_1),
    ._EVAL_2(fanin__EVAL_2),
    ._EVAL_3(fanin__EVAL_3),
    ._EVAL_4(fanin__EVAL_4),
    ._EVAL_5(fanin__EVAL_5),
    ._EVAL_6(fanin__EVAL_6),
    ._EVAL_7(fanin__EVAL_7),
    ._EVAL_8(fanin__EVAL_8),
    ._EVAL_9(fanin__EVAL_9),
    ._EVAL_10(fanin__EVAL_10),
    ._EVAL_11(fanin__EVAL_11),
    ._EVAL_12(fanin__EVAL_12),
    ._EVAL_13(fanin__EVAL_13),
    ._EVAL_14(fanin__EVAL_14),
    ._EVAL_15(fanin__EVAL_15),
    ._EVAL_16(fanin__EVAL_16),
    ._EVAL_17(fanin__EVAL_17),
    ._EVAL_18(fanin__EVAL_18),
    ._EVAL_19(fanin__EVAL_19),
    ._EVAL_20(fanin__EVAL_20),
    ._EVAL_21(fanin__EVAL_21),
    ._EVAL_22(fanin__EVAL_22),
    ._EVAL_23(fanin__EVAL_23),
    ._EVAL_24(fanin__EVAL_24),
    ._EVAL_25(fanin__EVAL_25),
    ._EVAL_26(fanin__EVAL_26),
    ._EVAL_27(fanin__EVAL_27),
    ._EVAL_28(fanin__EVAL_28),
    ._EVAL_29(fanin__EVAL_29),
    ._EVAL_30(fanin__EVAL_30),
    ._EVAL_31(fanin__EVAL_31),
    ._EVAL_32(fanin__EVAL_32),
    ._EVAL_33(fanin__EVAL_33),
    ._EVAL_34(fanin__EVAL_34),
    ._EVAL_35(fanin__EVAL_35),
    ._EVAL_36(fanin__EVAL_36),
    ._EVAL_37(fanin__EVAL_37),
    ._EVAL_38(fanin__EVAL_38),
    ._EVAL_39(fanin__EVAL_39),
    ._EVAL_40(fanin__EVAL_40),
    ._EVAL_41(fanin__EVAL_41),
    ._EVAL_42(fanin__EVAL_42),
    ._EVAL_43(fanin__EVAL_43),
    ._EVAL_44(fanin__EVAL_44),
    ._EVAL_45(fanin__EVAL_45),
    ._EVAL_46(fanin__EVAL_46),
    ._EVAL_47(fanin__EVAL_47),
    ._EVAL_48(fanin__EVAL_48),
    ._EVAL_49(fanin__EVAL_49),
    ._EVAL_50(fanin__EVAL_50),
    ._EVAL_51(fanin__EVAL_51),
    ._EVAL_52(fanin__EVAL_52),
    ._EVAL_53(fanin__EVAL_53),
    ._EVAL_54(fanin__EVAL_54),
    ._EVAL_55(fanin__EVAL_55),
    ._EVAL_56(fanin__EVAL_56),
    ._EVAL_57(fanin__EVAL_57),
    ._EVAL_58(fanin__EVAL_58),
    ._EVAL_59(fanin__EVAL_59),
    ._EVAL_60(fanin__EVAL_60),
    ._EVAL_61(fanin__EVAL_61),
    ._EVAL_62(fanin__EVAL_62),
    ._EVAL_63(fanin__EVAL_63),
    ._EVAL_64(fanin__EVAL_64),
    ._EVAL_65(fanin__EVAL_65),
    ._EVAL_66(fanin__EVAL_66),
    ._EVAL_67(fanin__EVAL_67),
    ._EVAL_68(fanin__EVAL_68),
    ._EVAL_69(fanin__EVAL_69),
    ._EVAL_70(fanin__EVAL_70),
    ._EVAL_71(fanin__EVAL_71),
    ._EVAL_72(fanin__EVAL_72),
    ._EVAL_73(fanin__EVAL_73),
    ._EVAL_74(fanin__EVAL_74),
    ._EVAL_75(fanin__EVAL_75),
    ._EVAL_76(fanin__EVAL_76),
    ._EVAL_77(fanin__EVAL_77),
    ._EVAL_78(fanin__EVAL_78),
    ._EVAL_79(fanin__EVAL_79),
    ._EVAL_80(fanin__EVAL_80),
    ._EVAL_81(fanin__EVAL_81),
    ._EVAL_82(fanin__EVAL_82),
    ._EVAL_83(fanin__EVAL_83),
    ._EVAL_84(fanin__EVAL_84),
    ._EVAL_85(fanin__EVAL_85),
    ._EVAL_86(fanin__EVAL_86),
    ._EVAL_87(fanin__EVAL_87),
    ._EVAL_88(fanin__EVAL_88),
    ._EVAL_89(fanin__EVAL_89),
    ._EVAL_90(fanin__EVAL_90),
    ._EVAL_91(fanin__EVAL_91),
    ._EVAL_92(fanin__EVAL_92),
    ._EVAL_93(fanin__EVAL_93),
    ._EVAL_94(fanin__EVAL_94),
    ._EVAL_95(fanin__EVAL_95),
    ._EVAL_96(fanin__EVAL_96),
    ._EVAL_97(fanin__EVAL_97),
    ._EVAL_98(fanin__EVAL_98),
    ._EVAL_99(fanin__EVAL_99),
    ._EVAL_100(fanin__EVAL_100),
    ._EVAL_101(fanin__EVAL_101),
    ._EVAL_102(fanin__EVAL_102),
    ._EVAL_103(fanin__EVAL_103),
    ._EVAL_104(fanin__EVAL_104),
    ._EVAL_105(fanin__EVAL_105),
    ._EVAL_106(fanin__EVAL_106),
    ._EVAL_107(fanin__EVAL_107),
    ._EVAL_108(fanin__EVAL_108),
    ._EVAL_109(fanin__EVAL_109),
    ._EVAL_110(fanin__EVAL_110),
    ._EVAL_111(fanin__EVAL_111),
    ._EVAL_112(fanin__EVAL_112),
    ._EVAL_113(fanin__EVAL_113),
    ._EVAL_114(fanin__EVAL_114),
    ._EVAL_115(fanin__EVAL_115),
    ._EVAL_116(fanin__EVAL_116),
    ._EVAL_117(fanin__EVAL_117),
    ._EVAL_118(fanin__EVAL_118),
    ._EVAL_119(fanin__EVAL_119),
    ._EVAL_120(fanin__EVAL_120),
    ._EVAL_121(fanin__EVAL_121),
    ._EVAL_122(fanin__EVAL_122),
    ._EVAL_123(fanin__EVAL_123),
    ._EVAL_124(fanin__EVAL_124),
    ._EVAL_125(fanin__EVAL_125),
    ._EVAL_126(fanin__EVAL_126),
    ._EVAL_127(fanin__EVAL_127),
    ._EVAL_128(fanin__EVAL_128)
  );
  _EVAL_96 gateways_gateway_29 (
    ._EVAL(gateways_gateway_29__EVAL),
    ._EVAL_0(gateways_gateway_29__EVAL_0),
    ._EVAL_1(gateways_gateway_29__EVAL_1),
    ._EVAL_2(gateways_gateway_29__EVAL_2),
    ._EVAL_3(gateways_gateway_29__EVAL_3),
    ._EVAL_4(gateways_gateway_29__EVAL_4)
  );
  _EVAL_96 gateways_gateway_79 (
    ._EVAL(gateways_gateway_79__EVAL),
    ._EVAL_0(gateways_gateway_79__EVAL_0),
    ._EVAL_1(gateways_gateway_79__EVAL_1),
    ._EVAL_2(gateways_gateway_79__EVAL_2),
    ._EVAL_3(gateways_gateway_79__EVAL_3),
    ._EVAL_4(gateways_gateway_79__EVAL_4)
  );
  _EVAL_96 gateways_gateway_106 (
    ._EVAL(gateways_gateway_106__EVAL),
    ._EVAL_0(gateways_gateway_106__EVAL_0),
    ._EVAL_1(gateways_gateway_106__EVAL_1),
    ._EVAL_2(gateways_gateway_106__EVAL_2),
    ._EVAL_3(gateways_gateway_106__EVAL_3),
    ._EVAL_4(gateways_gateway_106__EVAL_4)
  );
  _EVAL_96 gateways_gateway_121 (
    ._EVAL(gateways_gateway_121__EVAL),
    ._EVAL_0(gateways_gateway_121__EVAL_0),
    ._EVAL_1(gateways_gateway_121__EVAL_1),
    ._EVAL_2(gateways_gateway_121__EVAL_2),
    ._EVAL_3(gateways_gateway_121__EVAL_3),
    ._EVAL_4(gateways_gateway_121__EVAL_4)
  );
  _EVAL_96 gateways_gateway_35 (
    ._EVAL(gateways_gateway_35__EVAL),
    ._EVAL_0(gateways_gateway_35__EVAL_0),
    ._EVAL_1(gateways_gateway_35__EVAL_1),
    ._EVAL_2(gateways_gateway_35__EVAL_2),
    ._EVAL_3(gateways_gateway_35__EVAL_3),
    ._EVAL_4(gateways_gateway_35__EVAL_4)
  );
  _EVAL_96 gateways_gateway_74 (
    ._EVAL(gateways_gateway_74__EVAL),
    ._EVAL_0(gateways_gateway_74__EVAL_0),
    ._EVAL_1(gateways_gateway_74__EVAL_1),
    ._EVAL_2(gateways_gateway_74__EVAL_2),
    ._EVAL_3(gateways_gateway_74__EVAL_3),
    ._EVAL_4(gateways_gateway_74__EVAL_4)
  );
  _EVAL_96 gateways_gateway_66 (
    ._EVAL(gateways_gateway_66__EVAL),
    ._EVAL_0(gateways_gateway_66__EVAL_0),
    ._EVAL_1(gateways_gateway_66__EVAL_1),
    ._EVAL_2(gateways_gateway_66__EVAL_2),
    ._EVAL_3(gateways_gateway_66__EVAL_3),
    ._EVAL_4(gateways_gateway_66__EVAL_4)
  );
  _EVAL_96 gateways_gateway_56 (
    ._EVAL(gateways_gateway_56__EVAL),
    ._EVAL_0(gateways_gateway_56__EVAL_0),
    ._EVAL_1(gateways_gateway_56__EVAL_1),
    ._EVAL_2(gateways_gateway_56__EVAL_2),
    ._EVAL_3(gateways_gateway_56__EVAL_3),
    ._EVAL_4(gateways_gateway_56__EVAL_4)
  );
  _EVAL_96 gateways_gateway_107 (
    ._EVAL(gateways_gateway_107__EVAL),
    ._EVAL_0(gateways_gateway_107__EVAL_0),
    ._EVAL_1(gateways_gateway_107__EVAL_1),
    ._EVAL_2(gateways_gateway_107__EVAL_2),
    ._EVAL_3(gateways_gateway_107__EVAL_3),
    ._EVAL_4(gateways_gateway_107__EVAL_4)
  );
  _EVAL_96 gateways_gateway_8 (
    ._EVAL(gateways_gateway_8__EVAL),
    ._EVAL_0(gateways_gateway_8__EVAL_0),
    ._EVAL_1(gateways_gateway_8__EVAL_1),
    ._EVAL_2(gateways_gateway_8__EVAL_2),
    ._EVAL_3(gateways_gateway_8__EVAL_3),
    ._EVAL_4(gateways_gateway_8__EVAL_4)
  );
  _EVAL_96 gateways_gateway_11 (
    ._EVAL(gateways_gateway_11__EVAL),
    ._EVAL_0(gateways_gateway_11__EVAL_0),
    ._EVAL_1(gateways_gateway_11__EVAL_1),
    ._EVAL_2(gateways_gateway_11__EVAL_2),
    ._EVAL_3(gateways_gateway_11__EVAL_3),
    ._EVAL_4(gateways_gateway_11__EVAL_4)
  );
  _EVAL_96 gateways_gateway_12 (
    ._EVAL(gateways_gateway_12__EVAL),
    ._EVAL_0(gateways_gateway_12__EVAL_0),
    ._EVAL_1(gateways_gateway_12__EVAL_1),
    ._EVAL_2(gateways_gateway_12__EVAL_2),
    ._EVAL_3(gateways_gateway_12__EVAL_3),
    ._EVAL_4(gateways_gateway_12__EVAL_4)
  );
  _EVAL_96 gateways_gateway_57 (
    ._EVAL(gateways_gateway_57__EVAL),
    ._EVAL_0(gateways_gateway_57__EVAL_0),
    ._EVAL_1(gateways_gateway_57__EVAL_1),
    ._EVAL_2(gateways_gateway_57__EVAL_2),
    ._EVAL_3(gateways_gateway_57__EVAL_3),
    ._EVAL_4(gateways_gateway_57__EVAL_4)
  );
  _EVAL_96 gateways_gateway_43 (
    ._EVAL(gateways_gateway_43__EVAL),
    ._EVAL_0(gateways_gateway_43__EVAL_0),
    ._EVAL_1(gateways_gateway_43__EVAL_1),
    ._EVAL_2(gateways_gateway_43__EVAL_2),
    ._EVAL_3(gateways_gateway_43__EVAL_3),
    ._EVAL_4(gateways_gateway_43__EVAL_4)
  );
  _EVAL_96 gateways_gateway_4 (
    ._EVAL(gateways_gateway_4__EVAL),
    ._EVAL_0(gateways_gateway_4__EVAL_0),
    ._EVAL_1(gateways_gateway_4__EVAL_1),
    ._EVAL_2(gateways_gateway_4__EVAL_2),
    ._EVAL_3(gateways_gateway_4__EVAL_3),
    ._EVAL_4(gateways_gateway_4__EVAL_4)
  );
  _EVAL_96 gateways_gateway_36 (
    ._EVAL(gateways_gateway_36__EVAL),
    ._EVAL_0(gateways_gateway_36__EVAL_0),
    ._EVAL_1(gateways_gateway_36__EVAL_1),
    ._EVAL_2(gateways_gateway_36__EVAL_2),
    ._EVAL_3(gateways_gateway_36__EVAL_3),
    ._EVAL_4(gateways_gateway_36__EVAL_4)
  );
  _EVAL_96 gateways_gateway_5 (
    ._EVAL(gateways_gateway_5__EVAL),
    ._EVAL_0(gateways_gateway_5__EVAL_0),
    ._EVAL_1(gateways_gateway_5__EVAL_1),
    ._EVAL_2(gateways_gateway_5__EVAL_2),
    ._EVAL_3(gateways_gateway_5__EVAL_3),
    ._EVAL_4(gateways_gateway_5__EVAL_4)
  );
  _EVAL_96 gateways_gateway_18 (
    ._EVAL(gateways_gateway_18__EVAL),
    ._EVAL_0(gateways_gateway_18__EVAL_0),
    ._EVAL_1(gateways_gateway_18__EVAL_1),
    ._EVAL_2(gateways_gateway_18__EVAL_2),
    ._EVAL_3(gateways_gateway_18__EVAL_3),
    ._EVAL_4(gateways_gateway_18__EVAL_4)
  );
  _EVAL_96 gateways_gateway_50 (
    ._EVAL(gateways_gateway_50__EVAL),
    ._EVAL_0(gateways_gateway_50__EVAL_0),
    ._EVAL_1(gateways_gateway_50__EVAL_1),
    ._EVAL_2(gateways_gateway_50__EVAL_2),
    ._EVAL_3(gateways_gateway_50__EVAL_3),
    ._EVAL_4(gateways_gateway_50__EVAL_4)
  );
  _EVAL_96 gateways_gateway_60 (
    ._EVAL(gateways_gateway_60__EVAL),
    ._EVAL_0(gateways_gateway_60__EVAL_0),
    ._EVAL_1(gateways_gateway_60__EVAL_1),
    ._EVAL_2(gateways_gateway_60__EVAL_2),
    ._EVAL_3(gateways_gateway_60__EVAL_3),
    ._EVAL_4(gateways_gateway_60__EVAL_4)
  );
  _EVAL_96 gateways_gateway_95 (
    ._EVAL(gateways_gateway_95__EVAL),
    ._EVAL_0(gateways_gateway_95__EVAL_0),
    ._EVAL_1(gateways_gateway_95__EVAL_1),
    ._EVAL_2(gateways_gateway_95__EVAL_2),
    ._EVAL_3(gateways_gateway_95__EVAL_3),
    ._EVAL_4(gateways_gateway_95__EVAL_4)
  );
  _EVAL_96 gateways_gateway_13 (
    ._EVAL(gateways_gateway_13__EVAL),
    ._EVAL_0(gateways_gateway_13__EVAL_0),
    ._EVAL_1(gateways_gateway_13__EVAL_1),
    ._EVAL_2(gateways_gateway_13__EVAL_2),
    ._EVAL_3(gateways_gateway_13__EVAL_3),
    ._EVAL_4(gateways_gateway_13__EVAL_4)
  );
  _EVAL_96 gateways_gateway_20 (
    ._EVAL(gateways_gateway_20__EVAL),
    ._EVAL_0(gateways_gateway_20__EVAL_0),
    ._EVAL_1(gateways_gateway_20__EVAL_1),
    ._EVAL_2(gateways_gateway_20__EVAL_2),
    ._EVAL_3(gateways_gateway_20__EVAL_3),
    ._EVAL_4(gateways_gateway_20__EVAL_4)
  );
  _EVAL_96 gateways_gateway_25 (
    ._EVAL(gateways_gateway_25__EVAL),
    ._EVAL_0(gateways_gateway_25__EVAL_0),
    ._EVAL_1(gateways_gateway_25__EVAL_1),
    ._EVAL_2(gateways_gateway_25__EVAL_2),
    ._EVAL_3(gateways_gateway_25__EVAL_3),
    ._EVAL_4(gateways_gateway_25__EVAL_4)
  );
  _EVAL_96 gateways_gateway_19 (
    ._EVAL(gateways_gateway_19__EVAL),
    ._EVAL_0(gateways_gateway_19__EVAL_0),
    ._EVAL_1(gateways_gateway_19__EVAL_1),
    ._EVAL_2(gateways_gateway_19__EVAL_2),
    ._EVAL_3(gateways_gateway_19__EVAL_3),
    ._EVAL_4(gateways_gateway_19__EVAL_4)
  );
  _EVAL_96 gateways_gateway_32 (
    ._EVAL(gateways_gateway_32__EVAL),
    ._EVAL_0(gateways_gateway_32__EVAL_0),
    ._EVAL_1(gateways_gateway_32__EVAL_1),
    ._EVAL_2(gateways_gateway_32__EVAL_2),
    ._EVAL_3(gateways_gateway_32__EVAL_3),
    ._EVAL_4(gateways_gateway_32__EVAL_4)
  );
  _EVAL_96 gateways_gateway_67 (
    ._EVAL(gateways_gateway_67__EVAL),
    ._EVAL_0(gateways_gateway_67__EVAL_0),
    ._EVAL_1(gateways_gateway_67__EVAL_1),
    ._EVAL_2(gateways_gateway_67__EVAL_2),
    ._EVAL_3(gateways_gateway_67__EVAL_3),
    ._EVAL_4(gateways_gateway_67__EVAL_4)
  );
  _EVAL_96 gateways_gateway_93 (
    ._EVAL(gateways_gateway_93__EVAL),
    ._EVAL_0(gateways_gateway_93__EVAL_0),
    ._EVAL_1(gateways_gateway_93__EVAL_1),
    ._EVAL_2(gateways_gateway_93__EVAL_2),
    ._EVAL_3(gateways_gateway_93__EVAL_3),
    ._EVAL_4(gateways_gateway_93__EVAL_4)
  );
  _EVAL_96 gateways_gateway_52 (
    ._EVAL(gateways_gateway_52__EVAL),
    ._EVAL_0(gateways_gateway_52__EVAL_0),
    ._EVAL_1(gateways_gateway_52__EVAL_1),
    ._EVAL_2(gateways_gateway_52__EVAL_2),
    ._EVAL_3(gateways_gateway_52__EVAL_3),
    ._EVAL_4(gateways_gateway_52__EVAL_4)
  );
  _EVAL_96 gateways_gateway_109 (
    ._EVAL(gateways_gateway_109__EVAL),
    ._EVAL_0(gateways_gateway_109__EVAL_0),
    ._EVAL_1(gateways_gateway_109__EVAL_1),
    ._EVAL_2(gateways_gateway_109__EVAL_2),
    ._EVAL_3(gateways_gateway_109__EVAL_3),
    ._EVAL_4(gateways_gateway_109__EVAL_4)
  );
  _EVAL_96 gateways_gateway_64 (
    ._EVAL(gateways_gateway_64__EVAL),
    ._EVAL_0(gateways_gateway_64__EVAL_0),
    ._EVAL_1(gateways_gateway_64__EVAL_1),
    ._EVAL_2(gateways_gateway_64__EVAL_2),
    ._EVAL_3(gateways_gateway_64__EVAL_3),
    ._EVAL_4(gateways_gateway_64__EVAL_4)
  );
  _EVAL_96 gateways_gateway_80 (
    ._EVAL(gateways_gateway_80__EVAL),
    ._EVAL_0(gateways_gateway_80__EVAL_0),
    ._EVAL_1(gateways_gateway_80__EVAL_1),
    ._EVAL_2(gateways_gateway_80__EVAL_2),
    ._EVAL_3(gateways_gateway_80__EVAL_3),
    ._EVAL_4(gateways_gateway_80__EVAL_4)
  );
  _EVAL_96 gateways_gateway_85 (
    ._EVAL(gateways_gateway_85__EVAL),
    ._EVAL_0(gateways_gateway_85__EVAL_0),
    ._EVAL_1(gateways_gateway_85__EVAL_1),
    ._EVAL_2(gateways_gateway_85__EVAL_2),
    ._EVAL_3(gateways_gateway_85__EVAL_3),
    ._EVAL_4(gateways_gateway_85__EVAL_4)
  );
  _EVAL_96 gateways_gateway_48 (
    ._EVAL(gateways_gateway_48__EVAL),
    ._EVAL_0(gateways_gateway_48__EVAL_0),
    ._EVAL_1(gateways_gateway_48__EVAL_1),
    ._EVAL_2(gateways_gateway_48__EVAL_2),
    ._EVAL_3(gateways_gateway_48__EVAL_3),
    ._EVAL_4(gateways_gateway_48__EVAL_4)
  );
  _EVAL_96 gateways_gateway_26 (
    ._EVAL(gateways_gateway_26__EVAL),
    ._EVAL_0(gateways_gateway_26__EVAL_0),
    ._EVAL_1(gateways_gateway_26__EVAL_1),
    ._EVAL_2(gateways_gateway_26__EVAL_2),
    ._EVAL_3(gateways_gateway_26__EVAL_3),
    ._EVAL_4(gateways_gateway_26__EVAL_4)
  );
  _EVAL_96 gateways_gateway_65 (
    ._EVAL(gateways_gateway_65__EVAL),
    ._EVAL_0(gateways_gateway_65__EVAL_0),
    ._EVAL_1(gateways_gateway_65__EVAL_1),
    ._EVAL_2(gateways_gateway_65__EVAL_2),
    ._EVAL_3(gateways_gateway_65__EVAL_3),
    ._EVAL_4(gateways_gateway_65__EVAL_4)
  );
  _EVAL_96 gateways_gateway_62 (
    ._EVAL(gateways_gateway_62__EVAL),
    ._EVAL_0(gateways_gateway_62__EVAL_0),
    ._EVAL_1(gateways_gateway_62__EVAL_1),
    ._EVAL_2(gateways_gateway_62__EVAL_2),
    ._EVAL_3(gateways_gateway_62__EVAL_3),
    ._EVAL_4(gateways_gateway_62__EVAL_4)
  );
  assign fanin__EVAL_19 = _EVAL_355;
  assign _EVAL_2694 = {_EVAL_3242,_EVAL_1673,_EVAL_1944,_EVAL_2944,_EVAL_2268,_EVAL_902,_EVAL_3770,_EVAL_1576,_EVAL_3222
    };
  assign fanin__EVAL_68 = _EVAL_779;
  assign _EVAL_3847 = _EVAL_1193 ? _EVAL_826 : _EVAL_2061;
  assign _EVAL_1178 = out_back__EVAL_3[11];
  assign fanin__EVAL_29 = _EVAL_966;
  assign _EVAL_715 = _EVAL_1976 & _EVAL_2035;
  assign _EVAL_784 = _EVAL_3108 & _EVAL_826;
  assign _EVAL_2476 = _EVAL_1171 ? _EVAL_826 : _EVAL_2354;
  assign gateways_gateway_110__EVAL_2 = _EVAL_2917[111];
  assign _EVAL_2651 = _EVAL_203 & _EVAL_2035;
  assign _EVAL_383 = _EVAL_2686 | gateways_gateway_27__EVAL_4;
  assign gateways_gateway_105__EVAL_3 = _EVAL_110;
  assign _EVAL_2080 = 10'h72 == _EVAL_2998;
  assign _EVAL_3442 = _EVAL_647 ? {{29'd0}, _EVAL_1358} : _EVAL_2918;
  assign _EVAL_2142 = _EVAL_1325 & _EVAL_2035;
  assign gateways_gateway_21__EVAL_2 = _EVAL_2917[22];
  assign _EVAL_3485 = ~_EVAL_3174;
  assign _EVAL_386 = {_EVAL_1507,_EVAL_2297,_EVAL_2221,_EVAL_3199,_EVAL_1524,_EVAL_2153,_EVAL_2900,_EVAL_744,_EVAL_2682,
    _EVAL_3644};
  assign gateways_gateway_93__EVAL_3 = _EVAL_110;
  assign gateways_gateway_23__EVAL_1 = ~_EVAL_3129;
  assign _EVAL_1301 = _EVAL_910 & _EVAL_2035;
  assign gateways_gateway_74__EVAL_0 = _EVAL_9;
  assign gateways_gateway_73__EVAL_0 = _EVAL_9;
  assign _EVAL_1274 = 10'h1f == _EVAL_2998;
  assign _EVAL_1133 = _EVAL_1809 ? _EVAL_826 : _EVAL_975;
  assign gateways_gateway_56__EVAL = _EVAL_26;
  assign gateways_gateway_6__EVAL_2 = _EVAL_2917[7];
  assign _EVAL_1428 = _EVAL_3349[67];
  assign _EVAL_3587 = _EVAL_195 & _EVAL_1793;
  assign gateways_gateway_72__EVAL_1 = ~_EVAL_2719;
  assign _EVAL_1510 = ~_EVAL_2077;
  assign gateways_gateway_72__EVAL_0 = _EVAL_9;
  assign _EVAL_3416 = _EVAL_3367 ? _EVAL_826 : _EVAL_631;
  assign _EVAL_607 = _EVAL_2216 | gateways_gateway_54__EVAL_4;
  assign _EVAL_937 = ~_EVAL_3271;
  assign _EVAL_913 = _EVAL_195 & _EVAL_369;
  assign _EVAL_973 = ~_EVAL_1541;
  assign gateways_gateway_87__EVAL_3 = _EVAL_110;
  assign _EVAL_2534 = _EVAL_1998 & _EVAL_826;
  assign _EVAL_1036 = _EVAL_573 ? _EVAL_2979 : _EVAL_1130;
  assign gateways_gateway_58__EVAL_3 = _EVAL_110;
  assign gateways_gateway_14__EVAL_3 = _EVAL_110;
  assign gateways_gateway_17__EVAL_2 = _EVAL_2917[18];
  assign _EVAL_1754 = _EVAL_904 | gateways_gateway_112__EVAL_4;
  assign _EVAL_3450 = _EVAL_1902 ? _EVAL_826 : _EVAL_2131;
  assign gateways_gateway_25__EVAL_1 = ~_EVAL_3268;
  assign fanin__EVAL_31 = _EVAL_2921;
  assign gateways_gateway_46__EVAL_2 = _EVAL_2917[47];
  assign gateways_gateway_74__EVAL = _EVAL_31;
  assign fanin__EVAL_106 = _EVAL_3590;
  assign _EVAL_3408 = _EVAL_3030 & _EVAL_2957;
  assign _EVAL_2910 = _EVAL_285 | gateways_gateway_24__EVAL_4;
  assign _EVAL_2966 = ~_EVAL_3523;
  assign _EVAL_1946 = _EVAL_195 & _EVAL_3099;
  assign gateways_gateway_21__EVAL_1 = ~_EVAL_302;
  assign _EVAL_288 = _EVAL_2517 & _EVAL_2035;
  assign _EVAL_2494 = _EVAL_3030 & _EVAL_3266;
  assign _EVAL_1364 = _EVAL_2415 | gateways_gateway_88__EVAL_4;
  assign _EVAL_1833 = _EVAL_964 | gateways_gateway_41__EVAL_4;
  assign _EVAL_97 = _EVAL_3416 ? _EVAL_1299 : 32'h0;
  assign gateways_gateway_91__EVAL_2 = _EVAL_2917[92];
  assign gateways_gateway_7__EVAL_1 = ~_EVAL_780;
  assign _EVAL_3719 = _EVAL_667 & _EVAL_2035;
  assign _EVAL_1592 = _EVAL_195 & _EVAL_640;
  assign _EVAL_1072 = _EVAL_195 & _EVAL_2814;
  assign gateways_gateway_117__EVAL_2 = _EVAL_2917[118];
  assign gateways_gateway_99__EVAL_1 = ~_EVAL_3656;
  assign gateways_gateway_75__EVAL_1 = ~_EVAL_2900;
  assign _EVAL_979 = _EVAL_3599 | gateways_gateway_115__EVAL_4;
  assign gateways_gateway_27__EVAL_0 = _EVAL_9;
  assign _EVAL_2354 = _EVAL_499 ? _EVAL_826 : _EVAL_2929;
  assign _EVAL_873 = _EVAL_2671 & _EVAL_826;
  assign _EVAL_3061 = ~_EVAL_842;
  assign gateways_gateway_33__EVAL_0 = _EVAL_9;
  assign _EVAL_1973 = _EVAL_651[127];
  assign _EVAL_1738 = _EVAL_1237 & _EVAL_826;
  assign _EVAL_3378 = _EVAL_3349[82];
  assign _EVAL_3251 = 10'h44 == _EVAL_2998;
  assign _EVAL_3742 = _EVAL_3311 | gateways_gateway_103__EVAL_4;
  assign gateways_gateway_71__EVAL_0 = _EVAL_9;
  assign _EVAL_2410 = _EVAL_2728 & _EVAL_2035;
  assign _EVAL_2275 = _EVAL_2844 ? {{29'd0}, _EVAL_1843} : _EVAL_569;
  assign fanin__EVAL_77 = _EVAL_2981;
  assign _EVAL_1587 = _EVAL_3684 ? 8'hff : 8'h0;
  assign _EVAL_2308 = 10'ha == _EVAL_2998;
  assign _EVAL_381 = _EVAL_195 & _EVAL_2346;
  assign _EVAL_3642 = ~_EVAL_1180;
  assign _EVAL_1211 = _EVAL_195 & _EVAL_2798;
  assign _EVAL_1972 = _EVAL_3152 & _EVAL_2035;
  assign _EVAL_3034 = _EVAL_1923 ? _EVAL_826 : _EVAL_2759;
  assign _EVAL_3756 = _EVAL_1884 ? _EVAL_826 : _EVAL_752;
  assign _EVAL_2049 = _EVAL_2080 ? _EVAL_826 : _EVAL_1645;
  assign fanin__EVAL_117 = _EVAL_3513;
  assign gateways_gateway_55__EVAL_1 = ~_EVAL_2502;
  assign _EVAL_1015 = _EVAL_3341 | gateways_gateway_50__EVAL_4;
  assign gateways_gateway_24__EVAL = _EVAL_80;
  assign _EVAL_2451 = _EVAL_2308 ? {{29'd0}, _EVAL_966} : _EVAL_743;
  assign _EVAL_1707 = _EVAL_195 & _EVAL_1396;
  assign _EVAL_647 = 10'h33 == _EVAL_2998;
  assign _EVAL_1328 = _EVAL_3288 & _EVAL_2035;
  assign _EVAL_2217 = _EVAL_3278 & _EVAL_826;
  assign gateways_gateway_66__EVAL_1 = ~_EVAL_3387;
  assign _EVAL_2453 = _EVAL_2822 | gateways_gateway_30__EVAL_4;
  assign _EVAL_3637 = _EVAL_651[11];
  assign gateways_gateway_85__EVAL_3 = _EVAL_110;
  assign _EVAL_364 = _EVAL_2525 ? _EVAL_826 : _EVAL_2049;
  assign fanin__EVAL_34 = _EVAL_2477;
  assign gateways_gateway_86__EVAL_0 = _EVAL_9;
  assign gateways_gateway_97__EVAL_2 = _EVAL_2917[98];
  assign _EVAL_1899 = _EVAL_3616 & _EVAL_826;
  assign _EVAL_2846 = _EVAL_583 & _EVAL_2035;
  assign _EVAL_3206 = _EVAL_651[49];
  assign _EVAL_366 = _EVAL_164 ? {{29'd0}, _EVAL_3590} : _EVAL_1009;
  assign gateways_gateway_34__EVAL_2 = _EVAL_2917[35];
  assign _EVAL_3374 = _EVAL_195 & _EVAL_1532;
  assign _EVAL_238 = _EVAL_195 & _EVAL_1057;
  assign fanin__EVAL_88 = _EVAL_707;
  assign gateways_gateway__EVAL_0 = _EVAL_9;
  assign _EVAL_3122 = _EVAL_3349[107];
  assign _EVAL_2838 = _EVAL_404 ? {{29'd0}, _EVAL_1099} : _EVAL_1568;
  assign gateways_gateway_48__EVAL_0 = _EVAL_9;
  assign _EVAL_2385 = _EVAL_1918 ? {{29'd0}, _EVAL_355} : _EVAL_2628;
  assign _EVAL_2934 = _EVAL_1918 ? _EVAL_826 : _EVAL_241;
  assign _EVAL_1222 = ~_EVAL_1751;
  assign gateways_gateway_68__EVAL = _EVAL_98;
  assign _EVAL_3410 = _EVAL_2534 & _EVAL_2035;
  assign _EVAL_1854 = _EVAL_2985 ? {{29'd0}, _EVAL_1771} : _EVAL_1997;
  assign _EVAL_691 = _EVAL_648 & _EVAL_826;
  assign _EVAL_1061 = ~_EVAL_3393;
  assign _EVAL_1920 = 10'h100 == _EVAL_2998;
  assign _EVAL_3722 = _EVAL_691 & _EVAL_2035;
  assign _EVAL_2075 = _EVAL_2347 ? _EVAL_826 : _EVAL_1133;
  assign gateways_gateway_60__EVAL_2 = _EVAL_2917[61];
  assign gateways_gateway_15__EVAL_1 = ~_EVAL_911;
  assign gateways_gateway_55__EVAL_3 = _EVAL_110;
  assign fanin__EVAL_85 = _EVAL_1692;
  assign _EVAL_3433 = _EVAL_195 & _EVAL_3368;
  assign _EVAL_3286 = _EVAL_2313 & _EVAL_2035;
  assign gateways_gateway_124__EVAL_2 = _EVAL_2917[125];
  assign _EVAL_390 = ~_EVAL_3246;
  assign gateways_gateway_60__EVAL_3 = _EVAL_110;
  assign gateways_gateway_63__EVAL_1 = ~_EVAL_526;
  assign _EVAL_1443 = _EVAL_3476 ? _EVAL_826 : _EVAL_2094;
  assign gateways_gateway_99__EVAL_0 = _EVAL_9;
  assign _EVAL_1466 = _EVAL_3349[50];
  assign _EVAL_755 = ~_EVAL_3171;
  assign gateways_gateway_13__EVAL_3 = _EVAL_110;
  assign _EVAL_485 = _EVAL_2712 & _EVAL_2035;
  assign _EVAL_1447 = ~_EVAL_2904;
  assign _EVAL_1167 = _EVAL_3221 ? {{29'd0}, _EVAL_2030} : _EVAL_1374;
  assign gateways_gateway_63__EVAL = _EVAL_113;
  assign _EVAL_323 = _EVAL_195 & _EVAL_2234;
  assign _EVAL_817 = _EVAL_651[74];
  assign _EVAL_2623 = _EVAL_651[41];
  assign _EVAL_1949 = _EVAL_3349[14];
  assign _EVAL_3220 = _EVAL_195 & _EVAL_2103;
  assign _EVAL_3418 = _EVAL_2021 ? _EVAL_826 : _EVAL_3528;
  assign gateways_gateway_126__EVAL_3 = _EVAL_110;
  assign _EVAL_1184 = _EVAL_3349[81];
  assign gateways_gateway_69__EVAL_3 = _EVAL_110;
  assign gateways_gateway_75__EVAL_0 = _EVAL_9;
  assign _EVAL_1723 = _EVAL_165 ? 8'hff : 8'h0;
  assign _EVAL_190 = _EVAL_1666 ? _EVAL_175 : _EVAL_1659;
  assign _EVAL_1855 = ~_EVAL_2812;
  assign out_back__EVAL_14 = _EVAL_17;
  assign gateways_gateway_35__EVAL_3 = _EVAL_110;
  assign gateways_gateway_116__EVAL = _EVAL_90;
  assign _EVAL_2773 = _EVAL_3600 & _EVAL_2035;
  assign _EVAL_1645 = _EVAL_2397 ? _EVAL_826 : _EVAL_2659;
  assign gateways_gateway_24__EVAL_1 = ~_EVAL_2370;
  assign _EVAL_3393 = _EVAL_3349[20];
  assign _EVAL_1032 = _EVAL_3434 ? _EVAL_826 : _EVAL_1822;
  assign gateways_gateway_51__EVAL = _EVAL_20;
  assign _EVAL_910 = _EVAL_1072 & _EVAL_826;
  assign _EVAL_1809 = 10'h14 == _EVAL_2998;
  assign gateways_gateway_11__EVAL_0 = _EVAL_9;
  assign _EVAL_1250 = _EVAL_2977 & _EVAL_2035;
  assign gateways_gateway_86__EVAL_1 = ~_EVAL_1127;
  assign _EVAL_3339 = _EVAL_3328 & _EVAL_2957;
  assign _EVAL_3667 = ~out_back__EVAL;
  assign fanin__EVAL_124 = _EVAL_2853;
  assign _EVAL_2929 = _EVAL_1666 ? _EVAL_826 : _EVAL_2053;
  assign _EVAL_3443 = _EVAL_2885 & _EVAL_2035;
  assign _EVAL_2803 = 10'h3a == _EVAL_2998;
  assign _EVAL_688 = ~_EVAL_2366;
  assign _EVAL_2276 = ~_EVAL_1243;
  assign fanin__EVAL_28 = _EVAL_2309;
  assign gateways_gateway_47__EVAL_2 = _EVAL_2917[48];
  assign gateways_gateway_102__EVAL_3 = _EVAL_110;
  assign _EVAL_2879 = _EVAL_651[112];
  assign _EVAL_1544 = _EVAL_651[72];
  assign _EVAL_1339 = _EVAL_2607 | gateways_gateway_90__EVAL_4;
  assign _EVAL_3743 = _EVAL_1435 ? {{29'd0}, _EVAL_2988} : _EVAL_492;
  assign gateways_gateway_49__EVAL_3 = _EVAL_110;
  assign _EVAL_3354 = _EVAL_820 | gateways_gateway_73__EVAL_4;
  assign fanin__EVAL_59 = _EVAL_3290;
  assign _EVAL_906 = _EVAL_2616 & _EVAL_826;
  assign out_back__EVAL_4 = _EVAL_6 == 3'h4;
  assign gateways_gateway_109__EVAL_2 = _EVAL_2917[110];
  assign _EVAL_2957 = &_EVAL_2914;
  assign _EVAL_834 = _EVAL_3545 | gateways_gateway_86__EVAL_4;
  assign _EVAL_2724 = _EVAL_959 ? _EVAL_826 : _EVAL_699;
  assign gateways_gateway_49__EVAL_2 = _EVAL_2917[50];
  assign fanin__EVAL_7 = _EVAL_778;
  assign gateways_gateway_91__EVAL_0 = _EVAL_9;
  assign _EVAL_1441 = _EVAL_166 ? {{29'd0}, _EVAL_3653} : _EVAL_2385;
  assign gateways_gateway_54__EVAL_3 = _EVAL_110;
  assign _EVAL_487 = _EVAL_195 & _EVAL_709;
  assign gateways_gateway_98__EVAL_3 = _EVAL_110;
  assign _EVAL_2199 = _EVAL_2693 ? {{29'd0}, _EVAL_2518} : _EVAL_2226;
  assign _EVAL_775 = _EVAL_3201 ? _EVAL_826 : _EVAL_1631;
  assign _EVAL_1488 = _EVAL_3571 ? _EVAL_826 : _EVAL_2742;
  assign _EVAL_1875 = _EVAL_651[121];
  assign _EVAL_828 = _EVAL_2956 ? _EVAL_826 : _EVAL_954;
  assign _EVAL_1729 = _EVAL_2249 & _EVAL_2035;
  assign _EVAL_3147 = out_back__EVAL_3[4];
  assign _EVAL_3162 = _EVAL_2622 | gateways_gateway_15__EVAL_4;
  assign _EVAL_2561 = 10'h101 == _EVAL_2998;
  assign _EVAL_3725 = _EVAL_195 & _EVAL_1875;
  assign _EVAL_982 = {_EVAL_1638,_EVAL_1928,_EVAL_3059,_EVAL_3242,_EVAL_1673,_EVAL_1944,_EVAL_2944,_EVAL_2268,_EVAL_902,
    _EVAL_576};
  assign gateways_gateway_111__EVAL_3 = _EVAL_110;
  assign _EVAL_3312 = _EVAL_195 & _EVAL_2865;
  assign gateways_gateway_109__EVAL = _EVAL_64;
  assign _EVAL_693 = _EVAL_651[120];
  assign _EVAL_540 = _EVAL_195 & _EVAL_295;
  assign _EVAL_2175 = out_back__EVAL_1;
  assign gateways_gateway_47__EVAL_3 = _EVAL_110;
  assign fanin__EVAL_104 = _EVAL_3516;
  assign gateways_gateway_107__EVAL = _EVAL_108;
  assign _EVAL_1009 = _EVAL_3504 ? {{29'd0}, _EVAL_779} : _EVAL_3084;
  assign _EVAL_1371 = _EVAL_651[256];
  assign _EVAL_1990 = _EVAL_195 & _EVAL_3757;
  assign _EVAL_1282 = 10'h58 == _EVAL_2998;
  assign gateways_gateway_82__EVAL = _EVAL_92;
  assign gateways_gateway_97__EVAL_3 = _EVAL_110;
  assign gateways_gateway_94__EVAL_2 = _EVAL_2917[95];
  assign _EVAL_1023 = _EVAL_2099 | gateways_gateway_96__EVAL_4;
  assign _EVAL_3262 = _EVAL_1433 ? {{29'd0}, _EVAL_2477} : _EVAL_2284;
  assign _EVAL_3557 = _EVAL_3349[119];
  assign _EVAL_3108 = _EVAL_195 & _EVAL_840;
  assign _EVAL_2969 = _EVAL_3236 ? {{29'd0}, _EVAL_3072} : _EVAL_478;
  assign _EVAL_871 = _EVAL_627 & _EVAL_2035;
  assign _EVAL_2329 = _EVAL_2801 & _EVAL_2035;
  assign _EVAL_1935 = _EVAL_869 ? _EVAL_826 : _EVAL_3488;
  assign _EVAL_1942 = _EVAL_651[109];
  assign _EVAL_1903 = ~_EVAL_1828;
  assign _EVAL_3815 = _EVAL_2693 ? _EVAL_826 : _EVAL_1622;
  assign gateways_gateway_65__EVAL_3 = _EVAL_110;
  assign _EVAL_956 = _EVAL_195 & _EVAL_1712;
  assign gateways_gateway_114__EVAL_3 = _EVAL_110;
  assign _EVAL_3017 = _EVAL_2803 ? {{29'd0}, _EVAL_1569} : _EVAL_3370;
  assign _EVAL_164 = 10'h55 == _EVAL_2998;
  assign _EVAL_1892 = _EVAL_195 & _EVAL_3588;
  assign gateways_gateway_110__EVAL_0 = _EVAL_9;
  assign fanin__EVAL_122 = _EVAL_2531;
  assign _EVAL_2980 = _EVAL_195 & _EVAL_3489;
  assign gateways_gateway_50__EVAL_3 = _EVAL_110;
  assign _EVAL_3723 = _EVAL_2274 ? _EVAL_826 : _EVAL_1741;
  assign fanin__EVAL_72 = _EVAL_172;
  assign _EVAL_3064 = _EVAL_3205 & _EVAL_2035;
  assign gateways_gateway_18__EVAL_0 = _EVAL_9;
  assign _EVAL_60 = out_back__EVAL_2;
  assign _EVAL_1610 = _EVAL_195 & _EVAL_2233;
  assign _EVAL_2017 = _EVAL_3349[118];
  assign _EVAL_362 = _EVAL_3349[69];
  assign _EVAL_3152 = _EVAL_314 & _EVAL_826;
  assign gateways_gateway_89__EVAL = _EVAL_79;
  assign fanin__EVAL_110 = _EVAL_628;
  assign _EVAL_1446 = _EVAL_1211 & _EVAL_826;
  assign gateways_gateway_53__EVAL_2 = _EVAL_2917[54];
  assign _EVAL_3217 = _EVAL_195 & _EVAL_3462;
  assign gateways_gateway_61__EVAL_3 = _EVAL_110;
  assign gateways_gateway_95__EVAL_1 = ~_EVAL_415;
  assign fanin__EVAL_80 = _EVAL_1358;
  assign _EVAL_165 = out_back__EVAL_12[1];
  assign _EVAL_957 = _EVAL_446 ? {{29'd0}, _EVAL_3516} : _EVAL_892;
  assign _EVAL_643 = _EVAL_3349[58];
  assign _EVAL_759 = ~_EVAL_2604;
  assign _EVAL_3165 = _EVAL_651[66];
  assign _EVAL_573 = 10'h103 == _EVAL_2998;
  assign _EVAL_639 = ~_EVAL_3704;
  assign _EVAL_3684 = out_back__EVAL_12[3];
  assign _EVAL_751 = _EVAL_195 & _EVAL_3701;
  assign _EVAL_1239 = out_back__EVAL_3[10];
  assign _EVAL_337 = 10'h57 == _EVAL_2998;
  assign _EVAL_3651 = _EVAL_651[44];
  assign _EVAL_2758 = _EVAL_2377 >> _EVAL_1408;
  assign _EVAL_2633 = _EVAL_651[114];
  assign _EVAL_783 = ~_EVAL_1451;
  assign gateways_gateway_40__EVAL_2 = _EVAL_2917[41];
  assign _EVAL_3681 = _EVAL_651[22];
  assign _EVAL_1043 = _EVAL_3349[84];
  assign _EVAL_1698 = _EVAL_1269 | gateways_gateway_8__EVAL_4;
  assign gateways_gateway_122__EVAL_0 = _EVAL_9;
  assign gateways_gateway_13__EVAL = _EVAL_140;
  assign _EVAL_1112 = _EVAL_1021 & _EVAL_826;
  assign _EVAL_2499 = _EVAL_476 & _EVAL_2035;
  assign gateways_gateway_75__EVAL_3 = _EVAL_110;
  assign gateways_gateway_94__EVAL_3 = _EVAL_110;
  assign _EVAL_2616 = _EVAL_195 & _EVAL_3672;
  assign _EVAL_1103 = _EVAL_2150 & _EVAL_2035;
  assign gateways_gateway_27__EVAL_1 = ~_EVAL_2961;
  assign _EVAL_2915 = _EVAL_1880 | gateways_gateway_111__EVAL_4;
  assign gateways_gateway_104__EVAL_2 = _EVAL_2917[105];
  assign gateways_gateway_14__EVAL_1 = ~_EVAL_3213;
  assign gateways_gateway_13__EVAL_1 = ~_EVAL_1120;
  assign _EVAL_3793 = ~_EVAL_2558;
  assign _EVAL_2712 = _EVAL_1181 & _EVAL_826;
  assign fanin__EVAL_1 = _EVAL_2211;
  assign gateways_gateway_5__EVAL_3 = _EVAL_110;
  assign _EVAL_2650 = _EVAL_1670 ? {{29'd0}, _EVAL_2986} : _EVAL_2386;
  assign _EVAL_1755 = _EVAL_615 & _EVAL_3266;
  assign _EVAL_1238 = _EVAL_870 & _EVAL_826;
  assign _EVAL_1074 = _EVAL_195 & _EVAL_2168;
  assign _EVAL_2841 = _EVAL_1151 & _EVAL_826;
  assign gateways_gateway_19__EVAL_2 = _EVAL_2917[20];
  assign _EVAL_2942 = _EVAL_2676 & _EVAL_826;
  assign _EVAL_575 = _EVAL_876 & _EVAL_2035;
  assign gateways_gateway_112__EVAL_0 = _EVAL_9;
  assign _EVAL_2892 = _EVAL_1224 & _EVAL_826;
  assign gateways_gateway_54__EVAL_0 = _EVAL_9;
  assign gateways_gateway_28__EVAL_2 = _EVAL_2917[29];
  assign fanin__EVAL_125 = _EVAL_1876;
  assign _EVAL_1505 = _EVAL_651[24];
  assign _EVAL_161 = _EVAL_1812 ? _EVAL_826 : _EVAL_673;
  assign _EVAL_2525 = 10'h71 == _EVAL_2998;
  assign gateways_gateway_122__EVAL = _EVAL_85;
  assign _EVAL_1700 = &_EVAL_2850;
  assign _EVAL_3802 = _EVAL_2147 & _EVAL_826;
  assign _EVAL_3388 = _EVAL_997 ? _EVAL_826 : _EVAL_2075;
  assign _EVAL_905 = _EVAL_2936 ? {{29'd0}, _EVAL_2981} : _EVAL_2102;
  assign _EVAL_736 = _EVAL_195 & _EVAL_1248;
  assign _EVAL_3148 = _EVAL_651[77];
  assign _EVAL_3304 = ~_EVAL_285;
  assign gateways_gateway_35__EVAL_2 = _EVAL_2917[36];
  assign gateways_gateway_69__EVAL_2 = _EVAL_2917[70];
  assign _EVAL_482 = _EVAL_3349[45];
  assign gateways_gateway_2__EVAL_0 = _EVAL_9;
  assign _EVAL_2517 = _EVAL_3000 & _EVAL_826;
  assign _EVAL_1022 = _EVAL_1738 & _EVAL_2035;
  assign _EVAL_3402 = 10'h19 == _EVAL_2998;
  assign _EVAL_1039 = _EVAL_195 & _EVAL_2624;
  assign _EVAL_1536 = ~_EVAL_2216;
  assign _EVAL_1801 = _EVAL_1649 & _EVAL_3618;
  assign gateways_gateway_9__EVAL_2 = _EVAL_2917[10];
  assign fanin__EVAL_32 = _EVAL_3005;
  assign gateways_gateway__EVAL_3 = _EVAL_110;
  assign _EVAL_2833 = _EVAL_858 | gateways_gateway_102__EVAL_4;
  assign _EVAL_3237 = _EVAL_195 & _EVAL_2220;
  assign _EVAL_1102 = _EVAL_2455 & _EVAL_826;
  assign _EVAL_2263 = _EVAL_1190 | gateways_gateway_21__EVAL_4;
  assign _EVAL_1087 = _EVAL_195 & _EVAL_365;
  assign gateways_gateway_45__EVAL_1 = ~_EVAL_1673;
  assign _EVAL_3340 = _EVAL_195 & _EVAL_1338;
  assign _EVAL_411 = _EVAL_1172 ? _EVAL_826 : _EVAL_645;
  assign gateways_gateway_21__EVAL = _EVAL_46;
  assign _EVAL_1024 = _EVAL_3700 | gateways_gateway_47__EVAL_4;
  assign _EVAL_2922 = _EVAL_2987 & _EVAL_826;
  assign _EVAL_2728 = _EVAL_3029 & _EVAL_826;
  assign _EVAL_1031 = ~_EVAL_482;
  assign _EVAL_588 = out_back__EVAL_12[2];
  assign _EVAL_2122 = _EVAL_842 | gateways_gateway_4__EVAL_4;
  assign gateways_gateway_70__EVAL_3 = _EVAL_110;
  assign _EVAL_333 = _EVAL_1342 & _EVAL_2035;
  assign _EVAL_2667 = _EVAL_2604 | gateways_gateway_98__EVAL_4;
  assign gateways_gateway_58__EVAL_1 = ~_EVAL_1369;
  assign gateways_gateway_16__EVAL_1 = ~_EVAL_2165;
  assign _EVAL_3438 = 10'h5b == _EVAL_2998;
  assign _EVAL_1539 = _EVAL_615 & _EVAL_425;
  assign _EVAL_1953 = _EVAL_3468 & _EVAL_2035;
  assign _EVAL_1170 = _EVAL_651[5];
  assign gateways_gateway_1__EVAL_2 = _EVAL_2917[2];
  assign _EVAL_3081 = _EVAL_195 & _EVAL_3343;
  assign _EVAL_739 = _EVAL_3438 ? _EVAL_826 : _EVAL_2378;
  assign _EVAL_3130 = _EVAL_1707 & _EVAL_826;
  assign gateways_gateway_84__EVAL_3 = _EVAL_110;
  assign gateways_gateway_82__EVAL_2 = _EVAL_2917[83];
  assign _EVAL_3619 = _EVAL_651[115];
  assign gateways_gateway_15__EVAL_2 = _EVAL_2917[16];
  assign _EVAL_723 = _EVAL_1220 & _EVAL_2035;
  assign _EVAL_2738 = 10'h46 == _EVAL_2998;
  assign _EVAL_2671 = _EVAL_195 & _EVAL_3384;
  assign _EVAL_1689 = _EVAL_2264 | gateways_gateway_3__EVAL_4;
  assign _EVAL_3381 = _EVAL_3349[66];
  assign _EVAL_3844 = ~_EVAL_1499;
  assign _EVAL_2274 = 10'h7e == _EVAL_2998;
  assign _EVAL_2918 = _EVAL_959 ? {{29'd0}, _EVAL_1876} : _EVAL_2391;
  assign _EVAL_1547 = 10'h52 == _EVAL_2998;
  assign fanin__EVAL_54 = _EVAL_2711;
  assign _EVAL_3275 = _EVAL_195 & _EVAL_1354;
  assign gateways_gateway_78__EVAL_3 = _EVAL_110;
  assign gateways_gateway_99__EVAL_2 = _EVAL_2917[100];
  assign _EVAL_3214 = {_EVAL_2427,_EVAL_780,_EVAL_2344,_EVAL_2685,_EVAL_3151,_EVAL_276,_EVAL_594,_EVAL_1774,_EVAL_3643,1'h0
    };
  assign gateways_gateway_84__EVAL_2 = _EVAL_2917[85];
  assign gateways_gateway_123__EVAL_3 = _EVAL_110;
  assign _EVAL_1451 = _EVAL_3349[17];
  assign out_back__EVAL_9 = _EVAL_73;
  assign gateways_gateway_15__EVAL_0 = _EVAL_9;
  assign _EVAL_2428 = _EVAL_195 & _EVAL_1852;
  assign _EVAL_826 = _EVAL_2440 == 20'h0;
  assign _EVAL_278 = ~_EVAL_3311;
  assign _EVAL_2722 = _EVAL_955 ? {{29'd0}, _EVAL_692} : _EVAL_1605;
  assign gateways_gateway_22__EVAL_0 = _EVAL_9;
  assign _EVAL_3834 = _EVAL_3417 & _EVAL_826;
  assign _EVAL_3819 = 10'h20 == _EVAL_2998;
  assign fanin__EVAL_84 = _EVAL_1199;
  assign _EVAL_3084 = _EVAL_337 ? {{29'd0}, _EVAL_570} : _EVAL_2020;
  assign _EVAL_1560 = _EVAL_741 & _EVAL_3040;
  assign gateways_gateway_30__EVAL_3 = _EVAL_110;
  assign _EVAL_3166 = {_EVAL_2793,_EVAL_1565,_EVAL_2951,_EVAL_284,_EVAL_3627,_EVAL_3011,_EVAL_3107,_EVAL_2799,_EVAL_267,
    _EVAL_1994};
  assign _EVAL_2205 = _EVAL_3329 ? {{29'd0}, _EVAL_700} : _EVAL_2314;
  assign gateways_gateway_52__EVAL = _EVAL_131;
  assign _EVAL_3706 = _EVAL_849 ? {{29'd0}, _EVAL_3624} : _EVAL_1441;
  assign gateways_gateway_38__EVAL_1 = ~_EVAL_1138;
  assign fanin__EVAL_46 = _EVAL_1528;
  assign gateways_gateway_1__EVAL_0 = _EVAL_9;
  assign _EVAL_3386 = {_EVAL_1847,_EVAL_1434,_EVAL_1347,_EVAL_2961,_EVAL_3263};
  assign _EVAL_3291 = 10'h45 == _EVAL_2998;
  assign _EVAL_1594 = _EVAL_1052 ? _EVAL_826 : _EVAL_3034;
  assign _EVAL_330 = _EVAL_670 & _EVAL_826;
  assign _EVAL_299 = 10'h2b == _EVAL_2998;
  assign _EVAL_1578 = _EVAL_736 & _EVAL_826;
  assign _EVAL_3417 = _EVAL_195 & _EVAL_3524;
  assign gateways_gateway_27__EVAL_2 = _EVAL_2917[28];
  assign gateways_gateway_76__EVAL_0 = _EVAL_9;
  assign _EVAL_632 = _EVAL_282 & _EVAL_2035;
  assign _EVAL_2145 = ~_EVAL_410;
  assign _EVAL_1336 = _EVAL_3557 | gateways_gateway_118__EVAL_4;
  assign _EVAL_3615 = {_EVAL_3627,_EVAL_3011,_EVAL_3107,_EVAL_2799,_EVAL_1127,_EVAL_727,_EVAL_1937,_EVAL_1270,_EVAL_1175
    ,_EVAL_386};
  assign _EVAL_2533 = _EVAL_2936 ? _EVAL_826 : _EVAL_3115;
  assign gateways_gateway_76__EVAL_1 = ~_EVAL_2153;
  assign gateways_gateway_118__EVAL_3 = _EVAL_110;
  assign _EVAL_907 = _EVAL_2320 | gateways_gateway_87__EVAL_4;
  assign _EVAL_3476 = 10'h53 == _EVAL_2998;
  assign _EVAL_2425 = _EVAL_2739 & _EVAL_2035;
  assign _EVAL_3427 = _EVAL_1509 & _EVAL_826;
  assign _EVAL_3209 = _EVAL_638 ? _EVAL_826 : _EVAL_3450;
  assign gateways_gateway_115__EVAL_0 = _EVAL_9;
  assign gateways_gateway_41__EVAL = _EVAL_103;
  assign _EVAL_2252 = _EVAL_195 & _EVAL_2623;
  assign fanin__EVAL_66 = _EVAL_1655;
  assign _EVAL_2391 = _EVAL_1439 ? {{29'd0}, _EVAL_3284} : _EVAL_3075;
  assign _EVAL_374 = 10'h1e == _EVAL_2998;
  assign gateways_gateway_98__EVAL_2 = _EVAL_2917[99];
  assign _EVAL_726 = _EVAL_3349[57];
  assign gateways_gateway_8__EVAL_1 = ~_EVAL_2427;
  assign _EVAL_2945 = _EVAL_651[108];
  assign _EVAL_318 = _EVAL_195 & _EVAL_1830;
  assign _EVAL_772 = _EVAL_3427 & _EVAL_2957;
  assign gateways_gateway_126__EVAL_0 = _EVAL_9;
  assign fanin__EVAL_102 = _EVAL_3835;
  assign _EVAL_1731 = _EVAL_651[32];
  assign _EVAL_1486 = _EVAL_651[98];
  assign _EVAL_3002 = _EVAL_963 | gateways_gateway_14__EVAL_4;
  assign gateways_gateway_82__EVAL_0 = _EVAL_9;
  assign _EVAL_3456 = _EVAL_651[2];
  assign fanin__EVAL_100 = _EVAL_2575;
  assign gateways_gateway_81__EVAL_3 = _EVAL_110;
  assign gateways_gateway_81__EVAL_0 = _EVAL_9;
  assign _EVAL_2279 = _EVAL_195 & _EVAL_1012;
  assign _EVAL_2313 = _EVAL_3089 & _EVAL_826;
  assign gateways_gateway_100__EVAL_3 = _EVAL_110;
  assign gateways_gateway_100__EVAL_2 = _EVAL_2917[101];
  assign _EVAL_3571 = 10'h39 == _EVAL_2998;
  assign _EVAL_1310 = _EVAL_3828 ? {{29'd0}, _EVAL_2384} : _EVAL_3082;
  assign _EVAL_1624 = _EVAL_2904 | gateways_gateway_35__EVAL_4;
  assign _EVAL_1613 = _EVAL_1781 & _EVAL_2035;
  assign _EVAL_488 = 10'h2a == _EVAL_2998;
  assign _EVAL_3566 = 10'h6b == _EVAL_2998;
  assign _EVAL_1763 = _EVAL_651[125];
  assign _EVAL_2861 = _EVAL_3828 ? _EVAL_826 : _EVAL_2565;
  assign _EVAL_2191 = _EVAL_2465 & _EVAL_826;
  assign _EVAL_3455 = _EVAL_171 ? {{29'd0}, _EVAL_2211} : _EVAL_1310;
  assign _EVAL_2862 = out_back__EVAL_12[0];
  assign _EVAL_2144 = _EVAL_195 & _EVAL_1544;
  assign gateways_gateway_75__EVAL = _EVAL_129;
  assign _EVAL_3328 = _EVAL_1761 & _EVAL_826;
  assign gateways_gateway_9__EVAL_3 = _EVAL_110;
  assign _EVAL_1683 = ~_EVAL_753;
  assign _EVAL_1118 = 10'h28 == _EVAL_2998;
  assign _EVAL_3704 = _EVAL_3349[35];
  assign _EVAL_2249 = _EVAL_2989 & _EVAL_826;
  assign gateways_gateway_26__EVAL_0 = _EVAL_9;
  assign fanin__EVAL_118 = _EVAL_3711;
  assign gateways_gateway_2__EVAL_1 = ~_EVAL_594;
  assign gateways_gateway_84__EVAL = _EVAL_39;
  assign _EVAL_1010 = ~_EVAL_2788;
  assign _EVAL_342 = _EVAL_841 & _EVAL_826;
  assign gateways_gateway_114__EVAL_0 = _EVAL_9;
  assign gateways_gateway_98__EVAL_1 = ~_EVAL_3395;
  assign _EVAL_3686 = _EVAL_257 | gateways_gateway_85__EVAL_4;
  assign _EVAL_320 = _EVAL_1757 & _EVAL_2035;
  assign _EVAL_3102 = _EVAL_1438 ? {{29'd0}, _EVAL_2531} : _EVAL_1661;
  assign _EVAL_1172 = 10'h43 == _EVAL_2998;
  assign _EVAL_272 = _EVAL_3349[6];
  assign _EVAL_322 = ~_EVAL_3811;
  assign _EVAL_886 = _EVAL_195 & _EVAL_1780;
  assign _EVAL_3363 = _EVAL_856 ? _EVAL_826 : _EVAL_2462;
  assign _EVAL_3467 = 10'h5c == _EVAL_2998;
  assign gateways_gateway_88__EVAL_2 = _EVAL_2917[89];
  assign _EVAL_3412 = {_EVAL_202,_EVAL_1116,_EVAL_1948,_EVAL_3803,_EVAL_2193,_EVAL_2618,_EVAL_414,_EVAL_3366};
  assign _EVAL_2747 = _EVAL_651[96];
  assign _EVAL_585 = ~_EVAL_3700;
  assign gateways_gateway_57__EVAL_1 = ~_EVAL_3508;
  assign _EVAL_1020 = ~_EVAL_801;
  assign _EVAL_1976 = _EVAL_3587 & _EVAL_826;
  assign _EVAL_2881 = 10'h3c == _EVAL_2998;
  assign _EVAL_1957 = ~_EVAL_1485;
  assign _EVAL_569 = _EVAL_1017 ? {{29'd0}, _EVAL_1789} : _EVAL_313;
  assign _EVAL_1174 = 10'h18 == _EVAL_2998;
  assign gateways_gateway_65__EVAL_0 = _EVAL_9;
  assign gateways_gateway_8__EVAL = _EVAL_78;
  assign _EVAL_356 = _EVAL_3409 & _EVAL_2035;
  assign _EVAL_2855 = _EVAL_651[18];
  assign _EVAL_281 = 10'h2f == _EVAL_2998;
  assign gateways_gateway_58__EVAL_0 = _EVAL_9;
  assign _EVAL_1269 = _EVAL_3349[9];
  assign _EVAL_3480 = _EVAL_195 & _EVAL_2874;
  assign gateways_gateway_29__EVAL_0 = _EVAL_9;
  assign _EVAL_2784 = _EVAL_1367 ? _EVAL_826 : _EVAL_1593;
  assign _EVAL_1191 = _EVAL_3349[40];
  assign _EVAL_425 = &_EVAL_1016;
  assign gateways_gateway_103__EVAL_0 = _EVAL_9;
  assign fanin__EVAL_79 = _EVAL_1796;
  assign _EVAL_3104 = _EVAL_3349[109];
  assign _EVAL_353 = _EVAL_3219 & _EVAL_826;
  assign gateways_gateway_95__EVAL_2 = _EVAL_2917[96];
  assign _EVAL_1255 = _EVAL_1764 | gateways_gateway_40__EVAL_4;
  assign _EVAL_2054 = _EVAL_2133 & _EVAL_2035;
  assign _EVAL_695 = 10'h40 == _EVAL_2998;
  assign _EVAL_3644 = {_EVAL_2719,_EVAL_2509,_EVAL_1365,_EVAL_2737,_EVAL_811,_EVAL_3440,_EVAL_3387,_EVAL_3305,_EVAL_770,
    _EVAL_526};
  assign _EVAL_2779 = ~_EVAL_471;
  assign gateways_gateway_2__EVAL_3 = _EVAL_110;
  assign _EVAL_2832 = _EVAL_2017 | gateways_gateway_117__EVAL_4;
  assign gateways_gateway_6__EVAL_3 = _EVAL_110;
  assign _EVAL_3806 = _EVAL_651[50];
  assign _EVAL_2742 = _EVAL_2803 ? _EVAL_826 : _EVAL_3564;
  assign _EVAL_1237 = _EVAL_195 & _EVAL_2027;
  assign _EVAL_3142 = _EVAL_195 & _EVAL_3148;
  assign _EVAL_1440 = _EVAL_195 & _EVAL_3681;
  assign _EVAL_3568 = _EVAL_1809 ? {{29'd0}, _EVAL_2306} : _EVAL_2034;
  assign fanin__EVAL_67 = _EVAL_3559;
  assign _EVAL_3317 = _EVAL_1451 | gateways_gateway_16__EVAL_4;
  assign _EVAL_1411 = _EVAL_2123 ? _EVAL_2757 : 7'h0;
  assign _EVAL_2366 = _EVAL_3349[62];
  assign gateways_gateway_97__EVAL_0 = _EVAL_9;
  assign _EVAL_496 = _EVAL_3349[68];
  assign _EVAL_378 = _EVAL_195 & _EVAL_1942;
  assign _EVAL_166 = 10'h7 == _EVAL_2998;
  assign _EVAL_2965 = _EVAL_1867 ? _EVAL_826 : _EVAL_2720;
  assign gateways_gateway_117__EVAL_0 = _EVAL_9;
  assign gateways_gateway_25__EVAL_3 = _EVAL_110;
  assign _EVAL_2999 = _EVAL_3391 ? _EVAL_826 : _EVAL_2586;
  assign out_back__EVAL_10 = _EVAL_101;
  assign _EVAL_2686 = _EVAL_3349[28];
  assign _EVAL_2284 = _EVAL_3337 ? {{29'd0}, _EVAL_2753} : _EVAL_2871;
  assign gateways_gateway_25__EVAL_0 = _EVAL_9;
  assign _EVAL_1969 = ~_EVAL_2860;
  assign _EVAL_3123 = 10'h201 == _EVAL_2998;
  assign _EVAL_2852 = _EVAL_2696 & _EVAL_826;
  assign _EVAL_1359 = _EVAL_1499 | gateways_gateway_48__EVAL_4;
  assign gateways_gateway_3__EVAL_2 = _EVAL_2917[4];
  assign _EVAL_3299 = 10'h1b == _EVAL_2998;
  assign _EVAL_232 = _EVAL_2098 & _EVAL_826;
  assign fanin__EVAL_128 = _EVAL_1771;
  assign _EVAL_3555 = _EVAL_3577 & _EVAL_2035;
  assign _EVAL_696 = _EVAL_849 ? _EVAL_826 : _EVAL_1288;
  assign gateways_gateway_72__EVAL_2 = _EVAL_2917[73];
  assign _EVAL_2693 = 10'h27 == _EVAL_2998;
  assign _EVAL_1518 = _EVAL_1740 & _EVAL_826;
  assign _EVAL_3633 = _EVAL_3349[21];
  assign _EVAL_231 = ~_EVAL_3716;
  assign _EVAL_3548 = 10'h74 == _EVAL_2998;
  assign _EVAL_595 = 10'hb == _EVAL_2998;
  assign gateways_gateway_126__EVAL = _EVAL_3;
  assign gateways_gateway_106__EVAL_3 = _EVAL_110;
  assign gateways_gateway_107__EVAL_1 = ~_EVAL_872;
  assign gateways_gateway_54__EVAL_2 = _EVAL_2917[55];
  assign gateways_gateway_79__EVAL_2 = _EVAL_2917[80];
  assign gateways_gateway_95__EVAL_0 = _EVAL_9;
  assign _EVAL_1499 = _EVAL_3349[49];
  assign _EVAL_2231 = ~_EVAL_1428;
  assign _EVAL_2868 = 10'h79 == _EVAL_2998;
  assign _EVAL_1535 = _EVAL_2692 & _EVAL_2035;
  assign gateways_gateway_73__EVAL = _EVAL_34;
  assign gateways_gateway_82__EVAL_1 = ~_EVAL_1175;
  assign _EVAL_3504 = 10'h56 == _EVAL_2998;
  assign _EVAL_2896 = _EVAL_1292 | gateways_gateway_82__EVAL_4;
  assign _EVAL_2140 = _EVAL_3571 ? {{29'd0}, _EVAL_1988} : _EVAL_3017;
  assign _EVAL_2059 = _EVAL_2408 ? {{29'd0}, _EVAL_3744} : _EVAL_1008;
  assign gateways_gateway_77__EVAL_0 = _EVAL_9;
  assign _EVAL_2577 = _EVAL_2202 & _EVAL_2035;
  assign gateways_gateway_13__EVAL_0 = _EVAL_9;
  assign _EVAL_3610 = _EVAL_1541 | gateways_gateway_38__EVAL_4;
  assign _EVAL_921 = out_back__EVAL_3[0];
  assign gateways_gateway_14__EVAL_2 = _EVAL_2917[15];
  assign gateways_gateway_120__EVAL_3 = _EVAL_110;
  assign _EVAL_385 = 10'h200 == _EVAL_2998;
  assign _EVAL_909 = {_EVAL_2618,_EVAL_414,_EVAL_3366,_EVAL_3589,_EVAL_2396,_EVAL_1872,_EVAL_872,_EVAL_3043,_EVAL_168,
    _EVAL_224};
  assign _EVAL_1338 = _EVAL_651[113];
  assign _EVAL_3171 = _EVAL_3349[80];
  assign _EVAL_1688 = _EVAL_3244 & _EVAL_826;
  assign _EVAL_1787 = _EVAL_651[28];
  assign _EVAL_2617 = _EVAL_195 & _EVAL_1644;
  assign _EVAL_3105 = _EVAL_3349[96];
  assign _EVAL_787 = _EVAL_1485 | gateways_gateway_109__EVAL_4;
  assign _EVAL_3027 = ~_EVAL_2527;
  assign _EVAL_2348 = _EVAL_1191 | gateways_gateway_39__EVAL_4;
  assign _EVAL_1012 = _EVAL_651[118];
  assign gateways_gateway_19__EVAL_0 = _EVAL_9;
  assign _EVAL_3530 = _EVAL_1346 | gateways_gateway_110__EVAL_4;
  assign _EVAL_1534 = _EVAL_1824 ? _EVAL_826 : _EVAL_544;
  assign _EVAL_3241 = _EVAL_2862 ? 8'hff : 8'h0;
  assign _EVAL_3111 = _EVAL_1892 & _EVAL_826;
  assign _EVAL_3716 = _EVAL_3349[85];
  assign _EVAL_2375 = _EVAL_651[46];
  assign _EVAL_3708 = _EVAL_2970 ? _EVAL_826 : _EVAL_3307;
  assign _EVAL_1960 = _EVAL_195 & _EVAL_506;
  assign fanin__EVAL_24 = _EVAL_2982;
  assign fanin__EVAL_8 = _EVAL_2986;
  assign fanin__EVAL_107 = _EVAL_2988;
  assign _EVAL_3404 = _EVAL_3322 ? {{29'd0}, _EVAL_3218} : _EVAL_3848;
  assign gateways_gateway_94__EVAL_0 = _EVAL_9;
  assign _EVAL_1597 = _EVAL_3220 & _EVAL_826;
  assign _EVAL_3596 = 10'h77 == _EVAL_2998;
  assign _EVAL_1148 = _EVAL_1430 | gateways_gateway_107__EVAL_4;
  assign _EVAL_2431 = ~_EVAL_258;
  assign _EVAL_2593 = _EVAL_886 & _EVAL_826;
  assign _EVAL_3576 = _EVAL_3171 | gateways_gateway_79__EVAL_4;
  assign gateways_gateway_117__EVAL_1 = ~_EVAL_1116;
  assign fanin__EVAL_69 = _EVAL_1963;
  assign _EVAL_1398 = _EVAL_540 & _EVAL_826;
  assign _EVAL_903 = _EVAL_651[116];
  assign _EVAL_2601 = ~_EVAL_362;
  assign _EVAL_335 = _EVAL_873 & _EVAL_2035;
  assign _EVAL_1905 = _EVAL_1788 & _EVAL_2035;
  assign _EVAL_2805 = ~_EVAL_2316;
  assign _EVAL_3747 = _EVAL_651[89];
  assign gateways_gateway_89__EVAL_1 = ~_EVAL_3011;
  assign _EVAL_412 = _EVAL_404 ? _EVAL_826 : _EVAL_3363;
  assign _EVAL_1286 = ~_EVAL_643;
  assign _EVAL_170 = _EVAL_2347 ? {{29'd0}, _EVAL_936} : _EVAL_3568;
  assign gateways_gateway_83__EVAL_3 = _EVAL_110;
  assign _EVAL_3174 = _EVAL_3349[92];
  assign _EVAL_3560 = _EVAL_3337 ? _EVAL_826 : _EVAL_2008;
  assign _EVAL_876 = _EVAL_1946 & _EVAL_826;
  assign _EVAL_3038 = _EVAL_2850[15:8];
  assign gateways_gateway_67__EVAL_1 = ~_EVAL_3440;
  assign gateways_gateway_81__EVAL_1 = ~_EVAL_1507;
  assign _EVAL_254 = _EVAL_2322 | gateways_gateway_71__EVAL_4;
  assign gateways_gateway_1__EVAL = _EVAL_72;
  assign _EVAL_176 = 10'h7a == _EVAL_2998;
  assign _EVAL_1541 = _EVAL_3349[39];
  assign gateways_gateway_50__EVAL_2 = _EVAL_2917[51];
  assign _EVAL_2770 = _EVAL_2282 | gateways_gateway_58__EVAL_4;
  assign _EVAL_1608 = _EVAL_3438 ? {{29'd0}, _EVAL_1621} : _EVAL_1088;
  assign fanin__EVAL_41 = _EVAL_3657;
  assign _EVAL_504 = 10'h24 == _EVAL_2998;
  assign _EVAL_3579 = _EVAL_1506 ? _EVAL_826 : _EVAL_739;
  assign _EVAL_195 = _EVAL_2088 & _EVAL_3667;
  assign _EVAL_1997 = _EVAL_3533 ? {{29'd0}, _EVAL_3290} : _EVAL_3430;
  assign fanin__EVAL_71 = _EVAL_3357;
  assign _EVAL_241 = _EVAL_2974 ? _EVAL_826 : _EVAL_2236;
  assign _EVAL_1183 = _EVAL_3349[75];
  assign _EVAL_3683 = _EVAL_3782 | gateways_gateway_116__EVAL_4;
  assign _EVAL_3236 = 10'h1a == _EVAL_2998;
  assign gateways_gateway_16__EVAL_3 = _EVAL_110;
  assign _EVAL_343 = _EVAL_571 | gateways_gateway_77__EVAL_4;
  assign gateways_gateway_40__EVAL_1 = ~_EVAL_3770;
  assign gateways_gateway_119__EVAL_1 = ~_EVAL_965;
  assign gateways_gateway_45__EVAL_2 = _EVAL_2917[46];
  assign gateways_gateway_90__EVAL_0 = _EVAL_9;
  assign _EVAL_3593 = _EVAL_1512 | gateways_gateway_1__EVAL_4;
  assign gateways_gateway_34__EVAL = _EVAL_33;
  assign gateways_gateway_9__EVAL_1 = ~_EVAL_2627;
  assign fanin__EVAL_90 = _EVAL_1745;
  assign gateways_gateway_93__EVAL_2 = _EVAL_2917[94];
  assign _EVAL_1433 = 10'h65 == _EVAL_2998;
  assign gateways_gateway_19__EVAL_3 = _EVAL_110;
  assign _EVAL_1869 = 10'h3b == _EVAL_2998;
  assign gateways_gateway_120__EVAL_0 = _EVAL_9;
  assign _EVAL_2936 = 10'h6f == _EVAL_2998;
  assign fanin__EVAL_105 = _EVAL_2004;
  assign gateways_gateway_59__EVAL_1 = ~_EVAL_1392;
  assign _EVAL_2985 = 10'h1c == _EVAL_2998;
  assign _EVAL_827 = _EVAL_3716 | gateways_gateway_84__EVAL_4;
  assign _EVAL_862 = _EVAL_3067 & _EVAL_2035;
  assign _EVAL_1987 = 10'h5 == _EVAL_2998;
  assign _EVAL_265 = _EVAL_3322 ? _EVAL_826 : _EVAL_1056;
  assign _EVAL_975 = _EVAL_584 ? _EVAL_826 : _EVAL_3603;
  assign gateways_gateway_52__EVAL_1 = ~_EVAL_1749;
  assign _EVAL_3246 = _EVAL_3349[64];
  assign fanin__EVAL_64 = _EVAL_1634;
  assign _EVAL_1401 = _EVAL_1014 & _EVAL_2035;
  assign _EVAL_293 = _EVAL_2009 ? {{29'd0}, _EVAL_1407} : _EVAL_2946;
  assign _EVAL_2622 = _EVAL_3349[16];
  assign gateways_gateway_111__EVAL = _EVAL_23;
  assign _EVAL_2097 = _EVAL_3646 & _EVAL_2035;
  assign gateways_gateway_2__EVAL = _EVAL_18;
  assign _EVAL_1779 = _EVAL_2970 ? {{29'd0}, _EVAL_222} : _EVAL_2059;
  assign _EVAL_1540 = _EVAL_1438 ? _EVAL_826 : _EVAL_2417;
  assign gateways_gateway_116__EVAL_2 = _EVAL_2917[117];
  assign _EVAL_524 = _EVAL_3548 ? {{29'd0}, _EVAL_3446} : _EVAL_2791;
  assign _EVAL_1346 = _EVAL_3349[111];
  assign gateways_gateway_11__EVAL_1 = ~_EVAL_552;
  assign _EVAL_2438 = _EVAL_195 & _EVAL_2983;
  assign gateways_gateway_16__EVAL = _EVAL_86;
  assign _EVAL_679 = ~_EVAL_2196;
  assign _EVAL_1880 = _EVAL_3349[112];
  assign _EVAL_1733 = _EVAL_368 | gateways_gateway_75__EVAL_4;
  assign gateways_gateway_20__EVAL_1 = ~_EVAL_1467;
  assign _EVAL_820 = _EVAL_3349[74];
  assign _EVAL_47 = out_back__EVAL_7;
  assign fanin__EVAL_20 = _EVAL_1569;
  assign _EVAL_1886 = _EVAL_2515 & _EVAL_2035;
  assign _EVAL_510 = _EVAL_615 & _EVAL_2957;
  assign _EVAL_1158 = _EVAL_195 & _EVAL_3637;
  assign gateways_gateway_11__EVAL = _EVAL_11;
  assign _EVAL_274 = _EVAL_3349[24];
  assign gateways_gateway_63__EVAL_3 = _EVAL_110;
  assign _EVAL_1680 = _EVAL_195 & _EVAL_2375;
  assign _EVAL_3288 = _EVAL_422 & _EVAL_826;
  assign _EVAL_1180 = _EVAL_3349[71];
  assign gateways_gateway_121__EVAL_2 = _EVAL_2917[122];
  assign _EVAL_2087 = _EVAL_324 & _EVAL_2035;
  assign fanin__EVAL_14 = _EVAL_3505;
  assign _EVAL_592 = _EVAL_185 ? _EVAL_826 : _EVAL_1534;
  assign gateways_gateway_30__EVAL = _EVAL_68;
  assign _EVAL_3008 = _EVAL_1579 & _EVAL_2035;
  assign _EVAL_2236 = _EVAL_2308 ? _EVAL_826 : _EVAL_2312;
  assign _EVAL_3461 = _EVAL_3537 ? _EVAL_3386 : _EVAL_500;
  assign _EVAL_689 = _EVAL_3476 ? {{29'd0}, _EVAL_2853} : _EVAL_1678;
  assign _EVAL_534 = _EVAL_2005 | gateways_gateway_6__EVAL_4;
  assign _EVAL_462 = ~_EVAL_2341;
  assign _EVAL_2979 = {_EVAL_1471,_EVAL_2070,_EVAL_2418,_EVAL_1517};
  assign _EVAL_1591 = _EVAL_593 & _EVAL_2035;
  assign _EVAL_2257 = _EVAL_3490 & _EVAL_826;
  assign _EVAL_212 = _EVAL_651[259];
  assign gateways_gateway_109__EVAL_1 = ~_EVAL_2396;
  assign _EVAL_340 = _EVAL_651[111];
  assign _EVAL_2473 = _EVAL_195 & _EVAL_184;
  assign gateways_gateway_78__EVAL_2 = _EVAL_2917[79];
  assign gateways_gateway_37__EVAL = _EVAL_65;
  assign _EVAL_2810 = _EVAL_195 & _EVAL_1956;
  assign gateways_gateway_88__EVAL_3 = _EVAL_110;
  assign _EVAL_2992 = _EVAL_176 ? _EVAL_826 : _EVAL_2589;
  assign _EVAL_590 = _EVAL_3597 & _EVAL_2035;
  assign gateways_gateway_44__EVAL_1 = ~_EVAL_1944;
  assign _EVAL_2043 = _EVAL_1043 | gateways_gateway_83__EVAL_4;
  assign _EVAL_992 = ~_EVAL_1762;
  assign _EVAL_2102 = _EVAL_1482 ? {{29'd0}, _EVAL_3191} : _EVAL_2069;
  assign fanin__EVAL_42 = _EVAL_2873;
  assign _EVAL_368 = _EVAL_3349[76];
  assign _EVAL_2483 = ~_EVAL_1601;
  assign _EVAL_1439 = 10'h35 == _EVAL_2998;
  assign _EVAL_3489 = _EVAL_651[81];
  assign _EVAL_2171 = _EVAL_1554 ? {{29'd0}, _EVAL_642} : _EVAL_547;
  assign gateways_gateway_89__EVAL_3 = _EVAL_110;
  assign _EVAL_1554 = 10'h49 == _EVAL_2998;
  assign fanin__EVAL_74 = _EVAL_1459;
  assign _EVAL_520 = _EVAL_3349[38];
  assign _EVAL_3367 = 10'h1 == _EVAL_2998;
  assign gateways_gateway_108__EVAL = _EVAL_38;
  assign _EVAL_2094 = _EVAL_3270 ? _EVAL_826 : _EVAL_334;
  assign _EVAL_1783 = ~_EVAL_2907;
  assign _EVAL_2347 = 10'h13 == _EVAL_2998;
  assign gateways_gateway__EVAL = _EVAL_49;
  assign _EVAL_3069 = _EVAL_385 ? _EVAL_826 : _EVAL_2710;
  assign _EVAL_547 = _EVAL_860 ? {{29'd0}, _EVAL_3469} : _EVAL_1076;
  assign gateways_gateway_87__EVAL_0 = _EVAL_9;
  assign _EVAL_285 = _EVAL_3349[25];
  assign _EVAL_571 = _EVAL_3349[78];
  assign gateways_gateway_1__EVAL_1 = ~_EVAL_1774;
  assign gateways_gateway_12__EVAL_0 = _EVAL_9;
  assign _EVAL_1071 = _EVAL_3391 ? {{29'd0}, _EVAL_3315} : _EVAL_3743;
  assign _EVAL_3588 = _EVAL_651[14];
  assign fanin__EVAL_12 = _EVAL_3072;
  assign _EVAL_1430 = _EVAL_3349[108];
  assign gateways_gateway_96__EVAL_3 = _EVAL_110;
  assign gateways_gateway_85__EVAL_1 = ~_EVAL_727;
  assign _EVAL_3037 = _EVAL_3374 & _EVAL_826;
  assign _EVAL_3618 = _EVAL_651[513];
  assign _EVAL_1146 = _EVAL_615 & _EVAL_678;
  assign gateways_gateway_125__EVAL_3 = _EVAL_110;
  assign _EVAL_2159 = ~_EVAL_916;
  assign _EVAL_3454 = _EVAL_3256 ? {{29'd0}, _EVAL_1655} : _EVAL_1093;
  assign _EVAL_917 = _EVAL_614 & _EVAL_2035;
  assign _EVAL_3101 = _EVAL_3329 ? _EVAL_826 : _EVAL_828;
  assign _EVAL_851 = _EVAL_196 & _EVAL_2035;
  assign _EVAL_280 = _EVAL_2482 | gateways_gateway_45__EVAL_4;
  assign _EVAL_3219 = _EVAL_195 & _EVAL_3211;
  assign _EVAL_890 = ~_EVAL_2017;
  assign _EVAL_777 = _EVAL_1081 & _EVAL_2035;
  assign gateways_gateway_115__EVAL = _EVAL_121;
  assign _EVAL_1532 = _EVAL_651[56];
  assign _EVAL_2098 = _EVAL_195 & _EVAL_1973;
  assign _EVAL_490 = _EVAL_2788 | gateways_gateway_59__EVAL_4;
  assign gateways_gateway_18__EVAL_1 = ~_EVAL_498;
  assign gateways_gateway_90__EVAL_3 = _EVAL_110;
  assign _EVAL_3157 = _EVAL_3114 & _EVAL_826;
  assign _EVAL_3639 = ~_EVAL_571;
  assign _EVAL_3318 = _EVAL_2179 & _EVAL_826;
  assign _EVAL_996 = _EVAL_195 & _EVAL_2945;
  assign fanin__EVAL_33 = _EVAL_2518;
  assign gateways_gateway_38__EVAL_0 = _EVAL_9;
  assign gateways_gateway_38__EVAL = _EVAL_13;
  assign gateways_gateway_54__EVAL_1 = ~_EVAL_3346;
  assign _EVAL_151 = _EVAL_3007 & _EVAL_2035;
  assign _EVAL_1500 = 10'h17 == _EVAL_2998;
  assign gateways_gateway_33__EVAL_1 = ~_EVAL_2668;
  assign _EVAL_2346 = _EVAL_651[106];
  assign _EVAL_1000 = _EVAL_1902 ? {{29'd0}, _EVAL_1745} : _EVAL_978;
  assign _EVAL_844 = _EVAL_651[9];
  assign gateways_gateway_118__EVAL_1 = ~_EVAL_202;
  assign _EVAL_1752 = _EVAL_2366 | gateways_gateway_61__EVAL_4;
  assign _EVAL_2298 = _EVAL_3349[102];
  assign _EVAL_845 = {_EVAL_3420,_EVAL_3331,_EVAL_350,_EVAL_1392,_EVAL_1866};
  assign gateways_gateway_24__EVAL_0 = _EVAL_9;
  assign _EVAL_1762 = _EVAL_3349[114];
  assign _EVAL_2822 = _EVAL_3349[31];
  assign gateways_gateway_46__EVAL_3 = _EVAL_110;
  assign _EVAL_3762 = _EVAL_847 & _EVAL_826;
  assign _EVAL_3358 = _EVAL_3800 & _EVAL_826;
  assign gateways_gateway_85__EVAL = _EVAL_4;
  assign _EVAL_467 = _EVAL_2980 & _EVAL_826;
  assign _EVAL_338 = _EVAL_651[31];
  assign _EVAL_3359 = _EVAL_3328 & _EVAL_678;
  assign gateways_gateway_32__EVAL_3 = _EVAL_110;
  assign _EVAL_2149 = _EVAL_2279 & _EVAL_826;
  assign fanin__EVAL_119 = _EVAL_456;
  assign gateways_gateway_15__EVAL_3 = _EVAL_110;
  assign _EVAL_2700 = _EVAL_2251 | gateways_gateway_124__EVAL_4;
  assign _EVAL_2889 = {_EVAL_3213,_EVAL_1120,_EVAL_3824,_EVAL_552,_EVAL_3140,_EVAL_2627,_EVAL_2427,_EVAL_780,_EVAL_3475}
    ;
  assign _EVAL_1002 = _EVAL_195 & _EVAL_160;
  assign gateways_gateway_4__EVAL_3 = _EVAL_110;
  assign fanin__EVAL_30 = _EVAL_692;
  assign _EVAL_2987 = _EVAL_195 & _EVAL_3167;
  assign _EVAL_206 = _EVAL_195 & _EVAL_3165;
  assign _EVAL_1438 = 10'h25 == _EVAL_2998;
  assign gateways_gateway_1__EVAL_3 = _EVAL_110;
  assign _EVAL_3468 = _EVAL_318 & _EVAL_826;
  assign _EVAL_1485 = _EVAL_3349[110];
  assign gateways_gateway_113__EVAL_3 = _EVAL_110;
  assign _EVAL_2296 = {_EVAL_1471,_EVAL_2070,_EVAL_2418,_EVAL_1517,_EVAL_1340,_EVAL_1380,_EVAL_394,_EVAL_2877,_EVAL_2902
    };
  assign gateways_gateway_4__EVAL_2 = _EVAL_2917[5];
  assign fanin__EVAL_21 = _EVAL_167;
  assign gateways_gateway_7__EVAL_3 = _EVAL_110;
  assign gateways_gateway_111__EVAL_1 = ~_EVAL_3366;
  assign _EVAL_3182 = _EVAL_1278 & _EVAL_2035;
  assign _EVAL_3840 = _EVAL_784 & _EVAL_2035;
  assign _EVAL_2106 = ~_EVAL_274;
  assign gateways_gateway_104__EVAL_1 = ~_EVAL_2698;
  assign _EVAL_177 = _EVAL_496 | gateways_gateway_67__EVAL_4;
  assign _EVAL_712 = ~_EVAL_605;
  assign _EVAL_3538 = _EVAL_195 & _EVAL_3729;
  assign _EVAL_3394 = _EVAL_1367 ? {{29'd0}, _EVAL_3737} : _EVAL_1241;
  assign gateways_gateway_85__EVAL_0 = _EVAL_9;
  assign fanin__EVAL_58 = _EVAL_3342;
  assign _EVAL_1882 = _EVAL_1867 ? {{29'd0}, _EVAL_2012} : _EVAL_449;
  assign gateways_gateway_115__EVAL_2 = _EVAL_2917[116];
  assign _EVAL_1923 = 10'h76 == _EVAL_2998;
  assign _EVAL_2888 = _EVAL_2812 | gateways_gateway_123__EVAL_4;
  assign _EVAL_1702 = _EVAL_2868 ? {{29'd0}, _EVAL_1085} : _EVAL_2549;
  assign _EVAL_1144 = _EVAL_487 & _EVAL_826;
  assign gateways_gateway_112__EVAL = _EVAL_105;
  assign _EVAL_476 = _EVAL_206 & _EVAL_826;
  assign _EVAL_2772 = _EVAL_3349[121];
  assign _EVAL_1088 = _EVAL_3467 ? {{29'd0}, _EVAL_707} : _EVAL_1966;
  assign gateways_gateway_4__EVAL = _EVAL_7;
  assign _EVAL_1435 = 10'h2e == _EVAL_2998;
  assign gateways_gateway_108__EVAL_1 = ~_EVAL_1872;
  assign _EVAL_889 = ~_EVAL_2282;
  assign _EVAL_1681 = _EVAL_1900 & _EVAL_826;
  assign _EVAL_970 = _EVAL_1884 ? {{29'd0}, _EVAL_456} : _EVAL_2204;
  assign _EVAL_2549 = _EVAL_176 ? {{29'd0}, _EVAL_2996} : _EVAL_3077;
  assign _EVAL_1595 = _EVAL_3047 ? _EVAL_826 : _EVAL_3259;
  assign _EVAL_1101 = _EVAL_3142 & _EVAL_826;
  assign fanin__EVAL_109 = _EVAL_2828;
  assign gateways_gateway_11__EVAL_2 = _EVAL_2917[12];
  assign _EVAL_1267 = _EVAL_1578 & _EVAL_2035;
  assign _EVAL_3221 = 10'h51 == _EVAL_2998;
  assign _EVAL_489 = _EVAL_1144 & _EVAL_2035;
  assign gateways_gateway_55__EVAL = _EVAL_107;
  assign gateways_gateway_126__EVAL_1 = ~_EVAL_1710;
  assign _EVAL_2860 = _EVAL_3349[34];
  assign gateways_gateway_59__EVAL_2 = _EVAL_2917[60];
  assign gateways_gateway__EVAL_1 = ~_EVAL_3643;
  assign _EVAL_3692 = _EVAL_185 ? {{29'd0}, _EVAL_517} : _EVAL_3198;
  assign _EVAL_3409 = _EVAL_3612 & _EVAL_826;
  assign _EVAL_3732 = _EVAL_651[73];
  assign gateways_gateway_80__EVAL_2 = _EVAL_2917[81];
  assign gateways_gateway_2__EVAL_2 = _EVAL_2917[3];
  assign gateways_gateway_25__EVAL = _EVAL_111;
  assign gateways_gateway_70__EVAL_0 = _EVAL_9;
  assign gateways_gateway_40__EVAL_3 = _EVAL_110;
  assign fanin__EVAL_116 = _EVAL_1134;
  assign _EVAL_3528 = _EVAL_2009 ? _EVAL_826 : _EVAL_3695;
  assign gateways_gateway_119__EVAL_2 = _EVAL_2917[120];
  assign _EVAL_416 = _EVAL_651[124];
  assign _EVAL_2074 = _EVAL_1500 ? _EVAL_826 : _EVAL_1034;
  assign _EVAL_2152 = _EVAL_651[62];
  assign gateways_gateway_107__EVAL_0 = _EVAL_9;
  assign _EVAL_3071 = _EVAL_2428 & _EVAL_826;
  assign _EVAL_1342 = _EVAL_1087 & _EVAL_826;
  assign fanin__EVAL_51 = _EVAL_1252;
  assign _EVAL_2629 = _EVAL_3426 | gateways_gateway_42__EVAL_4;
  assign gateways_gateway_71__EVAL_3 = _EVAL_110;
  assign gateways_gateway_102__EVAL = _EVAL_15;
  assign gateways_gateway_35__EVAL = _EVAL_132;
  assign gateways_gateway_68__EVAL_0 = _EVAL_9;
  assign _EVAL_2732 = ~_EVAL_2264;
  assign _EVAL_3772 = _EVAL_281 ? _EVAL_826 : _EVAL_2763;
  assign gateways_gateway_112__EVAL_2 = _EVAL_2917[113];
  assign _EVAL_1248 = _EVAL_651[34];
  assign _EVAL_2998 = {_EVAL_2227,_EVAL_1178,_EVAL_1239,_EVAL_2490,_EVAL_792,_EVAL_3147,_EVAL_1550,_EVAL_2023,_EVAL_2660
    ,_EVAL_921};
  assign _EVAL_1419 = _EVAL_1418 ? _EVAL_826 : _EVAL_412;
  assign _EVAL_2027 = _EVAL_651[95];
  assign gateways_gateway_62__EVAL_0 = _EVAL_9;
  assign gateways_gateway_22__EVAL_1 = ~_EVAL_1964;
  assign _EVAL_3572 = _EVAL_651[51];
  assign _EVAL_954 = _EVAL_2349 ? _EVAL_826 : _EVAL_2521;
  assign _EVAL_3161 = _EVAL_751 & _EVAL_826;
  assign gateways_gateway_3__EVAL_1 = ~_EVAL_276;
  assign _EVAL_3564 = _EVAL_1869 ? _EVAL_826 : _EVAL_3474;
  assign _EVAL_1418 = 10'h4e == _EVAL_2998;
  assign gateways_gateway_108__EVAL_3 = _EVAL_110;
  assign _EVAL_2361 = _EVAL_499 ? _EVAL_2576 : _EVAL_190;
  assign gateways_gateway_37__EVAL_0 = _EVAL_9;
  assign fanin__EVAL_43 = _EVAL_570;
  assign _EVAL_2576 = {_EVAL_2793,_EVAL_1565,_EVAL_2951,_EVAL_284,_EVAL_3615};
  assign _EVAL_1658 = _EVAL_3122 | gateways_gateway_106__EVAL_4;
  assign _EVAL_2315 = _EVAL_3523 | gateways_gateway_55__EVAL_4;
  assign _EVAL_602 = _EVAL_195 & _EVAL_3806;
  assign _EVAL_1879 = 10'h23 == _EVAL_2998;
  assign _EVAL_2659 = _EVAL_3548 ? _EVAL_826 : _EVAL_1594;
  assign _EVAL_1314 = ~_EVAL_1413;
  assign _EVAL_3015 = 128'h1 << _EVAL_1408;
  assign _EVAL_583 = _EVAL_473 & _EVAL_826;
  assign gateways_gateway_116__EVAL_0 = _EVAL_9;
  assign _EVAL_673 = _EVAL_1697 ? _EVAL_826 : _EVAL_1537;
  assign _EVAL_1308 = _EVAL_195 & _EVAL_3696;
  assign _EVAL_1220 = _EVAL_3538 & _EVAL_826;
  assign _EVAL_2264 = _EVAL_3349[4];
  assign gateways_gateway_60__EVAL_0 = _EVAL_9;
  assign gateways_gateway_84__EVAL_0 = _EVAL_9;
  assign fanin__EVAL_57 = _EVAL_3437;
  assign _EVAL_1631 = _EVAL_1433 ? _EVAL_826 : _EVAL_3560;
  assign _EVAL_3804 = _EVAL_2144 & _EVAL_826;
  assign _EVAL_939 = _EVAL_1158 & _EVAL_826;
  assign _EVAL_3335 = _EVAL_1418 ? {{29'd0}, _EVAL_2281} : _EVAL_2838;
  assign _EVAL_3326 = _EVAL_446 ? _EVAL_826 : _EVAL_1637;
  assign _EVAL_3612 = _EVAL_195 & _EVAL_560;
  assign _EVAL_1333 = _EVAL_195 & _EVAL_3622;
  assign _EVAL_2720 = _EVAL_3204 ? _EVAL_826 : _EVAL_2533;
  assign _EVAL_3760 = _EVAL_3349[98];
  assign _EVAL_2282 = _EVAL_3349[59];
  assign _EVAL_2555 = _EVAL_3797 & _EVAL_826;
  assign _EVAL_3343 = _EVAL_651[88];
  assign _EVAL_796 = _EVAL_3804 & _EVAL_2035;
  assign _EVAL_3488 = _EVAL_3153 ? _EVAL_826 : _EVAL_3723;
  assign _EVAL_3089 = _EVAL_195 & _EVAL_1135;
  assign _EVAL_2906 = _EVAL_651[117];
  assign _EVAL_609 = ~_EVAL_1618;
  assign gateways_gateway_16__EVAL_0 = _EVAL_9;
  assign _EVAL_987 = 10'h2c == _EVAL_2998;
  assign fanin__EVAL_73 = _EVAL_3080;
  assign _EVAL_3849 = _EVAL_3349[30];
  assign _EVAL_3341 = _EVAL_3349[51];
  assign _EVAL_2345 = _EVAL_2503 | gateways_gateway_31__EVAL_4;
  assign _EVAL_1902 = 10'h4c == _EVAL_2998;
  assign _EVAL_1008 = _EVAL_3047 ? {{29'd0}, _EVAL_2575} : _EVAL_434;
  assign gateways_gateway_78__EVAL_1 = ~_EVAL_3199;
  assign gateways_gateway_26__EVAL = _EVAL_100;
  assign _EVAL_150 = _EVAL_1697 ? {{29'd0}, _EVAL_3798} : _EVAL_2171;
  assign fanin__EVAL_127 = _EVAL_2621;
  assign _EVAL_2624 = _EVAL_651[103];
  assign _EVAL_1395 = _EVAL_1857 ? {{29'd0}, _EVAL_1758} : _EVAL_3404;
  assign _EVAL_334 = _EVAL_164 ? _EVAL_826 : _EVAL_1472;
  assign gateways_gateway_33__EVAL = _EVAL;
  assign _EVAL_214 = _EVAL_3725 & _EVAL_826;
  assign _EVAL_1251 = _EVAL_776 & _EVAL_826;
  assign gateways_gateway_121__EVAL_3 = _EVAL_110;
  assign gateways_gateway_80__EVAL_0 = _EVAL_9;
  assign _EVAL_2055 = _EVAL_1592 & _EVAL_826;
  assign gateways_gateway_43__EVAL_0 = _EVAL_9;
  assign _EVAL_3222 = {_EVAL_1138,_EVAL_3527,_EVAL_3145,_EVAL_1368,_EVAL_677,_EVAL_2668,_EVAL_193,_EVAL_3112};
  assign _EVAL_2872 = _EVAL_2080 ? {{29'd0}, _EVAL_2982} : _EVAL_683;
  assign _EVAL_2103 = _EVAL_651[85];
  assign _EVAL_3475 = {_EVAL_2344,_EVAL_2685,_EVAL_3151,_EVAL_276,_EVAL_594,_EVAL_1774,_EVAL_3643};
  assign _EVAL_1871 = _EVAL_2274 ? {{29'd0}, _EVAL_189} : _EVAL_2230;
  assign _EVAL_3337 = 10'h66 == _EVAL_2998;
  assign _EVAL_1512 = _EVAL_3349[2];
  assign gateways_gateway_45__EVAL_0 = _EVAL_9;
  assign fanin__EVAL_38 = _EVAL_3218;
  assign _EVAL_3483 = _EVAL_2298 | gateways_gateway_101__EVAL_4;
  assign gateways_gateway_104__EVAL_3 = _EVAL_110;
  assign _EVAL_1292 = _EVAL_3349[83];
  assign _EVAL_2989 = _EVAL_195 & _EVAL_3619;
  assign gateways_gateway_106__EVAL_2 = _EVAL_2917[107];
  assign _EVAL_3266 = &_EVAL_3038;
  assign fanin__EVAL_16 = _EVAL_1621;
  assign gateways_gateway_44__EVAL_3 = _EVAL_110;
  assign _EVAL_184 = _EVAL_651[64];
  assign gateways_gateway_67__EVAL = _EVAL_48;
  assign _EVAL_2148 = _EVAL_1187 | gateways_gateway_93__EVAL_4;
  assign gateways_gateway_29__EVAL_3 = _EVAL_110;
  assign _EVAL_3347 = _EVAL_3328 & _EVAL_3266;
  assign _EVAL_3519 = _EVAL_232 & _EVAL_2035;
  assign _EVAL_908 = _EVAL_1739 & _EVAL_2035;
  assign fanin__EVAL_70 = _EVAL_240;
  assign _EVAL_3391 = 10'h2d == _EVAL_2998;
  assign _EVAL_2628 = _EVAL_2974 ? {{29'd0}, _EVAL_1341} : _EVAL_2451;
  assign _EVAL_3259 = _EVAL_3566 ? _EVAL_826 : _EVAL_1254;
  assign _EVAL_1994 = {_EVAL_3199,_EVAL_1524,_EVAL_2153,_EVAL_2900,_EVAL_744,_EVAL_2682,_EVAL_2719,_EVAL_2509,_EVAL_2520
    };
  assign _EVAL_2320 = _EVAL_3349[88];
  assign _EVAL_3193 = _EVAL_573 ? _EVAL_826 : _EVAL_3069;
  assign gateways_gateway_86__EVAL = _EVAL_24;
  assign _EVAL_1472 = _EVAL_3504 ? _EVAL_826 : _EVAL_3534;
  assign _EVAL_3007 = _EVAL_3275 & _EVAL_826;
  assign gateways_gateway_125__EVAL = _EVAL_41;
  assign gateways_gateway_14__EVAL = _EVAL_55;
  assign gateways_gateway_41__EVAL_1 = ~_EVAL_902;
  assign _EVAL_2800 = _EVAL_695 ? {{29'd0}, _EVAL_2580} : _EVAL_2938;
  assign _EVAL_2034 = _EVAL_584 ? {{29'd0}, _EVAL_2621} : _EVAL_3454;
  assign _EVAL_422 = _EVAL_195 & _EVAL_2906;
  assign gateways_gateway_6__EVAL = _EVAL_137;
  assign _EVAL_625 = _EVAL_651[53];
  assign gateways_gateway_57__EVAL_2 = _EVAL_2917[58];
  assign _EVAL_2035 = &_EVAL_2084;
  assign gateways_gateway_118__EVAL_2 = _EVAL_2917[119];
  assign fanin__EVAL_0 = _EVAL_1968;
  assign gateways_gateway_31__EVAL_0 = _EVAL_9;
  assign _EVAL_1182 = _EVAL_471 | gateways_gateway_7__EVAL_4;
  assign _EVAL_593 = _EVAL_3237 & _EVAL_826;
  assign fanin__EVAL_76 = _EVAL_2637;
  assign _EVAL_1195 = _EVAL_362 | gateways_gateway_68__EVAL_4;
  assign _EVAL_1489 = ~_EVAL_1190;
  assign gateways_gateway_113__EVAL_2 = _EVAL_2917[114];
  assign gateways_gateway_52__EVAL_3 = _EVAL_110;
  assign gateways_gateway_80__EVAL_3 = _EVAL_110;
  assign _EVAL_3545 = _EVAL_3349[87];
  assign gateways_gateway_56__EVAL_1 = ~_EVAL_423;
  assign _EVAL_3426 = _EVAL_3349[43];
  assign _EVAL_2515 = _EVAL_209 & _EVAL_826;
  assign gateways_gateway_42__EVAL_3 = _EVAL_110;
  assign _EVAL_257 = _EVAL_3349[86];
  assign gateways_gateway_78__EVAL_0 = _EVAL_9;
  assign _EVAL_495 = ~_EVAL_3381;
  assign gateways_gateway_62__EVAL_2 = _EVAL_2917[63];
  assign _EVAL_408 = 10'h61 == _EVAL_2998;
  assign _EVAL_3463 = 10'h67 == _EVAL_2998;
  assign fanin__EVAL_99 = _EVAL_189;
  assign _EVAL_3179 = _EVAL_2149 & _EVAL_2035;
  assign gateways_gateway_50__EVAL_1 = ~_EVAL_819;
  assign _EVAL_1480 = _EVAL_3349[123];
  assign _EVAL_2649 = _EVAL_2196 | gateways_gateway_53__EVAL_4;
  assign fanin__EVAL_91 = _EVAL_3446;
  assign _EVAL_2155 = _EVAL_1343 & _EVAL_826;
  assign _EVAL_1264 = _EVAL_3349[61];
  assign gateways_gateway_106__EVAL_0 = _EVAL_9;
  assign _EVAL_683 = _EVAL_2397 ? {{29'd0}, _EVAL_167} : _EVAL_524;
  assign _EVAL_19 = _EVAL_809 > _EVAL_3156;
  assign _EVAL_3696 = _EVAL_651[10];
  assign _EVAL_2865 = _EVAL_651[7];
  assign _EVAL_2206 = _EVAL_1677 & _EVAL_2035;
  assign _EVAL_1057 = _EVAL_651[100];
  assign _EVAL_614 = _EVAL_1203 & _EVAL_826;
  assign _EVAL_463 = _EVAL_651[63];
  assign _EVAL_1677 = _EVAL_2252 & _EVAL_826;
  assign _EVAL_1096 = 10'h7b == _EVAL_2998;
  assign _EVAL_1853 = _EVAL_1033 | gateways_gateway_125__EVAL_4;
  assign gateways_gateway_9__EVAL_0 = _EVAL_9;
  assign _EVAL_1066 = _EVAL_651[69];
  assign _EVAL_1579 = _EVAL_3340 & _EVAL_826;
  assign gateways_gateway_101__EVAL_1 = ~_EVAL_2160;
  assign fanin__EVAL_48 = _EVAL_2296 & _EVAL_304;
  assign _EVAL_2710 = _EVAL_3123 ? _EVAL_826 : 1'h1;
  assign _EVAL_2216 = _EVAL_3349[55];
  assign _EVAL_3134 = _EVAL_3819 ? {{29'd0}, _EVAL_1796} : _EVAL_2650;
  assign _EVAL_2520 = {_EVAL_1365,_EVAL_2737,_EVAL_811,_EVAL_3440,_EVAL_3387,_EVAL_3305,_EVAL_770,_EVAL_526};
  assign _EVAL_3201 = 10'h64 == _EVAL_2998;
  assign _EVAL_944 = ~_EVAL_3122;
  assign fanin__EVAL_13 = _EVAL_3055;
  assign _EVAL_2061 = _EVAL_1912 ? _EVAL_826 : _EVAL_411;
  assign gateways_gateway_60__EVAL_1 = ~_EVAL_350;
  assign _EVAL_1320 = _EVAL_1238 & _EVAL_2035;
  assign _EVAL_3531 = _EVAL_1751 | gateways_gateway_100__EVAL_4;
  assign _EVAL_1257 = ~_EVAL_1346;
  assign _EVAL_2486 = _EVAL_3402 ? {{29'd0}, _EVAL_2079} : _EVAL_2969;
  assign _EVAL_369 = _EVAL_651[94];
  assign _EVAL_3595 = ~_EVAL_1140;
  assign gateways_gateway_109__EVAL_0 = _EVAL_9;
  assign _EVAL_1224 = _EVAL_195 & _EVAL_515;
  assign gateways_gateway_90__EVAL_2 = _EVAL_2917[91];
  assign _EVAL_126 = out_back__EVAL_6;
  assign gateways_gateway_49__EVAL_0 = _EVAL_9;
  assign gateways_gateway_124__EVAL_0 = _EVAL_9;
  assign _EVAL_1051 = _EVAL_3161 & _EVAL_2035;
  assign _EVAL_2632 = _EVAL_860 ? _EVAL_826 : _EVAL_3209;
  assign gateways_gateway_47__EVAL_0 = _EVAL_9;
  assign gateways_gateway_67__EVAL_0 = _EVAL_9;
  assign _EVAL_124 = out_back__EVAL_11;
  assign _EVAL_3777 = _EVAL_3392 | gateways_gateway_22__EVAL_4;
  assign fanin__EVAL_115 = _EVAL_1687;
  assign _EVAL_2589 = _EVAL_1096 ? _EVAL_826 : _EVAL_1935;
  assign _EVAL_2739 = _EVAL_3399 & _EVAL_826;
  assign _EVAL_735 = _EVAL_3349[70];
  assign _EVAL_1033 = _EVAL_3349[126];
  assign gateways_gateway_48__EVAL_2 = _EVAL_2917[49];
  assign gateways_gateway_96__EVAL_0 = _EVAL_9;
  assign _EVAL_2777 = _EVAL_3811 | gateways_gateway_18__EVAL_4;
  assign _EVAL_3401 = _EVAL_225 ? _EVAL_826 : _EVAL_3193;
  assign gateways_gateway_93__EVAL = _EVAL_128;
  assign fanin__EVAL_37 = _EVAL_3216;
  assign _EVAL_2028 = ~_EVAL_2503;
  assign gateways_gateway_121__EVAL = _EVAL_112;
  assign gateways_gateway_12__EVAL_2 = _EVAL_2917[13];
  assign gateways_gateway_100__EVAL = _EVAL_77;
  assign gateways_gateway_90__EVAL = _EVAL_2;
  assign _EVAL_3486 = _EVAL_2860 | gateways_gateway_33__EVAL_4;
  assign gateways_gateway_35__EVAL_1 = ~_EVAL_1368;
  assign _EVAL_842 = _EVAL_3349[5];
  assign _EVAL_1011 = _EVAL_3349[120];
  assign _EVAL_838 = _EVAL_651[47];
  assign gateways_gateway_32__EVAL_2 = _EVAL_2917[33];
  assign _EVAL_2150 = _EVAL_378 & _EVAL_826;
  assign _EVAL_2196 = _EVAL_3349[54];
  assign gateways_gateway_6__EVAL_1 = ~_EVAL_2344;
  assign _EVAL_1081 = _EVAL_1333 & _EVAL_826;
  assign fanin__EVAL_3 = _EVAL_3744;
  assign _EVAL_1288 = _EVAL_166 ? _EVAL_826 : _EVAL_2934;
  assign gateways_gateway_5__EVAL_0 = _EVAL_9;
  assign _EVAL_2380 = _EVAL_2222 | gateways_gateway_25__EVAL_4;
  assign gateways_gateway_7__EVAL_2 = _EVAL_2917[8];
  assign _EVAL_1670 = 10'h21 == _EVAL_2998;
  assign gateways_gateway_90__EVAL_1 = ~_EVAL_3627;
  assign _EVAL_1026 = 10'h22 == _EVAL_2998;
  assign gateways_gateway_101__EVAL = _EVAL_142;
  assign _EVAL_245 = _EVAL_195 & _EVAL_2484;
  assign _EVAL_2312 = _EVAL_595 ? _EVAL_826 : _EVAL_3620;
  assign _EVAL_1254 = _EVAL_179 ? _EVAL_826 : _EVAL_2965;
  assign _EVAL_989 = _EVAL_1618 | gateways_gateway_11__EVAL_4;
  assign _EVAL_492 = _EVAL_281 ? {{29'd0}, _EVAL_854} : _EVAL_3455;
  assign _EVAL_2556 = _EVAL_1122 | gateways_gateway_28__EVAL_4;
  assign _EVAL_2406 = _EVAL_651[101];
  assign _EVAL_2812 = _EVAL_3349[124];
  assign _EVAL_1793 = _EVAL_651[38];
  assign _EVAL_3278 = _EVAL_195 & _EVAL_1094;
  assign _EVAL_978 = _EVAL_1799 ? {{29'd0}, _EVAL_3005} : _EVAL_3335;
  assign gateways_gateway_126__EVAL_2 = _EVAL_2917[127];
  assign _EVAL_2289 = _EVAL_1762 | gateways_gateway_113__EVAL_4;
  assign gateways_gateway_5__EVAL_2 = _EVAL_2917[6];
  assign _EVAL_2251 = _EVAL_3349[125];
  assign _EVAL_471 = _EVAL_3349[8];
  assign fanin__EVAL_22 = _EVAL_2012;
  assign _EVAL_3030 = _EVAL_2342 & _EVAL_826;
  assign gateways_gateway_24__EVAL_2 = _EVAL_2917[25];
  assign _EVAL_2285 = _EVAL_504 ? {{29'd0}, _EVAL_3055} : _EVAL_3102;
  assign _EVAL_3729 = _EVAL_651[83];
  assign gateways_gateway_58__EVAL = _EVAL_104;
  assign _EVAL_3368 = _EVAL_651[52];
  assign _EVAL_3324 = ~_EVAL_1187;
  assign _EVAL_1415 = _EVAL_2881 ? {{29'd0}, _EVAL_1283} : _EVAL_2205;
  assign _EVAL_531 = _EVAL_468 & _EVAL_826;
  assign _EVAL_741 = _EVAL_2155 & _EVAL_1700;
  assign _EVAL_2482 = _EVAL_3349[46];
  assign _EVAL_2062 = _EVAL_1274 ? {{29'd0}, _EVAL_240} : _EVAL_3134;
  assign _EVAL_1281 = _EVAL_236 & _EVAL_826;
  assign gateways_gateway_79__EVAL_1 = ~_EVAL_2221;
  assign _EVAL_3036 = _EVAL_651[3];
  assign _EVAL_1828 = _EVAL_3349[105];
  assign _EVAL_2676 = _EVAL_195 & _EVAL_2152;
  assign _EVAL_1907 = ~_EVAL_3378;
  assign _EVAL_2914 = _EVAL_2850[31:24];
  assign _EVAL_2224 = _EVAL_651[4];
  assign _EVAL_3319 = _EVAL_651[15];
  assign _EVAL_899 = _EVAL_2907 | gateways_gateway_114__EVAL_4;
  assign _EVAL_1768 = _EVAL_195 & _EVAL_3319;
  assign _EVAL_1867 = 10'h6d == _EVAL_2998;
  assign _EVAL_652 = _EVAL_3802 & _EVAL_2035;
  assign gateways_gateway_104__EVAL = _EVAL_82;
  assign _EVAL_3481 = 10'h59 == _EVAL_2998;
  assign _EVAL_2479 = _EVAL_482 | gateways_gateway_44__EVAL_4;
  assign gateways_gateway_68__EVAL_3 = _EVAL_110;
  assign _EVAL_3797 = _EVAL_195 & _EVAL_2733;
  assign _EVAL_3261 = _EVAL_1264 | gateways_gateway_60__EVAL_4;
  assign _EVAL_2218 = _EVAL_2817 & _EVAL_826;
  assign _EVAL_3399 = _EVAL_195 & _EVAL_2406;
  assign gateways_gateway_36__EVAL_1 = ~_EVAL_3145;
  assign gateways_gateway_54__EVAL = _EVAL_56;
  assign gateways_gateway_10__EVAL = _EVAL_138;
  assign _EVAL_3718 = _EVAL_2619 & _EVAL_826;
  assign _EVAL_1209 = _EVAL_646 | gateways_gateway_2__EVAL_4;
  assign _EVAL_3316 = ~_EVAL_1292;
  assign _EVAL_776 = _EVAL_195 & _EVAL_903;
  assign _EVAL_2619 = _EVAL_195 & _EVAL_1090;
  assign _EVAL_1021 = _EVAL_195 & _EVAL_3456;
  assign _EVAL_3285 = ~_EVAL_904;
  assign _EVAL_1666 = 10'h83 == _EVAL_2998;
  assign _EVAL_1549 = ~_EVAL_2099;
  assign _EVAL_3390 = _EVAL_3071 & _EVAL_2035;
  assign gateways_gateway_116__EVAL_1 = ~_EVAL_1948;
  assign gateways_gateway_124__EVAL_1 = ~_EVAL_1417;
  assign _EVAL_536 = _EVAL_2653 & _EVAL_826;
  assign _EVAL_2559 = _EVAL_3480 & _EVAL_826;
  assign gateways_gateway_33__EVAL_2 = _EVAL_2917[34];
  assign _EVAL_296 = ~_EVAL_2607;
  assign _EVAL_765 = _EVAL_3030 & _EVAL_644;
  assign _EVAL_3204 = 10'h6e == _EVAL_2998;
  assign _EVAL_1857 = 10'hd == _EVAL_2998;
  assign _EVAL_2011 = _EVAL_2702 & _EVAL_2035;
  assign _EVAL_3243 = _EVAL_651[60];
  assign gateways_gateway_12__EVAL_3 = _EVAL_110;
  assign _EVAL_3720 = _EVAL_382 & _EVAL_2035;
  assign _EVAL_709 = _EVAL_651[104];
  assign gateways_gateway_65__EVAL_2 = _EVAL_2917[66];
  assign _EVAL_1171 = 10'h81 == _EVAL_2998;
  assign gateways_gateway_51__EVAL_3 = _EVAL_110;
  assign gateways_gateway_114__EVAL = _EVAL_12;
  assign _EVAL_2195 = _EVAL_1722 & _EVAL_826;
  assign gateways_gateway_43__EVAL_2 = _EVAL_2917[44];
  assign _EVAL_2392 = _EVAL_2558 | gateways_gateway_126__EVAL_4;
  assign gateways_gateway_17__EVAL = _EVAL_10;
  assign gateways_gateway_79__EVAL_3 = _EVAL_110;
  assign _EVAL_810 = out_back__EVAL_1[2:0];
  assign _EVAL_3375 = _EVAL_753 | gateways_gateway_12__EVAL_4;
  assign gateways_gateway_36__EVAL_2 = _EVAL_2917[37];
  assign gateways_gateway_112__EVAL_1 = ~_EVAL_414;
  assign _EVAL_3355 = {_EVAL_1964,_EVAL_302,_EVAL_1467,_EVAL_612,_EVAL_498,_EVAL_2174,_EVAL_2165,_EVAL_911};
  assign gateways_gateway_39__EVAL_1 = ~_EVAL_1576;
  assign _EVAL_849 = 10'h6 == _EVAL_2998;
  assign gateways_gateway_102__EVAL_0 = _EVAL_9;
  assign gateways_gateway_56__EVAL_2 = _EVAL_2917[57];
  assign gateways_gateway_27__EVAL = _EVAL_25;
  assign _EVAL_236 = _EVAL_195 & _EVAL_1763;
  assign _EVAL_2053 = _EVAL_1920 ? _EVAL_826 : _EVAL_1627;
  assign _EVAL_2060 = _EVAL_1987 ? {{29'd0}, _EVAL_1293} : _EVAL_3706;
  assign gateways_gateway_75__EVAL_2 = _EVAL_2917[76];
  assign gateways_gateway_18__EVAL_3 = _EVAL_110;
  assign _EVAL_1153 = _EVAL_1826 | gateways_gateway_36__EVAL_4;
  assign _EVAL_282 = _EVAL_301 & _EVAL_826;
  assign _EVAL_815 = _EVAL_2349 ? {{29'd0}, _EVAL_1252} : _EVAL_2800;
  assign _EVAL_2450 = {_EVAL_1847,_EVAL_1434,_EVAL_1347,_EVAL_2961,_EVAL_2143,_EVAL_3268,_EVAL_2370,_EVAL_3129,
    _EVAL_3355,_EVAL_2889};
  assign _EVAL_244 = _EVAL_2852 & _EVAL_2035;
  assign _EVAL_855 = _EVAL_3271 | gateways_gateway_17__EVAL_4;
  assign _EVAL_3845 = _EVAL_3246 | gateways_gateway_63__EVAL_4;
  assign gateways_gateway_47__EVAL_1 = ~_EVAL_3059;
  assign out_back__EVAL_5 = _EVAL_84;
  assign _EVAL_1564 = _EVAL_916 | gateways_gateway_121__EVAL_4;
  assign gateways_gateway_69__EVAL_1 = ~_EVAL_2737;
  assign _EVAL_2970 = 10'h68 == _EVAL_2998;
  assign _EVAL_2956 = 10'h3e == _EVAL_2998;
  assign _EVAL_1408 = _EVAL_2175[6:0];
  assign fanin__EVAL_25 = _EVAL_1805;
  assign gateways_gateway_53__EVAL_3 = _EVAL_110;
  assign _EVAL_3695 = _EVAL_3074 ? _EVAL_826 : _EVAL_2784;
  assign gateways_gateway_65__EVAL_1 = ~_EVAL_3305;
  assign gateways_gateway_74__EVAL_1 = ~_EVAL_744;
  assign gateways_gateway_119__EVAL_0 = _EVAL_9;
  assign _EVAL_2190 = _EVAL_988 & _EVAL_2035;
  assign _EVAL_219 = _EVAL_1140 | gateways_gateway_52__EVAL_4;
  assign _EVAL_3138 = _EVAL_3349[93];
  assign gateways_gateway_62__EVAL_3 = _EVAL_110;
  assign _EVAL_576 = {_EVAL_3770,_EVAL_1576,_EVAL_1138,_EVAL_3527,_EVAL_3145,_EVAL_1368,_EVAL_677,_EVAL_2668,_EVAL_193,
    _EVAL_3112};
  assign gateways_gateway_82__EVAL_3 = _EVAL_110;
  assign gateways_gateway_14__EVAL_0 = _EVAL_9;
  assign _EVAL_2408 = 10'h69 == _EVAL_2998;
  assign gateways_gateway_64__EVAL_1 = ~_EVAL_770;
  assign gateways_gateway_117__EVAL = _EVAL_83;
  assign _EVAL_2474 = _EVAL_3444 & _EVAL_826;
  assign _EVAL_2903 = {_EVAL_2655,_EVAL_668,_EVAL_2167,_EVAL_965,_EVAL_202,_EVAL_1116,_EVAL_1948,_EVAL_3803,_EVAL_2193,
    _EVAL_909};
  assign _EVAL_1812 = 10'h47 == _EVAL_2998;
  assign _EVAL_3600 = _EVAL_2617 & _EVAL_826;
  assign _EVAL_3714 = _EVAL_1923 ? {{29'd0}, _EVAL_1695} : _EVAL_894;
  assign _EVAL_1017 = 10'h63 == _EVAL_2998;
  assign _EVAL_1385 = _EVAL_1801 & _EVAL_826;
  assign _EVAL_1794 = _EVAL_3081 & _EVAL_826;
  assign _EVAL_295 = _EVAL_651[17];
  assign _EVAL_509 = _EVAL_342 & _EVAL_2035;
  assign fanin__EVAL_89 = _EVAL_2753;
  assign _EVAL_1664 = _EVAL_3127 & _EVAL_2035;
  assign gateways_gateway_8__EVAL_2 = _EVAL_2917[9];
  assign _EVAL_2314 = _EVAL_2956 ? {{29'd0}, _EVAL_2845} : _EVAL_815;
  assign _EVAL_1761 = _EVAL_195 & _EVAL_1304;
  assign _EVAL_1826 = _EVAL_3349[37];
  assign _EVAL_3039 = _EVAL_3349[44];
  assign gateways_gateway_20__EVAL = _EVAL_122;
  assign _EVAL_1506 = 10'h5a == _EVAL_2998;
  assign gateways_gateway_30__EVAL_2 = _EVAL_2917[31];
  assign gateways_gateway_28__EVAL = _EVAL_43;
  assign gateways_gateway_23__EVAL = _EVAL_40;
  assign _EVAL_1792 = ~_EVAL_1764;
  assign gateways_gateway_12__EVAL = _EVAL_54;
  assign _EVAL_3848 = _EVAL_2557 ? {{29'd0}, _EVAL_797} : _EVAL_957;
  assign _EVAL_179 = 10'h6c == _EVAL_2998;
  assign _EVAL_2689 = _EVAL_3111 & _EVAL_2035;
  assign _EVAL_1325 = _EVAL_3529 & _EVAL_826;
  assign _EVAL_3616 = _EVAL_195 & _EVAL_838;
  assign gateways_gateway_43__EVAL = _EVAL_69;
  assign _EVAL_533 = _EVAL_2389 & _EVAL_2035;
  assign _EVAL_2088 = out_back__EVAL_7 & _EVAL_136;
  assign gateways_gateway_20__EVAL_0 = _EVAL_9;
  assign _EVAL_2077 = _EVAL_3349[106];
  assign _EVAL_2842 = _EVAL_195 & _EVAL_3747;
  assign gateways_gateway_80__EVAL = _EVAL_95;
  assign gateways_gateway_108__EVAL_2 = _EVAL_2917[109];
  assign gateways_gateway_123__EVAL_1 = ~_EVAL_2178;
  assign _EVAL_645 = _EVAL_3251 ? _EVAL_826 : _EVAL_3361;
  assign gateways_gateway_122__EVAL_1 = ~_EVAL_2655;
  assign gateways_gateway_125__EVAL_1 = ~_EVAL_1147;
  assign _EVAL_1678 = _EVAL_3270 ? {{29'd0}, _EVAL_3835} : _EVAL_366;
  assign _EVAL_655 = _EVAL_3349[100];
  assign _EVAL_466 = _EVAL_1828 | gateways_gateway_104__EVAL_4;
  assign _EVAL_2386 = _EVAL_1026 ? {{29'd0}, _EVAL_3216} : _EVAL_1623;
  assign _EVAL_1780 = _EVAL_651[93];
  assign gateways_gateway_65__EVAL = _EVAL_134;
  assign gateways_gateway_33__EVAL_3 = _EVAL_110;
  assign gateways_gateway_102__EVAL_2 = _EVAL_2917[103];
  assign gateways_gateway_10__EVAL_1 = ~_EVAL_3140;
  assign gateways_gateway_17__EVAL_1 = ~_EVAL_2174;
  assign _EVAL_2204 = _EVAL_488 ? {{29'd0}, _EVAL_2186} : _EVAL_2095;
  assign gateways_gateway_84__EVAL_1 = ~_EVAL_1937;
  assign _EVAL_1769 = _EVAL_3030 & _EVAL_425;
  assign _EVAL_1140 = _EVAL_3349[53];
  assign fanin__EVAL_60 = _EVAL_865;
  assign _EVAL_1315 = _EVAL_3123 ? _EVAL_2639 : 32'h0;
  assign gateways_gateway_112__EVAL_3 = _EVAL_110;
  assign _EVAL_3471 = _EVAL_1912 ? {{29'd0}, _EVAL_2466} : _EVAL_3680;
  assign _EVAL_1413 = _EVAL_3349[11];
  assign gateways_gateway_92__EVAL_2 = _EVAL_2917[93];
  assign _EVAL_1568 = _EVAL_856 ? {{29'd0}, _EVAL_953} : _EVAL_1167;
  assign _EVAL_1751 = _EVAL_3349[101];
  assign gateways_gateway_114__EVAL_2 = _EVAL_2917[115];
  assign _EVAL_752 = _EVAL_488 ? _EVAL_826 : _EVAL_850;
  assign _EVAL_2300 = _EVAL_2561 ? _EVAL_3336 : _EVAL_3076;
  assign gateways_gateway_110__EVAL = _EVAL_135;
  assign _EVAL_2377 = {_EVAL_1471,_EVAL_2070,_EVAL_2418,_EVAL_1517,_EVAL_1340,_EVAL_1380,_EVAL_394,_EVAL_2877,_EVAL_2902
    ,1'h0};
  assign _EVAL_458 = _EVAL_1243 | gateways_gateway_94__EVAL_4;
  assign _EVAL_2871 = _EVAL_3463 ? {{29'd0}, _EVAL_2873} : _EVAL_1779;
  assign _EVAL_988 = _EVAL_1610 & _EVAL_826;
  assign _EVAL_1593 = _EVAL_408 ? _EVAL_826 : _EVAL_1307;
  assign gateways_gateway_42__EVAL_2 = _EVAL_2917[43];
  assign _EVAL_1550 = out_back__EVAL_3[3];
  assign gateways_gateway_61__EVAL_0 = _EVAL_9;
  assign fanin__EVAL_87 = _EVAL_3469;
  assign _EVAL_3435 = _EVAL_651[80];
  assign _EVAL_341 = _EVAL_3349[65];
  assign _EVAL_1764 = _EVAL_3349[41];
  assign _EVAL_967 = _EVAL_1480 | gateways_gateway_122__EVAL_4;
  assign gateways_gateway_28__EVAL_0 = _EVAL_9;
  assign _EVAL_2417 = _EVAL_451 ? _EVAL_826 : _EVAL_3815;
  assign gateways_gateway_123__EVAL_0 = _EVAL_9;
  assign gateways_gateway_31__EVAL_2 = _EVAL_2917[32];
  assign _EVAL_1674 = ~_EVAL_2415;
  assign _EVAL_3510 = _EVAL_374 ? _EVAL_826 : _EVAL_2303;
  assign _EVAL_382 = _EVAL_2473 & _EVAL_826;
  assign _EVAL_2730 = _EVAL_3174 | gateways_gateway_91__EVAL_4;
  assign _EVAL_365 = _EVAL_651[123];
  assign gateways_gateway_120__EVAL_2 = _EVAL_2917[121];
  assign _EVAL_667 = _EVAL_956 & _EVAL_826;
  assign gateways_gateway_122__EVAL_3 = _EVAL_110;
  assign _EVAL_1307 = _EVAL_2844 ? _EVAL_826 : _EVAL_3567;
  assign _EVAL_1382 = _EVAL_2341 | gateways_gateway_26__EVAL_4;
  assign _EVAL_1241 = _EVAL_408 ? {{29'd0}, _EVAL_3096} : _EVAL_2275;
  assign _EVAL_758 = _EVAL_3819 ? _EVAL_826 : _EVAL_3569;
  assign _EVAL_1623 = _EVAL_1879 ? {{29'd0}, _EVAL_3635} : _EVAL_2285;
  assign _EVAL_2234 = _EVAL_651[97];
  assign _EVAL_1866 = {_EVAL_1369,_EVAL_3508,_EVAL_423,_EVAL_2502,_EVAL_3346,_EVAL_3150,_EVAL_1749,_EVAL_3014,_EVAL_819,
    _EVAL_982};
  assign gateways_gateway_96__EVAL = _EVAL_120;
  assign _EVAL_1722 = _EVAL_195 & _EVAL_1877;
  assign gateways_gateway_93__EVAL_0 = _EVAL_9;
  assign gateways_gateway_92__EVAL_3 = _EVAL_110;
  assign _EVAL_2399 = ~_EVAL_1043;
  assign fanin__EVAL_92 = _EVAL_3734;
  assign gateways_gateway_22__EVAL_3 = _EVAL_110;
  assign _EVAL_1304 = _EVAL_651[257];
  assign gateways_gateway_83__EVAL_1 = ~_EVAL_1270;
  assign _EVAL_627 = _EVAL_1765 & _EVAL_826;
  assign _EVAL_646 = _EVAL_3349[3];
  assign _EVAL_2095 = _EVAL_299 ? {{29'd0}, _EVAL_3559} : _EVAL_1496;
  assign _EVAL_2527 = _EVAL_3349[10];
  assign _EVAL_344 = _EVAL_1542 | gateways_gateway_32__EVAL_4;
  assign gateways_gateway_30__EVAL_1 = ~_EVAL_1847;
  assign _EVAL_3794 = ~_EVAL_1542;
  assign _EVAL_1483 = _EVAL_2842 & _EVAL_826;
  assign _EVAL_2379 = out_back__EVAL_1[23:16];
  assign _EVAL_955 = 10'h37 == _EVAL_2998;
  assign _EVAL_3663 = ~_EVAL_964;
  assign _EVAL_3828 = 10'h31 == _EVAL_2998;
  assign fanin__EVAL_40 = _EVAL_3737;
  assign gateways_gateway_116__EVAL_3 = _EVAL_110;
  assign gateways_gateway_122__EVAL_2 = _EVAL_2917[123];
  assign fanin__EVAL_96 = _EVAL_936;
  assign gateways_gateway_94__EVAL = _EVAL_30;
  assign _EVAL_1788 = _EVAL_421 & _EVAL_826;
  assign _EVAL_2928 = _EVAL_341 | gateways_gateway_64__EVAL_4;
  assign gateways_gateway_42__EVAL_1 = ~_EVAL_2268;
  assign gateways_gateway_101__EVAL_3 = _EVAL_110;
  assign _EVAL_3533 = 10'h1d == _EVAL_2998;
  assign gateways_gateway_20__EVAL_3 = _EVAL_110;
  assign gateways_gateway_111__EVAL_0 = _EVAL_9;
  assign gateways_gateway_56__EVAL_3 = _EVAL_110;
  assign gateways_gateway_97__EVAL_1 = ~_EVAL_325;
  assign gateways_gateway_118__EVAL = _EVAL_45;
  assign gateways_gateway_34__EVAL_1 = ~_EVAL_677;
  assign _EVAL_1661 = _EVAL_451 ? {{29'd0}, _EVAL_628} : _EVAL_2199;
  assign _EVAL_3270 = 10'h54 == _EVAL_2998;
  assign _EVAL_3622 = _EVAL_651[16];
  assign _EVAL_3329 = 10'h3d == _EVAL_2998;
  assign _EVAL_1900 = _EVAL_195 & _EVAL_3133;
  assign _EVAL_3444 = _EVAL_195 & _EVAL_2747;
  assign _EVAL_1649 = _EVAL_2088 & out_back__EVAL;
  assign _EVAL_3791 = ~_EVAL_2772;
  assign _EVAL_1482 = 10'h70 == _EVAL_2998;
  assign _EVAL_32 = {{2'd0}, _EVAL_367};
  assign fanin__EVAL_27 = _EVAL_1988;
  assign _EVAL_697 = _EVAL_651[40];
  assign gateways_gateway_101__EVAL_0 = _EVAL_9;
  assign _EVAL_468 = _EVAL_195 & _EVAL_3732;
  assign _EVAL_160 = _EVAL_651[35];
  assign gateways_gateway_66__EVAL_3 = _EVAL_110;
  assign _EVAL_2974 = 10'h9 == _EVAL_2998;
  assign _EVAL_478 = _EVAL_3299 ? {{29'd0}, _EVAL_172} : _EVAL_1854;
  assign gateways_gateway_50__EVAL_0 = _EVAL_9;
  assign _EVAL_1962 = _EVAL_1516 ? _EVAL_826 : _EVAL_1488;
  assign _EVAL_3811 = _EVAL_3349[19];
  assign _EVAL_3245 = out_back__EVAL_1[31:24];
  assign _EVAL_3210 = ~_EVAL_1826;
  assign _EVAL_1190 = _EVAL_3349[22];
  assign _EVAL_837 = _EVAL_3449 & _EVAL_2035;
  assign _EVAL_1918 = 10'h8 == _EVAL_2998;
  assign fanin__EVAL_81 = _EVAL_1407;
  assign _EVAL_3462 = _EVAL_651[39];
  assign _EVAL_2294 = ~_EVAL_496;
  assign _EVAL_1280 = _EVAL_651[92];
  assign _EVAL_963 = _EVAL_3349[15];
  assign _EVAL_300 = _EVAL_3318 & _EVAL_2035;
  assign _EVAL_1644 = _EVAL_651[8];
  assign gateways_gateway_3__EVAL_0 = _EVAL_9;
  assign gateways_gateway_92__EVAL_1 = ~_EVAL_2951;
  assign gateways_gateway_103__EVAL_2 = _EVAL_2917[104];
  assign _EVAL_2756 = _EVAL_1398 & _EVAL_2035;
  assign gateways_gateway_32__EVAL_1 = ~_EVAL_193;
  assign gateways_gateway_125__EVAL_2 = _EVAL_2917[126];
  assign _EVAL_3434 = 10'h36 == _EVAL_2998;
  assign _EVAL_3303 = ~_EVAL_257;
  assign _EVAL_2349 = 10'h3f == _EVAL_2998;
  assign _EVAL_670 = _EVAL_195 & _EVAL_3572;
  assign gateways_gateway_79__EVAL_0 = _EVAL_9;
  assign gateways_gateway_96__EVAL_2 = _EVAL_2917[97];
  assign _EVAL_1090 = _EVAL_651[126];
  assign _EVAL_638 = 10'h4b == _EVAL_2998;
  assign _EVAL_2511 = _EVAL_2922 & _EVAL_2035;
  assign _EVAL_2253 = ~_EVAL_2322;
  assign gateways_gateway_107__EVAL_2 = _EVAL_2917[108];
  assign _EVAL_2727 = _EVAL_195 & _EVAL_2633;
  assign _EVAL_3757 = _EVAL_651[75];
  assign _EVAL_3465 = _EVAL_647 ? _EVAL_826 : _EVAL_2724;
  assign gateways_gateway_31__EVAL_3 = _EVAL_110;
  assign gateways_gateway_62__EVAL = _EVAL_125;
  assign _EVAL_3646 = _EVAL_2856 & _EVAL_826;
  assign _EVAL_2558 = _EVAL_3349[127];
  assign fanin__EVAL_17 = _EVAL_3096;
  assign _EVAL_2465 = _EVAL_195 & _EVAL_1731;
  assign _EVAL_1824 = 10'h4 == _EVAL_2998;
  assign gateways_gateway_77__EVAL_2 = _EVAL_2917[78];
  assign _EVAL_267 = {_EVAL_1127,_EVAL_727,_EVAL_1937,_EVAL_1270,_EVAL_1175,_EVAL_1507,_EVAL_2297,_EVAL_2221};
  assign gateways_gateway_43__EVAL_3 = _EVAL_110;
  assign gateways_gateway_69__EVAL_0 = _EVAL_9;
  assign _EVAL_253 = _EVAL_258 | gateways_gateway_72__EVAL_4;
  assign _EVAL_3685 = ~_EVAL_3426;
  assign _EVAL_631 = _EVAL_3086 ? _EVAL_826 : _EVAL_592;
  assign _EVAL_3852 = _EVAL_651[13];
  assign _EVAL_1367 = 10'h60 == _EVAL_2998;
  assign _EVAL_1164 = _EVAL_2841 & _EVAL_2035;
  assign _EVAL_721 = _EVAL_1466 | gateways_gateway_49__EVAL_4;
  assign gateways_gateway_55__EVAL_2 = _EVAL_2917[56];
  assign gateways_gateway_40__EVAL = _EVAL_14;
  assign _EVAL_3599 = _EVAL_3349[116];
  assign gateways_gateway_64__EVAL = _EVAL_66;
  assign _EVAL_1202 = _EVAL_1518 & _EVAL_2035;
  assign _EVAL_208 = _EVAL_3481 ? _EVAL_826 : _EVAL_3579;
  assign fanin__EVAL_93 = _EVAL_1758;
  assign _EVAL_273 = _EVAL_3575 & _EVAL_826;
  assign _EVAL_1016 = _EVAL_2850[23:16];
  assign _EVAL_331 = _EVAL_1601 | gateways_gateway_46__EVAL_4;
  assign _EVAL_2604 = _EVAL_3349[99];
  assign _EVAL_1630 = _EVAL_3349[90];
  assign _EVAL_2913 = _EVAL_1630 | gateways_gateway_89__EVAL_4;
  assign gateways_gateway_41__EVAL_0 = _EVAL_9;
  assign _EVAL_3115 = _EVAL_1482 ? _EVAL_826 : _EVAL_364;
  assign _EVAL_2542 = _EVAL_3393 | gateways_gateway_19__EVAL_4;
  assign gateways_gateway_89__EVAL_2 = _EVAL_2917[90];
  assign _EVAL_1622 = _EVAL_1118 ? _EVAL_826 : _EVAL_3756;
  assign _EVAL_3311 = _EVAL_3349[104];
  assign _EVAL_1785 = _EVAL_735 | gateways_gateway_69__EVAL_4;
  assign _EVAL_3575 = _EVAL_195 & _EVAL_402;
  assign _EVAL_3807 = _EVAL_1413 | gateways_gateway_10__EVAL_4;
  assign _EVAL_3068 = _EVAL_939 & _EVAL_2035;
  assign gateways_gateway_64__EVAL_3 = _EVAL_110;
  assign gateways_gateway_115__EVAL_3 = _EVAL_110;
  assign gateways_gateway_7__EVAL_0 = _EVAL_9;
  assign _EVAL_644 = &_EVAL_3702;
  assign _EVAL_3133 = _EVAL_651[119];
  assign _EVAL_2789 = _EVAL_2019 ? {{29'd0}, _EVAL_3513} : _EVAL_1395;
  assign _EVAL_3702 = _EVAL_2850[7:1];
  assign gateways_gateway_120__EVAL_1 = ~_EVAL_2167;
  assign _EVAL_449 = _EVAL_3204 ? {{29'd0}, _EVAL_1634} : _EVAL_905;
  assign fanin__EVAL_61 = _EVAL_2845;
  assign _EVAL_959 = 10'h34 == _EVAL_2998;
  assign gateways_gateway_5__EVAL = _EVAL_37;
  assign gateways_gateway_67__EVAL_2 = _EVAL_2917[68];
  assign _EVAL_2919 = _EVAL_214 & _EVAL_2035;
  assign gateways_gateway_61__EVAL_1 = ~_EVAL_3331;
  assign gateways_gateway_91__EVAL_1 = ~_EVAL_284;
  assign gateways_gateway_95__EVAL_3 = _EVAL_110;
  assign gateways_gateway_32__EVAL = _EVAL_16;
  assign _EVAL_3271 = _EVAL_3349[18];
  assign _EVAL_156 = _EVAL_2316 | gateways_gateway_78__EVAL_4;
  assign _EVAL_2005 = _EVAL_3349[7];
  assign fanin__EVAL_63 = _EVAL_1843;
  assign fanin__EVAL_95 = _EVAL_3635;
  assign _EVAL_1366 = ~_EVAL_2005;
  assign gateways_gateway_27__EVAL_3 = _EVAL_110;
  assign _EVAL_1520 = _EVAL_3849 | gateways_gateway_29__EVAL_4;
  assign _EVAL_719 = ~_EVAL_1466;
  assign fanin__EVAL_53 = _EVAL_222;
  assign gateways_gateway_61__EVAL = _EVAL_29;
  assign _EVAL_1151 = _EVAL_195 & _EVAL_697;
  assign _EVAL_1740 = _EVAL_195 & _EVAL_416;
  assign gateways_gateway_95__EVAL = _EVAL_81;
  assign gateways_gateway_120__EVAL = _EVAL_96;
  assign gateways_gateway_115__EVAL_1 = ~_EVAL_3803;
  assign gateways_gateway_28__EVAL_1 = ~_EVAL_1347;
  assign _EVAL_2607 = _EVAL_3349[91];
  assign _EVAL_1627 = _EVAL_2561 ? _EVAL_826 : _EVAL_3401;
  assign _EVAL_2441 = _EVAL_1282 ? _EVAL_826 : _EVAL_208;
  assign gateways_gateway_51__EVAL_2 = _EVAL_2917[52];
  assign gateways_gateway_48__EVAL_3 = _EVAL_110;
  assign gateways_gateway_50__EVAL = _EVAL_106;
  assign gateways_gateway_51__EVAL_1 = ~_EVAL_3014;
  assign _EVAL_603 = ~_EVAL_1512;
  assign _EVAL_2018 = _EVAL_3801 & _EVAL_826;
  assign _EVAL_3851 = _EVAL_1184 | gateways_gateway_80__EVAL_4;
  assign _EVAL_2083 = ~_EVAL_3138;
  assign _EVAL_3321 = _EVAL_2195 & _EVAL_2035;
  assign _EVAL_1832 = _EVAL_980 | gateways_gateway_76__EVAL_4;
  assign gateways_gateway_63__EVAL_2 = _EVAL_2917[64];
  assign gateways_gateway_106__EVAL_1 = ~_EVAL_3043;
  assign _EVAL_1193 = 10'h41 == _EVAL_2998;
  assign gateways_gateway_83__EVAL_2 = _EVAL_2917[84];
  assign gateways_gateway_68__EVAL_1 = ~_EVAL_811;
  assign gateways_gateway_70__EVAL_2 = _EVAL_2917[71];
  assign _EVAL_2844 = 10'h62 == _EVAL_2998;
  assign gateways_gateway_110__EVAL_3 = _EVAL_110;
  assign _EVAL_792 = out_back__EVAL_3[5];
  assign _EVAL_933 = _EVAL_3633 | gateways_gateway_20__EVAL_4;
  assign _EVAL_428 = {_EVAL_2488,_EVAL_2160,_EVAL_2197,_EVAL_3656,_EVAL_3395,_EVAL_325,_EVAL_3200,_EVAL_415};
  assign gateways_gateway_39__EVAL = _EVAL_1;
  assign _EVAL_2696 = _EVAL_195 & _EVAL_3255;
  assign _EVAL_2254 = _EVAL_1026 ? _EVAL_826 : _EVAL_2612;
  assign gateways_gateway_4__EVAL_1 = ~_EVAL_3151;
  assign fanin__EVAL_44 = _EVAL_1527;
  assign gateways_gateway_94__EVAL_1 = ~_EVAL_2793;
  assign gateways_gateway_93__EVAL_1 = ~_EVAL_1565;
  assign _EVAL_669 = _EVAL_869 ? {{29'd0}, _EVAL_3342} : _EVAL_3591;
  assign _EVAL_2817 = _EVAL_195 & _EVAL_1170;
  assign _EVAL_1203 = _EVAL_195 & _EVAL_1444;
  assign fanin__EVAL_75 = _EVAL_700;
  assign _EVAL_916 = _EVAL_3349[122];
  assign fanin__EVAL_98 = _EVAL_2384;
  assign gateways_gateway_52__EVAL_0 = _EVAL_9;
  assign fanin__EVAL_9 = _EVAL_2030;
  assign _EVAL_1504 = _EVAL_1949 | gateways_gateway_13__EVAL_4;
  assign _EVAL_1605 = _EVAL_1516 ? {{29'd0}, _EVAL_2309} : _EVAL_2140;
  assign _EVAL_870 = _EVAL_195 & _EVAL_2224;
  assign gateways_gateway_44__EVAL = _EVAL_71;
  assign _EVAL_1516 = 10'h38 == _EVAL_2998;
  assign _EVAL_980 = _EVAL_3349[77];
  assign _EVAL_440 = _EVAL_3251 ? {{29'd0}, _EVAL_3063} : _EVAL_1481;
  assign _EVAL_294 = _EVAL_651[37];
  assign gateways_gateway_40__EVAL_0 = _EVAL_9;
  assign _EVAL_567 = ~_EVAL_3782;
  assign _EVAL_321 = _EVAL_997 ? {{29'd0}, _EVAL_3711} : _EVAL_170;
  assign gateways_gateway_109__EVAL_3 = _EVAL_110;
  assign gateways_gateway_38__EVAL_2 = _EVAL_2917[39];
  assign gateways_gateway_101__EVAL_2 = _EVAL_2917[102];
  assign gateways_gateway_105__EVAL_1 = ~_EVAL_168;
  assign _EVAL_2147 = _EVAL_195 & _EVAL_1311;
  assign fanin__EVAL_62 = _EVAL_1789;
  assign _EVAL_753 = _EVAL_3349[13];
  assign gateways_gateway_35__EVAL_0 = _EVAL_9;
  assign gateways_gateway_60__EVAL = _EVAL_36;
  assign _EVAL_213 = _EVAL_651[512];
  assign _EVAL_1444 = _EVAL_651[99];
  assign _EVAL_771 = ~_EVAL_520;
  assign _EVAL_2653 = _EVAL_195 & _EVAL_3223;
  assign _EVAL_1954 = ~_EVAL_1122;
  assign gateways_gateway_66__EVAL = _EVAL_22;
  assign gateways_gateway_49__EVAL = _EVAL_127;
  assign _EVAL_2745 = out_back__EVAL_1[7:0];
  assign gateways_gateway_89__EVAL_0 = _EVAL_9;
  assign gateways_gateway_10__EVAL_0 = _EVAL_9;
  assign gateways_gateway_39__EVAL_3 = _EVAL_110;
  assign _EVAL_1765 = _EVAL_195 & _EVAL_3651;
  assign _EVAL_3205 = _EVAL_602 & _EVAL_826;
  assign _EVAL_3225 = {{28'd0}, _EVAL_2352};
  assign _EVAL_2938 = _EVAL_1193 ? {{29'd0}, _EVAL_2921} : _EVAL_3471;
  assign _EVAL_434 = _EVAL_3566 ? {{29'd0}, _EVAL_1459} : _EVAL_309;
  assign _EVAL_3775 = _EVAL_3652 & _EVAL_826;
  assign _EVAL_1773 = _EVAL_2772 | gateways_gateway_120__EVAL_4;
  assign gateways_gateway_111__EVAL_2 = _EVAL_2917[112];
  assign _EVAL_2227 = out_back__EVAL_3[19];
  assign _EVAL_2328 = _EVAL_3762 & _EVAL_2035;
  assign _EVAL_404 = 10'h4f == _EVAL_2998;
  assign _EVAL_847 = _EVAL_195 & _EVAL_1066;
  assign _EVAL_3626 = ~_EVAL_2482;
  assign gateways_gateway_121__EVAL_1 = ~_EVAL_668;
  assign _EVAL_2672 = _EVAL_3533 ? _EVAL_826 : _EVAL_3510;
  assign _EVAL_2460 = ~_EVAL_1184;
  assign _EVAL_1014 = _EVAL_323 & _EVAL_826;
  assign _EVAL_148 = _EVAL_3039 | gateways_gateway_43__EVAL_4;
  assign _EVAL_2440 = out_back__EVAL_3 & 20'h7f380;
  assign _EVAL_1243 = _EVAL_3349[95];
  assign gateways_gateway_88__EVAL = _EVAL_28;
  assign gateways_gateway_18__EVAL = _EVAL_102;
  assign _EVAL_2230 = _EVAL_1046 ? {{29'd0}, _EVAL_513} : _EVAL_3461;
  assign _EVAL_304 = {_EVAL_2469,_EVAL_3166,_EVAL_3397,_EVAL_2450};
  assign gateways_gateway_41__EVAL_3 = _EVAL_110;
  assign _EVAL_3056 = _EVAL_467 & _EVAL_2035;
  assign _EVAL_3349 = 128'h1 << _EVAL_1411;
  assign _EVAL_2904 = _EVAL_3349[36];
  assign gateways_gateway_97__EVAL = _EVAL_75;
  assign _EVAL_3186 = 10'h32 == _EVAL_2998;
  assign _EVAL_2658 = _EVAL_1281 & _EVAL_2035;
  assign gateways_gateway_25__EVAL_2 = _EVAL_2917[26];
  assign _EVAL_3567 = _EVAL_1017 ? _EVAL_826 : _EVAL_775;
  assign _EVAL_3801 = _EVAL_195 & _EVAL_2855;
  assign _EVAL_2069 = _EVAL_2525 ? {{29'd0}, _EVAL_2004} : _EVAL_2872;
  assign gateways_gateway_119__EVAL = _EVAL_50;
  assign _EVAL_3035 = ~_EVAL_3104;
  assign _EVAL_640 = _EVAL_651[30];
  assign _EVAL_3127 = _EVAL_1002 & _EVAL_826;
  assign gateways_gateway_91__EVAL_3 = _EVAL_110;
  assign _EVAL_3597 = _EVAL_2438 & _EVAL_826;
  assign _EVAL_3001 = _EVAL_245 & _EVAL_826;
  assign gateways_gateway_31__EVAL_1 = ~_EVAL_3112;
  assign _EVAL_339 = _EVAL_1812 ? {{29'd0}, _EVAL_1199} : _EVAL_150;
  assign _EVAL_2661 = _EVAL_2892 & _EVAL_2035;
  assign _EVAL_1278 = _EVAL_1768 & _EVAL_826;
  assign _EVAL_1422 = ~_EVAL_1191;
  assign _EVAL_3155 = _EVAL_410 | gateways_gateway__EVAL_4;
  assign _EVAL_1056 = _EVAL_2557 ? _EVAL_826 : _EVAL_3326;
  assign _EVAL_313 = _EVAL_3201 ? {{29'd0}, _EVAL_3080} : _EVAL_3262;
  assign _EVAL_3523 = _EVAL_3349[56];
  assign _EVAL_3265 = out_back__EVAL_1[15:8];
  assign gateways_gateway_53__EVAL_1 = ~_EVAL_3150;
  assign fanin__EVAL_45 = _EVAL_3653;
  assign gateways_gateway_18__EVAL_2 = _EVAL_2917[19];
  assign gateways_gateway_21__EVAL_0 = _EVAL_9;
  assign _EVAL_3717 = _EVAL_651[122];
  assign gateways_gateway_105__EVAL_2 = _EVAL_2917[106];
  assign _EVAL_2856 = _EVAL_195 & _EVAL_1505;
  assign gateways_gateway_19__EVAL_1 = ~_EVAL_612;
  assign _EVAL_3537 = 10'h80 == _EVAL_2998;
  assign gateways_gateway_117__EVAL_3 = _EVAL_110;
  assign gateways_gateway_105__EVAL_0 = _EVAL_9;
  assign _EVAL_2008 = _EVAL_3463 ? _EVAL_826 : _EVAL_3708;
  assign fanin__EVAL_112 = _EVAL_854;
  assign gateways_gateway_71__EVAL_1 = ~_EVAL_2509;
  assign _EVAL_1143 = _EVAL_2868 ? _EVAL_826 : _EVAL_2992;
  assign _EVAL_1956 = _EVAL_651[78];
  assign fanin__EVAL_36 = _EVAL_1695;
  assign _EVAL_3430 = _EVAL_374 ? {{29'd0}, _EVAL_1005} : _EVAL_2062;
  assign _EVAL_2303 = _EVAL_1274 ? _EVAL_826 : _EVAL_758;
  assign gateways_gateway_57__EVAL = _EVAL_61;
  assign gateways_gateway_28__EVAL_3 = _EVAL_110;
  assign _EVAL_962 = ~_EVAL_1264;
  assign gateways_gateway_74__EVAL_3 = _EVAL_110;
  assign _EVAL_1741 = _EVAL_1046 ? _EVAL_826 : _EVAL_991;
  assign fanin__EVAL_50 = _EVAL_517;
  assign gateways_gateway_100__EVAL_1 = ~_EVAL_2197;
  assign gateways_gateway_48__EVAL_1 = ~_EVAL_1928;
  assign _EVAL_2478 = _EVAL_130[27:2];
  assign gateways_gateway_76__EVAL_2 = _EVAL_2917[77];
  assign gateways_gateway_37__EVAL_1 = ~_EVAL_3527;
  assign _EVAL_2168 = _EVAL_651[91];
  assign _EVAL_1396 = _EVAL_651[12];
  assign gateways_gateway_70__EVAL = _EVAL_109;
  assign gateways_gateway_83__EVAL_0 = _EVAL_9;
  assign gateways_gateway_23__EVAL_2 = _EVAL_2917[24];
  assign _EVAL_354 = _EVAL_381 & _EVAL_826;
  assign gateways_gateway_59__EVAL_3 = _EVAL_110;
  assign _EVAL_3077 = _EVAL_1096 ? {{29'd0}, _EVAL_3734} : _EVAL_669;
  assign _EVAL_995 = ~_EVAL_858;
  assign _EVAL_1896 = _EVAL_2559 & _EVAL_2035;
  assign fanin__EVAL_94 = _EVAL_1647;
  assign out_back__EVAL_0 = _EVAL_2478[19:0];
  assign gateways_gateway_38__EVAL_3 = _EVAL_110;
  assign gateways_gateway_32__EVAL_0 = _EVAL_9;
  assign _EVAL_2462 = _EVAL_3221 ? _EVAL_826 : _EVAL_2537;
  assign _EVAL_1697 = 10'h48 == _EVAL_2998;
  assign gateways_gateway_113__EVAL = _EVAL_74;
  assign _EVAL_2734 = _EVAL_330 & _EVAL_2035;
  assign _EVAL_225 = 10'h102 == _EVAL_2998;
  assign _EVAL_1601 = _EVAL_3349[47];
  assign gateways_gateway_78__EVAL = _EVAL_52;
  assign _EVAL_801 = _EVAL_3349[52];
  assign gateways_gateway_26__EVAL_1 = ~_EVAL_2143;
  assign gateways_gateway_103__EVAL_1 = ~_EVAL_813;
  assign gateways_gateway_98__EVAL_0 = _EVAL_9;
  assign _EVAL_2114 = {_EVAL_3346,_EVAL_3150,_EVAL_1749,_EVAL_3014,_EVAL_819,_EVAL_1638,_EVAL_1928,_EVAL_3059};
  assign _EVAL_446 = 10'h10 == _EVAL_2998;
  assign fanin__EVAL_78 = _EVAL_3191;
  assign gateways_gateway_124__EVAL_3 = _EVAL_110;
  assign _EVAL_904 = _EVAL_3349[113];
  assign _EVAL_205 = _EVAL_531 & _EVAL_2035;
  assign _EVAL_224 = {_EVAL_2698,_EVAL_813,_EVAL_2488,_EVAL_2160,_EVAL_2197,_EVAL_3656,_EVAL_3395,_EVAL_325,_EVAL_3200,
    _EVAL_415};
  assign _EVAL_3361 = _EVAL_3291 ? _EVAL_826 : _EVAL_925;
  assign _EVAL_2484 = _EVAL_651[57];
  assign _EVAL_858 = _EVAL_3349[103];
  assign _EVAL_3397 = {_EVAL_3420,_EVAL_3331,_EVAL_350,_EVAL_1392,_EVAL_1369,_EVAL_3508,_EVAL_423,_EVAL_2502,_EVAL_2114,
    _EVAL_2694};
  assign gateways_gateway_46__EVAL_0 = _EVAL_9;
  assign _EVAL_3524 = _EVAL_651[48];
  assign gateways_gateway_22__EVAL = _EVAL_42;
  assign _EVAL_604 = _EVAL_1101 & _EVAL_2035;
  assign _EVAL_2917 = _EVAL_1560 ? _EVAL_3015 : 128'h0;
  assign _EVAL_2787 = ~_EVAL_2222;
  assign _EVAL_2454 = _EVAL_3775 & _EVAL_2035;
  assign gateways_gateway_76__EVAL_3 = _EVAL_110;
  assign _EVAL_3000 = _EVAL_195 & _EVAL_1053;
  assign _EVAL_2791 = _EVAL_1052 ? {{29'd0}, _EVAL_1527} : _EVAL_3714;
  assign _EVAL_544 = _EVAL_1987 ? _EVAL_826 : _EVAL_696;
  assign _EVAL_1596 = _EVAL_1794 & _EVAL_2035;
  assign gateways_gateway_103__EVAL_3 = _EVAL_110;
  assign _EVAL_3652 = _EVAL_195 & _EVAL_294;
  assign gateways_gateway_8__EVAL_0 = _EVAL_9;
  assign _EVAL_3490 = _EVAL_195 & _EVAL_340;
  assign _EVAL_2472 = {_EVAL_2174,_EVAL_2165,_EVAL_911,_EVAL_3213,_EVAL_1120,_EVAL_3824,_EVAL_552,_EVAL_3140,_EVAL_2627,
    _EVAL_3214};
  assign _EVAL_2626 = _EVAL_2811 ? _EVAL_826 : _EVAL_1143;
  assign _EVAL_703 = ~_EVAL_1183;
  assign gateways_gateway_8__EVAL_3 = _EVAL_110;
  assign _EVAL_2064 = _EVAL_3104 | gateways_gateway_108__EVAL_4;
  assign _EVAL_1830 = _EVAL_651[65];
  assign _EVAL_180 = _EVAL_1597 & _EVAL_2035;
  assign _EVAL_1093 = _EVAL_1500 ? {{29'd0}, _EVAL_3505} : _EVAL_2078;
  assign _EVAL_314 = _EVAL_195 & _EVAL_3414;
  assign _EVAL_3370 = _EVAL_1869 ? {{29'd0}, _EVAL_2182} : _EVAL_1415;
  assign gateways_gateway_61__EVAL_2 = _EVAL_2917[62];
  assign _EVAL_1720 = _EVAL_3037 & _EVAL_2035;
  assign _EVAL_2811 = 10'h78 == _EVAL_2998;
  assign gateways_gateway_77__EVAL_1 = ~_EVAL_1524;
  assign gateways_gateway_73__EVAL_2 = _EVAL_2917[74];
  assign gateways_gateway_26__EVAL_3 = _EVAL_110;
  assign _EVAL_3153 = 10'h7d == _EVAL_2998;
  assign _EVAL_2397 = 10'h73 == _EVAL_2998;
  assign _EVAL_270 = _EVAL_3381 | gateways_gateway_65__EVAL_4;
  assign gateways_gateway_45__EVAL_3 = _EVAL_110;
  assign _EVAL_2439 = _EVAL_272 | gateways_gateway_5__EVAL_4;
  assign _EVAL_451 = 10'h26 == _EVAL_2998;
  assign _EVAL_2874 = _EVAL_651[29];
  assign _EVAL_3494 = _EVAL_1483 & _EVAL_2035;
  assign _EVAL_793 = ~_EVAL_2622;
  assign _EVAL_2927 = _EVAL_987 ? _EVAL_826 : _EVAL_2999;
  assign _EVAL_2233 = _EVAL_651[23];
  assign _EVAL_2350 = ~_EVAL_341;
  assign _EVAL_3700 = _EVAL_3349[48];
  assign gateways_gateway_58__EVAL_2 = _EVAL_2917[59];
  assign gateways_gateway_96__EVAL_1 = ~_EVAL_3200;
  assign _EVAL_1952 = _EVAL_504 ? _EVAL_826 : _EVAL_1540;
  assign _EVAL_991 = _EVAL_3537 ? _EVAL_826 : _EVAL_2476;
  assign _EVAL_3436 = ~_EVAL_1880;
  assign _EVAL_2759 = _EVAL_3596 ? _EVAL_826 : _EVAL_2626;
  assign gateways_gateway_108__EVAL_0 = _EVAL_9;
  assign _EVAL_196 = _EVAL_2727 & _EVAL_826;
  assign gateways_gateway_100__EVAL_0 = _EVAL_9;
  assign _EVAL_2403 = _EVAL_3328 & _EVAL_425;
  assign _EVAL_3474 = _EVAL_2881 ? _EVAL_826 : _EVAL_3101;
  assign gateways_gateway_20__EVAL_2 = _EVAL_2917[21];
  assign _EVAL_2198 = _EVAL_2555 & _EVAL_2035;
  assign gateways_gateway_34__EVAL_0 = _EVAL_9;
  assign gateways_gateway_87__EVAL_2 = _EVAL_2917[88];
  assign _EVAL_2226 = _EVAL_1118 ? {{29'd0}, _EVAL_1692} : _EVAL_970;
  assign _EVAL_2902 = {_EVAL_445,_EVAL_2121,_EVAL_3850,_EVAL_3654,_EVAL_1030,_EVAL_1548,_EVAL_930,_EVAL_1925};
  assign _EVAL_2131 = _EVAL_1799 ? _EVAL_826 : _EVAL_1419;
  assign gateways_gateway_34__EVAL_3 = _EVAL_110;
  assign _EVAL_1637 = _EVAL_994 ? _EVAL_826 : _EVAL_3388;
  assign gateways_gateway_59__EVAL_0 = _EVAL_9;
  assign gateways_gateway_88__EVAL_0 = _EVAL_9;
  assign _EVAL_1750 = _EVAL_3427 & _EVAL_425;
  assign _EVAL_1094 = _EVAL_651[59];
  assign _EVAL_1684 = _EVAL_1428 | gateways_gateway_66__EVAL_4;
  assign _EVAL_848 = ~_EVAL_3633;
  assign _EVAL_324 = _EVAL_1990 & _EVAL_826;
  assign _EVAL_228 = ~_EVAL_1269;
  assign _EVAL_685 = ~_EVAL_1949;
  assign gateways_gateway_114__EVAL_1 = ~_EVAL_2193;
  assign _EVAL_850 = _EVAL_299 ? _EVAL_826 : _EVAL_2927;
  assign gateways_gateway_24__EVAL_3 = _EVAL_110;
  assign _EVAL_3449 = _EVAL_1308 & _EVAL_826;
  assign _EVAL_2521 = _EVAL_695 ? _EVAL_826 : _EVAL_3847;
  assign _EVAL_2498 = ~_EVAL_655;
  assign gateways_gateway_29__EVAL_1 = ~_EVAL_1434;
  assign gateways_gateway_72__EVAL_3 = _EVAL_110;
  assign _EVAL_2321 = _EVAL_1960 & _EVAL_826;
  assign _EVAL_3106 = ~_EVAL_963;
  assign _EVAL_794 = _EVAL_651[84];
  assign gateways_gateway_121__EVAL_0 = _EVAL_9;
  assign _EVAL_2015 = _EVAL_1688 & _EVAL_2035;
  assign gateways_gateway_119__EVAL_3 = _EVAL_110;
  assign _EVAL_1303 = _EVAL_1680 & _EVAL_826;
  assign _EVAL_1473 = _EVAL_643 | gateways_gateway_57__EVAL_4;
  assign gateways_gateway_81__EVAL_2 = _EVAL_2917[82];
  assign _EVAL_3040 = _EVAL_2758[0];
  assign gateways_gateway_99__EVAL_3 = _EVAL_110;
  assign fanin__EVAL_4 = _EVAL_2281;
  assign fanin__EVAL_82 = _EVAL_2996;
  assign _EVAL_410 = _EVAL_3349[1];
  assign _EVAL_3033 = _EVAL_2738 ? {{29'd0}, _EVAL_289} : _EVAL_339;
  assign _EVAL_2342 = _EVAL_195 & _EVAL_1371;
  assign _EVAL_856 = 10'h50 == _EVAL_2998;
  assign gateways_gateway_9__EVAL = _EVAL_27;
  assign _EVAL_3094 = _EVAL_195 & _EVAL_3717;
  assign _EVAL_1852 = _EVAL_651[87];
  assign _EVAL_3172 = _EVAL_195 & _EVAL_3249;
  assign gateways_gateway_69__EVAL = _EVAL_117;
  assign _EVAL_3529 = _EVAL_195 & _EVAL_3243;
  assign _EVAL_2352 = {1'h0,_EVAL_3156};
  assign _EVAL_2697 = out_back__EVAL_1[7:1];
  assign gateways_gateway_48__EVAL = _EVAL_63;
  assign gateways_gateway_10__EVAL_2 = _EVAL_2917[11];
  assign gateways_gateway_6__EVAL_0 = _EVAL_9;
  assign _EVAL_657 = _EVAL_3402 ? _EVAL_826 : _EVAL_1089;
  assign gateways_gateway_7__EVAL = _EVAL_0;
  assign _EVAL_560 = _EVAL_651[61];
  assign _EVAL_3322 = 10'he == _EVAL_2998;
  assign _EVAL_171 = 10'h30 == _EVAL_2998;
  assign _EVAL_2977 = _EVAL_1718 & _EVAL_826;
  assign _EVAL_804 = ~_EVAL_1430;
  assign _EVAL_3076 = _EVAL_225 ? _EVAL_832 : _EVAL_1036;
  assign gateways_gateway_68__EVAL_2 = _EVAL_2917[69];
  assign _EVAL_3124 = _EVAL_3086 ? {{29'd0}, _EVAL_2637} : _EVAL_3692;
  assign _EVAL_3680 = _EVAL_1172 ? {{29'd0}, _EVAL_2262} : _EVAL_440;
  assign _EVAL_2530 = ~_EVAL_3341;
  assign _EVAL_3240 = {_EVAL_3589,_EVAL_2396,_EVAL_1872,_EVAL_872,_EVAL_3043,_EVAL_168,_EVAL_2698,_EVAL_813,_EVAL_428};
  assign _EVAL_2134 = _EVAL_1183 | gateways_gateway_74__EVAL_4;
  assign gateways_gateway_12__EVAL_1 = ~_EVAL_3824;
  assign _EVAL_2952 = _EVAL_3157 & _EVAL_2035;
  assign _EVAL_2885 = _EVAL_996 & _EVAL_826;
  assign _EVAL_2537 = _EVAL_1547 ? _EVAL_826 : _EVAL_1443;
  assign fanin__EVAL_2 = _EVAL_2466;
  assign gateways_gateway_42__EVAL_0 = _EVAL_9;
  assign fanin__EVAL_126 = _EVAL_853;
  assign fanin__EVAL_6 = _EVAL_2262;
  assign gateways_gateway_39__EVAL_2 = _EVAL_2917[40];
  assign fanin__EVAL_18 = _EVAL_797;
  assign fanin__EVAL = _EVAL_2182;
  assign gateways_gateway_99__EVAL = _EVAL_53;
  assign _EVAL_2009 = 10'h5e == _EVAL_2998;
  assign fanin__EVAL_111 = _EVAL_2306;
  assign _EVAL_868 = _EVAL_1112 & _EVAL_2035;
  assign _EVAL_699 = _EVAL_1439 ? _EVAL_826 : _EVAL_1032;
  assign gateways_gateway_22__EVAL_2 = _EVAL_2917[23];
  assign _EVAL_2270 = _EVAL_2191 & _EVAL_2035;
  assign gateways_gateway_21__EVAL_3 = _EVAL_110;
  assign _EVAL_584 = 10'h15 == _EVAL_2998;
  assign _EVAL_3211 = _EVAL_651[76];
  assign _EVAL_2795 = _EVAL_651[27];
  assign gateways_gateway_74__EVAL_2 = _EVAL_2917[75];
  assign gateways_gateway_44__EVAL_2 = _EVAL_2917[45];
  assign _EVAL_3735 = _EVAL_2055 & _EVAL_2035;
  assign _EVAL_2702 = _EVAL_3312 & _EVAL_826;
  assign _EVAL_3099 = _EVAL_651[20];
  assign gateways_gateway_77__EVAL = _EVAL_35;
  assign fanin__EVAL_103 = _EVAL_461;
  assign _EVAL_2222 = _EVAL_3349[26];
  assign fanin__EVAL_47 = _EVAL_513;
  assign gateways_gateway_91__EVAL = _EVAL_62;
  assign _EVAL_3307 = _EVAL_2408 ? _EVAL_826 : _EVAL_1595;
  assign gateways_gateway_113__EVAL_1 = ~_EVAL_2618;
  assign _EVAL_3787 = _EVAL_3185 & _EVAL_2035;
  assign _EVAL_918 = ~_EVAL_2822;
  assign fanin__EVAL_114 = _EVAL_2580;
  assign gateways_gateway_15__EVAL = _EVAL_88;
  assign _EVAL_2316 = _EVAL_3349[79];
  assign _EVAL_1426 = _EVAL_3427 & _EVAL_678;
  assign _EVAL_832 = {_EVAL_1340,_EVAL_1380,_EVAL_394,_EVAL_2877};
  assign _EVAL_3198 = _EVAL_1824 ? {{29'd0}, _EVAL_1805} : _EVAL_2060;
  assign _EVAL_2880 = _EVAL_195 & _EVAL_3036;
  assign _EVAL_1374 = _EVAL_1547 ? {{29'd0}, _EVAL_853} : _EVAL_689;
  assign _EVAL_500 = _EVAL_1171 ? _EVAL_845 : _EVAL_2361;
  assign gateways_gateway_49__EVAL_1 = ~_EVAL_1638;
  assign _EVAL_799 = _EVAL_3130 & _EVAL_2035;
  assign fanin__EVAL_83 = _EVAL_3063;
  assign gateways_gateway_53__EVAL = _EVAL_76;
  assign gateways_gateway__EVAL_2 = _EVAL_2917[1];
  assign _EVAL_506 = _EVAL_651[21];
  assign gateways_gateway_13__EVAL_2 = _EVAL_2917[14];
  assign fanin__EVAL_39 = _EVAL_3624;
  assign _EVAL_3715 = _EVAL_1303 & _EVAL_2035;
  assign gateways_gateway_123__EVAL = _EVAL_94;
  assign fanin__EVAL_101 = _EVAL_2186;
  assign gateways_gateway_63__EVAL_0 = _EVAL_9;
  assign _EVAL_1034 = _EVAL_1174 ? _EVAL_826 : _EVAL_657;
  assign _EVAL_2801 = _EVAL_1039 & _EVAL_826;
  assign _EVAL_3591 = _EVAL_3153 ? {{29'd0}, _EVAL_1268} : _EVAL_1871;
  assign _EVAL_275 = _EVAL_273 & _EVAL_2035;
  assign _EVAL_1349 = ~_EVAL_3557;
  assign _EVAL_2503 = _EVAL_3349[32];
  assign gateways_gateway_30__EVAL_0 = _EVAL_9;
  assign _EVAL_2983 = _EVAL_651[68];
  assign _EVAL_1130 = _EVAL_385 ? _EVAL_3225 : _EVAL_1315;
  assign _EVAL_2318 = _EVAL_536 & _EVAL_2035;
  assign _EVAL_1476 = _EVAL_3718 & _EVAL_2035;
  assign _EVAL_2568 = _EVAL_1857 ? _EVAL_826 : _EVAL_265;
  assign gateways_gateway_39__EVAL_0 = _EVAL_9;
  assign fanin__EVAL_10 = _EVAL_289;
  assign gateways_gateway_23__EVAL_3 = _EVAL_110;
  assign gateways_gateway_125__EVAL_0 = _EVAL_9;
  assign _EVAL_3534 = _EVAL_337 ? _EVAL_826 : _EVAL_2441;
  assign gateways_gateway_62__EVAL_1 = ~_EVAL_3420;
  assign _EVAL_653 = _EVAL_2527 | gateways_gateway_9__EVAL_4;
  assign _EVAL_2615 = _EVAL_1899 & _EVAL_2035;
  assign _EVAL_1555 = ~_EVAL_2320;
  assign fanin__EVAL_123 = _EVAL_3315;
  assign _EVAL_2084 = _EVAL_2850[2:0];
  assign gateways_gateway_105__EVAL = _EVAL_93;
  assign _EVAL_1135 = _EVAL_651[36];
  assign _EVAL_1542 = _EVAL_3349[33];
  assign gateways_gateway_86__EVAL_2 = _EVAL_2917[87];
  assign _EVAL_894 = _EVAL_3596 ? {{29'd0}, _EVAL_865} : _EVAL_2663;
  assign gateways_gateway_118__EVAL_0 = _EVAL_9;
  assign _EVAL_2322 = _EVAL_3349[72];
  assign gateways_gateway_46__EVAL_1 = ~_EVAL_3242;
  assign fanin__EVAL_35 = _EVAL_2079;
  assign _EVAL_175 = {_EVAL_1710,_EVAL_1147,_EVAL_1417,_EVAL_2178,_EVAL_2903};
  assign _EVAL_223 = _EVAL_2218 & _EVAL_2035;
  assign _EVAL_402 = _EVAL_651[33];
  assign _EVAL_892 = _EVAL_994 ? {{29'd0}, _EVAL_2711} : _EVAL_321;
  assign _EVAL_1218 = _EVAL_2942 & _EVAL_2035;
  assign gateways_gateway_80__EVAL_1 = ~_EVAL_2297;
  assign _EVAL_3263 = {_EVAL_2143,_EVAL_3268,_EVAL_2370,_EVAL_3129,_EVAL_1964,_EVAL_302,_EVAL_1467,_EVAL_612,_EVAL_498,
    _EVAL_2472};
  assign _EVAL_2565 = _EVAL_3186 ? _EVAL_826 : _EVAL_3465;
  assign _EVAL_3701 = _EVAL_651[42];
  assign gateways_gateway_19__EVAL = _EVAL_99;
  assign _EVAL_1711 = _EVAL_3299 ? _EVAL_826 : _EVAL_2926;
  assign _EVAL_2455 = _EVAL_195 & _EVAL_2795;
  assign _EVAL_1932 = {_EVAL_1030,_EVAL_1548,_EVAL_930,_EVAL_1925,1'h0};
  assign _EVAL_2612 = _EVAL_1879 ? _EVAL_826 : _EVAL_1952;
  assign _EVAL_259 = _EVAL_3834 & _EVAL_2035;
  assign gateways_gateway_70__EVAL_1 = ~_EVAL_1365;
  assign _EVAL_3189 = _EVAL_2880 & _EVAL_826;
  assign gateways_gateway_64__EVAL_2 = _EVAL_2917[65];
  assign _EVAL_1657 = _EVAL_3105 | gateways_gateway_95__EVAL_4;
  assign _EVAL_1187 = _EVAL_3349[94];
  assign _EVAL_1712 = _EVAL_651[45];
  assign _EVAL_3086 = 10'h2 == _EVAL_2998;
  assign _EVAL_1086 = _EVAL_651[105];
  assign fanin__EVAL_49 = _EVAL_1005;
  assign _EVAL_687 = _EVAL_1446 & _EVAL_2035;
  assign _EVAL_2586 = _EVAL_1435 ? _EVAL_826 : _EVAL_3772;
  assign _EVAL_258 = _EVAL_3349[73];
  assign _EVAL_2814 = _EVAL_651[25];
  assign _EVAL_2132 = _EVAL_1011 | gateways_gateway_119__EVAL_4;
  assign gateways_gateway_79__EVAL = _EVAL_118;
  assign gateways_gateway_57__EVAL_0 = _EVAL_9;
  assign _EVAL_610 = _EVAL_655 | gateways_gateway_99__EVAL_4;
  assign _EVAL_613 = _EVAL_354 & _EVAL_2035;
  assign out_back__EVAL_13 = _EVAL_110;
  assign _EVAL_762 = ~_EVAL_1480;
  assign gateways_gateway_86__EVAL_3 = _EVAL_110;
  assign _EVAL_3422 = ~_EVAL_1011;
  assign _EVAL_1537 = _EVAL_1554 ? _EVAL_826 : _EVAL_2632;
  assign _EVAL_3809 = _EVAL_3427 & _EVAL_3266;
  assign _EVAL_3662 = _EVAL_2321 & _EVAL_2035;
  assign gateways_gateway_71__EVAL_2 = _EVAL_2917[72];
  assign gateways_gateway_16__EVAL_2 = _EVAL_2917[17];
  assign gateways_gateway_87__EVAL = _EVAL_144;
  assign _EVAL_3526 = |_EVAL_2850;
  assign _EVAL_615 = _EVAL_1452 & _EVAL_826;
  assign _EVAL_2220 = _EVAL_651[67];
  assign _EVAL_3384 = _EVAL_651[102];
  assign gateways_gateway_5__EVAL_1 = ~_EVAL_2685;
  assign _EVAL_2130 = ~_EVAL_2686;
  assign _EVAL_2179 = _EVAL_195 & _EVAL_338;
  assign gateways_gateway_37__EVAL_2 = _EVAL_2917[38];
  assign _EVAL_2078 = _EVAL_1174 ? {{29'd0}, _EVAL_1528} : _EVAL_2486;
  assign gateways_gateway_17__EVAL_3 = _EVAL_110;
  assign gateways_gateway_107__EVAL_3 = _EVAL_110;
  assign _EVAL_3577 = _EVAL_1813 & _EVAL_826;
  assign _EVAL_1739 = _EVAL_2810 & _EVAL_826;
  assign gateways_gateway_29__EVAL_2 = _EVAL_2917[30];
  assign _EVAL_1065 = ~_EVAL_3599;
  assign _EVAL_2788 = _EVAL_3349[60];
  assign _EVAL_710 = ~_EVAL_1630;
  assign _EVAL_301 = _EVAL_195 & _EVAL_693;
  assign _EVAL_3620 = _EVAL_2019 ? _EVAL_826 : _EVAL_2568;
  assign _EVAL_309 = _EVAL_179 ? {{29'd0}, _EVAL_1968} : _EVAL_1882;
  assign _EVAL_3632 = _EVAL_3378 | gateways_gateway_81__EVAL_4;
  assign _EVAL_2554 = _EVAL_195 & _EVAL_213;
  assign _EVAL_2663 = _EVAL_2811 ? {{29'd0}, _EVAL_2878} : _EVAL_1702;
  assign _EVAL_743 = _EVAL_595 ? {{29'd0}, _EVAL_1687} : _EVAL_2789;
  assign gateways_gateway_87__EVAL_1 = ~_EVAL_2799;
  assign _EVAL_1985 = ~_EVAL_980;
  assign _EVAL_3414 = _EVAL_651[110];
  assign _EVAL_1815 = ~_EVAL_726;
  assign _EVAL_2123 = _EVAL_1385 & _EVAL_3526;
  assign _EVAL_1529 = _EVAL_3172 & _EVAL_826;
  assign _EVAL_247 = _EVAL_1180 | gateways_gateway_70__EVAL_4;
  assign _EVAL_3067 = _EVAL_1074 & _EVAL_826;
  assign _EVAL_2798 = _EVAL_651[19];
  assign _EVAL_1618 = _EVAL_3349[12];
  assign gateways_gateway_81__EVAL = _EVAL_116;
  assign _EVAL_733 = _EVAL_913 & _EVAL_826;
  assign fanin__EVAL_26 = _EVAL_2878;
  assign gateways_gateway_98__EVAL = _EVAL_141;
  assign _EVAL_2090 = _EVAL_2077 | gateways_gateway_105__EVAL_4;
  assign fanin__EVAL_121 = _EVAL_3798;
  assign _EVAL_3075 = _EVAL_3434 ? {{29'd0}, _EVAL_3013} : _EVAL_2722;
  assign gateways_gateway_102__EVAL_1 = ~_EVAL_2488;
  assign _EVAL_2327 = _EVAL_3001 & _EVAL_2035;
  assign _EVAL_3569 = _EVAL_1670 ? _EVAL_826 : _EVAL_2254;
  assign _EVAL_641 = ~_EVAL_1033;
  assign gateways_gateway_73__EVAL_1 = ~_EVAL_2682;
  assign _EVAL_2362 = _EVAL_733 & _EVAL_2035;
  assign _EVAL_3376 = ~_EVAL_3392;
  assign _EVAL_2850 = {_EVAL_1587,_EVAL_1696,_EVAL_1723,_EVAL_3241};
  assign _EVAL_209 = _EVAL_195 & _EVAL_1280;
  assign _EVAL_2113 = _EVAL_1251 & _EVAL_2035;
  assign _EVAL_1877 = _EVAL_651[43];
  assign gateways_gateway_47__EVAL = _EVAL_133;
  assign gateways_gateway_23__EVAL_0 = _EVAL_9;
  assign _EVAL_2389 = _EVAL_3433 & _EVAL_826;
  assign _EVAL_1521 = _EVAL_2217 & _EVAL_2035;
  assign gateways_gateway_45__EVAL = _EVAL_139;
  assign gateways_gateway_92__EVAL_0 = _EVAL_9;
  assign _EVAL_1053 = _EVAL_651[70];
  assign _EVAL_925 = _EVAL_2738 ? _EVAL_826 : _EVAL_161;
  assign _EVAL_3255 = _EVAL_651[1];
  assign _EVAL_1299 = _EVAL_3367 ? {{29'd0}, _EVAL_1134} : _EVAL_3124;
  assign _EVAL_3782 = _EVAL_3349[117];
  assign _EVAL_3603 = _EVAL_3256 ? _EVAL_826 : _EVAL_2074;
  assign _EVAL_841 = _EVAL_195 & _EVAL_1086;
  assign _EVAL_515 = _EVAL_651[107];
  assign _EVAL_2378 = _EVAL_3467 ? _EVAL_826 : _EVAL_3418;
  assign _EVAL_2639 = {{25'd0}, _EVAL_2757};
  assign gateways_gateway_37__EVAL_3 = _EVAL_110;
  assign _EVAL_3786 = _EVAL_195 & _EVAL_1787;
  assign _EVAL_1076 = _EVAL_638 ? {{29'd0}, _EVAL_3825} : _EVAL_1000;
  assign _EVAL_2020 = _EVAL_1282 ? {{29'd0}, _EVAL_3657} : _EVAL_2654;
  assign gateways_gateway_4__EVAL_0 = _EVAL_9;
  assign fanin__EVAL_15 = _EVAL_3825;
  assign _EVAL_3249 = _EVAL_651[58];
  assign _EVAL_3074 = 10'h5f == _EVAL_2998;
  assign gateways_gateway_17__EVAL_0 = _EVAL_9;
  assign _EVAL_499 = 10'h82 == _EVAL_2998;
  assign _EVAL_371 = ~_EVAL_368;
  assign _EVAL_651 = 1024'h1 << _EVAL_2998;
  assign gateways_gateway_66__EVAL_2 = _EVAL_2917[67];
  assign _EVAL_964 = _EVAL_3349[42];
  assign _EVAL_1659 = _EVAL_1920 ? _EVAL_1932 : _EVAL_2300;
  assign _EVAL_2099 = _EVAL_3349[97];
  assign gateways_gateway_11__EVAL_3 = _EVAL_110;
  assign _EVAL_1046 = 10'h7f == _EVAL_2998;
  assign _EVAL_1998 = _EVAL_195 & _EVAL_3287;
  assign gateways_gateway_56__EVAL_0 = _EVAL_9;
  assign _EVAL_605 = _EVAL_3349[63];
  assign gateways_gateway_66__EVAL_0 = _EVAL_9;
  assign _EVAL_2021 = 10'h5d == _EVAL_2998;
  assign gateways_gateway_29__EVAL = _EVAL_115;
  assign gateways_gateway_123__EVAL_2 = _EVAL_2917[124];
  assign _EVAL_3082 = _EVAL_3186 ? {{29'd0}, _EVAL_3437} : _EVAL_3442;
  assign _EVAL_1797 = _EVAL_2474 & _EVAL_2035;
  assign _EVAL_2341 = _EVAL_3349[27];
  assign gateways_gateway_88__EVAL_1 = ~_EVAL_3107;
  assign gateways_gateway_77__EVAL_3 = _EVAL_110;
  assign gateways_gateway_53__EVAL_0 = _EVAL_9;
  assign gateways_gateway_72__EVAL = _EVAL_57;
  assign _EVAL_203 = _EVAL_3786 & _EVAL_826;
  assign _EVAL_3745 = _EVAL_1681 & _EVAL_2035;
  assign out_back__EVAL_16 = _EVAL_5;
  assign _EVAL_2660 = out_back__EVAL_3[1];
  assign _EVAL_469 = _EVAL_2850[7:0];
  assign _EVAL_2337 = _EVAL_274 | gateways_gateway_23__EVAL_4;
  assign _EVAL_2654 = _EVAL_3481 ? {{29'd0}, _EVAL_3357} : _EVAL_532;
  assign _EVAL_1496 = _EVAL_987 ? {{29'd0}, _EVAL_461} : _EVAL_1071;
  assign fanin__EVAL_23 = _EVAL_642;
  assign _EVAL_678 = &_EVAL_469;
  assign _EVAL_3185 = _EVAL_238 & _EVAL_826;
  assign gateways_gateway_83__EVAL = _EVAL_143;
  assign _EVAL_1181 = _EVAL_195 & _EVAL_2879;
  assign _EVAL_3800 = _EVAL_195 & _EVAL_625;
  assign gateways_gateway_43__EVAL_1 = ~_EVAL_2944;
  assign _EVAL_3029 = _EVAL_195 & _EVAL_817;
  assign _EVAL_2990 = _EVAL_1529 & _EVAL_2035;
  assign gateways_gateway_42__EVAL = _EVAL_114;
  assign gateways_gateway_26__EVAL_2 = _EVAL_2917[27];
  assign _EVAL_869 = 10'h7c == _EVAL_2998;
  assign _EVAL_1904 = _EVAL_2018 & _EVAL_2035;
  assign fanin__EVAL_56 = _EVAL_1341;
  assign gateways_gateway_67__EVAL_3 = _EVAL_110;
  assign gateways_gateway_41__EVAL_2 = _EVAL_2917[42];
  assign gateways_gateway_46__EVAL = _EVAL_21;
  assign _EVAL_480 = _EVAL_520 | gateways_gateway_37__EVAL_4;
  assign gateways_gateway_73__EVAL_3 = _EVAL_110;
  assign out_back__EVAL_15 = _EVAL_9;
  assign _EVAL_1509 = _EVAL_195 & _EVAL_212;
  assign gateways_gateway_113__EVAL_0 = _EVAL_9;
  assign gateways_gateway_36__EVAL_3 = _EVAL_110;
  assign gateways_gateway_52__EVAL_2 = _EVAL_2917[53];
  assign gateways_gateway_10__EVAL_3 = _EVAL_110;
  assign fanin__EVAL_52 = _EVAL_1085;
  assign gateways_gateway_55__EVAL_0 = _EVAL_9;
  assign _EVAL_2202 = _EVAL_3217 & _EVAL_826;
  assign _EVAL_1696 = _EVAL_588 ? 8'hff : 8'h0;
  assign _EVAL_3457 = ~_EVAL_3105;
  assign gateways_gateway_51__EVAL_0 = _EVAL_9;
  assign _EVAL_2907 = _EVAL_3349[115];
  assign _EVAL_1757 = _EVAL_2554 & _EVAL_826;
  assign _EVAL_403 = _EVAL_651[79];
  assign gateways_gateway_3__EVAL_3 = _EVAL_110;
  assign gateways_gateway_104__EVAL_0 = _EVAL_9;
  assign gateways_gateway_103__EVAL = _EVAL_58;
  assign _EVAL_3353 = ~_EVAL_272;
  assign _EVAL_1966 = _EVAL_2021 ? {{29'd0}, _EVAL_2828} : _EVAL_293;
  assign _EVAL_1040 = _EVAL_195 & _EVAL_1486;
  assign _EVAL_648 = _EVAL_195 & _EVAL_794;
  assign _EVAL_3264 = _EVAL_3138 | gateways_gateway_92__EVAL_4;
  assign _EVAL_1890 = ~_EVAL_3545;
  assign _EVAL_3183 = ~_EVAL_2251;
  assign gateways_gateway_3__EVAL = _EVAL_44;
  assign _EVAL_3244 = _EVAL_195 & _EVAL_3206;
  assign _EVAL_185 = 10'h3 == _EVAL_2998;
  assign _EVAL_473 = _EVAL_195 & _EVAL_463;
  assign gateways_gateway_85__EVAL_2 = _EVAL_2917[86];
  assign _EVAL_3392 = _EVAL_3349[23];
  assign _EVAL_2946 = _EVAL_3074 ? {{29'd0}, _EVAL_778} : _EVAL_3394;
  assign _EVAL_1452 = _EVAL_195 & _EVAL_379;
  assign _EVAL_1311 = _EVAL_651[90];
  assign _EVAL_3047 = 10'h6a == _EVAL_2998;
  assign _EVAL_2701 = ~_EVAL_735;
  assign _EVAL_3223 = _EVAL_651[71];
  assign _EVAL_1481 = _EVAL_3291 ? {{29'd0}, _EVAL_1963} : _EVAL_3033;
  assign _EVAL_2369 = ~_EVAL_2298;
  assign _EVAL_840 = _EVAL_651[6];
  assign _EVAL_2692 = _EVAL_1440 & _EVAL_826;
  assign _EVAL_3260 = ~_EVAL_646;
  assign _EVAL_1662 = _EVAL_1102 & _EVAL_2035;
  assign _EVAL_1781 = _EVAL_3094 & _EVAL_826;
  assign _EVAL_1715 = _EVAL_2257 & _EVAL_2035;
  assign gateways_gateway_36__EVAL_0 = _EVAL_9;
  assign _EVAL_1813 = _EVAL_195 & _EVAL_3435;
  assign fanin__EVAL_108 = _EVAL_1099;
  assign _EVAL_2926 = _EVAL_2985 ? _EVAL_826 : _EVAL_2672;
  assign _EVAL_860 = 10'h4a == _EVAL_2998;
  assign _EVAL_215 = _EVAL_726 | gateways_gateway_56__EVAL_4;
  assign fanin__EVAL_11 = _EVAL_3013;
  assign _EVAL_1089 = _EVAL_3236 ? _EVAL_826 : _EVAL_1711;
  assign gateways_gateway_31__EVAL = _EVAL_51;
  assign out_back__EVAL_8 = _EVAL_136;
  assign gateways_gateway_36__EVAL = _EVAL_59;
  assign fanin__EVAL_97 = _EVAL_1283;
  assign _EVAL_2557 = 10'hf == _EVAL_2998;
  assign _EVAL_3336 = {_EVAL_445,_EVAL_2121,_EVAL_3850,_EVAL_3654};
  assign _EVAL_997 = 10'h12 == _EVAL_2998;
  assign _EVAL_2415 = _EVAL_3349[89];
  assign _EVAL_421 = _EVAL_195 & _EVAL_844;
  assign _EVAL_2911 = _EVAL_801 | gateways_gateway_51__EVAL_4;
  assign fanin__EVAL_55 = _EVAL_1268;
  assign _EVAL_3114 = _EVAL_195 & _EVAL_403;
  assign _EVAL_2023 = out_back__EVAL_3[2];
  assign _EVAL_367 = out_back__EVAL;
  assign gateways_gateway_92__EVAL = _EVAL_123;
  assign _EVAL_379 = _EVAL_651[258];
  assign fanin__EVAL_113 = _EVAL_953;
  assign _EVAL_1052 = 10'h75 == _EVAL_2998;
  assign _EVAL_1912 = 10'h42 == _EVAL_2998;
  assign gateways_gateway_106__EVAL = _EVAL_89;
  assign _EVAL_2978 = _EVAL_3704 | gateways_gateway_34__EVAL_4;
  assign gateways_gateway_59__EVAL = _EVAL_8;
  assign _EVAL_3256 = 10'h16 == _EVAL_2998;
  assign _EVAL_1718 = _EVAL_195 & _EVAL_3852;
  assign _EVAL_2963 = _EVAL_3358 & _EVAL_2035;
  assign gateways_gateway_64__EVAL_0 = _EVAL_9;
  assign _EVAL_1354 = _EVAL_651[82];
  assign fanin__EVAL_120 = _EVAL_3284;
  assign _EVAL_2774 = _EVAL_906 & _EVAL_2035;
  assign _EVAL_2492 = _EVAL_3760 | gateways_gateway_97__EVAL_4;
  assign _EVAL_435 = ~_EVAL_3760;
  assign fanin__EVAL_5 = _EVAL_1293;
  assign _EVAL_505 = ~_EVAL_820;
  assign _EVAL_994 = 10'h11 == _EVAL_2998;
  assign gateways_gateway_44__EVAL_0 = _EVAL_9;
  assign gateways_gateway_57__EVAL_3 = _EVAL_110;
  assign _EVAL_2733 = _EVAL_651[26];
  assign _EVAL_3097 = _EVAL_353 & _EVAL_2035;
  assign gateways_gateway_76__EVAL = _EVAL_67;
  assign _EVAL_3287 = _EVAL_651[54];
  assign gateways_gateway_71__EVAL = _EVAL_87;
  assign gateways_gateway_124__EVAL = _EVAL_91;
  assign _EVAL_532 = _EVAL_1506 ? {{29'd0}, _EVAL_1647} : _EVAL_1608;
  assign _EVAL_2019 = 10'hc == _EVAL_2998;
  assign _EVAL_1263 = _EVAL_2593 & _EVAL_2035;
  assign _EVAL_2119 = _EVAL_3189 & _EVAL_2035;
  assign _EVAL_1343 = _EVAL_195 & _EVAL_3618;
  assign _EVAL_2763 = _EVAL_171 ? _EVAL_826 : _EVAL_2861;
  assign _EVAL_3672 = _EVAL_651[55];
  assign _EVAL_1122 = _EVAL_3349[29];
  assign _EVAL_3167 = _EVAL_651[86];
  assign _EVAL_630 = ~_EVAL_3849;
  assign _EVAL_1822 = _EVAL_955 ? _EVAL_826 : _EVAL_1962;
  assign _EVAL_2444 = ~_EVAL_3039;
  assign _EVAL_2133 = _EVAL_1040 & _EVAL_826;
  assign _EVAL_1799 = 10'h4d == _EVAL_2998;
  assign _EVAL_1884 = 10'h29 == _EVAL_2998;
  assign _EVAL_2490 = out_back__EVAL_3[6];
  assign _EVAL_2469 = {_EVAL_1710,_EVAL_1147,_EVAL_1417,_EVAL_2178,_EVAL_2655,_EVAL_668,_EVAL_2167,_EVAL_965,_EVAL_3412,
    _EVAL_3240};
  assign gateways_gateway_110__EVAL_1 = ~_EVAL_3589;
  assign _EVAL_3521 = _EVAL_605 | gateways_gateway_62__EVAL_4;
  always @(posedge _EVAL_9) begin
    if (_EVAL_1729) begin
      _EVAL_167 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_168 <= 1'h0;
    end else if (_EVAL_2090) begin
      _EVAL_168 <= _EVAL_1510;
    end
    if (_EVAL_1662) begin
      _EVAL_172 <= _EVAL_810;
    end
    if (_EVAL_1476) begin
      _EVAL_189 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_193 <= 1'h0;
    end else if (_EVAL_344) begin
      _EVAL_193 <= _EVAL_3794;
    end
    if (_EVAL_110) begin
      _EVAL_202 <= 1'h0;
    end else if (_EVAL_1336) begin
      _EVAL_202 <= _EVAL_1349;
    end
    if (_EVAL_489) begin
      _EVAL_222 <= _EVAL_810;
    end
    if (_EVAL_300) begin
      _EVAL_240 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_276 <= 1'h0;
    end else if (_EVAL_1689) begin
      _EVAL_276 <= _EVAL_2732;
    end
    if (_EVAL_110) begin
      _EVAL_284 <= 1'h0;
    end else if (_EVAL_2730) begin
      _EVAL_284 <= _EVAL_3485;
    end
    if (_EVAL_288) begin
      _EVAL_289 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_302 <= 1'h0;
    end else if (_EVAL_2263) begin
      _EVAL_302 <= _EVAL_1489;
    end
    if (_EVAL_110) begin
      _EVAL_325 <= 1'h0;
    end else if (_EVAL_2492) begin
      _EVAL_325 <= _EVAL_435;
    end
    if (_EVAL_110) begin
      _EVAL_350 <= 1'h0;
    end else if (_EVAL_3261) begin
      _EVAL_350 <= _EVAL_962;
    end
    if (_EVAL_2773) begin
      _EVAL_355 <= _EVAL_810;
    end
    if (_EVAL_1755) begin
      _EVAL_394 <= _EVAL_3265;
    end
    if (_EVAL_110) begin
      _EVAL_414 <= 1'h0;
    end else if (_EVAL_1754) begin
      _EVAL_414 <= _EVAL_3285;
    end
    if (_EVAL_110) begin
      _EVAL_415 <= 1'h0;
    end else if (_EVAL_1657) begin
      _EVAL_415 <= _EVAL_3457;
    end
    if (_EVAL_110) begin
      _EVAL_423 <= 1'h0;
    end else if (_EVAL_215) begin
      _EVAL_423 <= _EVAL_1815;
    end
    if (_EVAL_3339) begin
      _EVAL_445 <= _EVAL_3245;
    end
    if (_EVAL_2206) begin
      _EVAL_456 <= _EVAL_810;
    end
    if (_EVAL_871) begin
      _EVAL_461 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_498 <= 1'h0;
    end else if (_EVAL_2777) begin
      _EVAL_498 <= _EVAL_322;
    end
    if (_EVAL_3519) begin
      _EVAL_513 <= _EVAL_810;
    end
    if (_EVAL_2119) begin
      _EVAL_517 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_526 <= 1'h0;
    end else if (_EVAL_3845) begin
      _EVAL_526 <= _EVAL_390;
    end
    if (_EVAL_110) begin
      _EVAL_552 <= 1'h0;
    end else if (_EVAL_989) begin
      _EVAL_552 <= _EVAL_609;
    end
    if (_EVAL_3390) begin
      _EVAL_570 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_594 <= 1'h0;
    end else if (_EVAL_1209) begin
      _EVAL_594 <= _EVAL_3260;
    end
    if (_EVAL_110) begin
      _EVAL_612 <= 1'h0;
    end else if (_EVAL_2542) begin
      _EVAL_612 <= _EVAL_1061;
    end
    if (_EVAL_715) begin
      _EVAL_628 <= _EVAL_810;
    end
    if (_EVAL_205) begin
      _EVAL_642 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_668 <= 1'h0;
    end else if (_EVAL_1564) begin
      _EVAL_668 <= _EVAL_2159;
    end
    if (_EVAL_110) begin
      _EVAL_677 <= 1'h0;
    end else if (_EVAL_2978) begin
      _EVAL_677 <= _EVAL_639;
    end
    if (_EVAL_2774) begin
      _EVAL_692 <= _EVAL_810;
    end
    if (_EVAL_356) begin
      _EVAL_700 <= _EVAL_810;
    end
    if (_EVAL_1886) begin
      _EVAL_707 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_727 <= 1'h0;
    end else if (_EVAL_3686) begin
      _EVAL_727 <= _EVAL_3303;
    end
    if (_EVAL_110) begin
      _EVAL_744 <= 1'h0;
    end else if (_EVAL_2134) begin
      _EVAL_744 <= _EVAL_703;
    end
    if (_EVAL_110) begin
      _EVAL_770 <= 1'h0;
    end else if (_EVAL_2928) begin
      _EVAL_770 <= _EVAL_2350;
    end
    if (_EVAL_1022) begin
      _EVAL_778 <= _EVAL_810;
    end
    if (_EVAL_2511) begin
      _EVAL_779 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_780 <= 1'h0;
    end else if (_EVAL_1182) begin
      _EVAL_780 <= _EVAL_2779;
    end
    if (_EVAL_3182) begin
      _EVAL_797 <= _EVAL_810;
    end
    _EVAL_809 <= fanin__EVAL_65;
    if (_EVAL_110) begin
      _EVAL_811 <= 1'h0;
    end else if (_EVAL_1195) begin
      _EVAL_811 <= _EVAL_2601;
    end
    if (_EVAL_110) begin
      _EVAL_813 <= 1'h0;
    end else if (_EVAL_3742) begin
      _EVAL_813 <= _EVAL_278;
    end
    if (_EVAL_110) begin
      _EVAL_819 <= 1'h0;
    end else if (_EVAL_1015) begin
      _EVAL_819 <= _EVAL_2530;
    end
    if (_EVAL_151) begin
      _EVAL_853 <= _EVAL_810;
    end
    if (_EVAL_2615) begin
      _EVAL_854 <= _EVAL_810;
    end
    if (_EVAL_3745) begin
      _EVAL_865 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_872 <= 1'h0;
    end else if (_EVAL_1148) begin
      _EVAL_872 <= _EVAL_804;
    end
    if (_EVAL_110) begin
      _EVAL_902 <= 1'h0;
    end else if (_EVAL_1833) begin
      _EVAL_902 <= _EVAL_3663;
    end
    if (_EVAL_110) begin
      _EVAL_911 <= 1'h0;
    end else if (_EVAL_3162) begin
      _EVAL_911 <= _EVAL_793;
    end
    if (_EVAL_2494) begin
      _EVAL_930 <= _EVAL_3265;
    end
    if (_EVAL_687) begin
      _EVAL_936 <= _EVAL_810;
    end
    if (_EVAL_3555) begin
      _EVAL_953 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_965 <= 1'h0;
    end else if (_EVAL_2132) begin
      _EVAL_965 <= _EVAL_3422;
    end
    if (_EVAL_837) begin
      _EVAL_966 <= _EVAL_810;
    end
    if (_EVAL_3735) begin
      _EVAL_1005 <= _EVAL_810;
    end
    if (_EVAL_3408) begin
      _EVAL_1030 <= _EVAL_3245;
    end
    if (_EVAL_2919) begin
      _EVAL_1085 <= _EVAL_810;
    end
    if (_EVAL_2952) begin
      _EVAL_1099 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_1116 <= 1'h0;
    end else if (_EVAL_2832) begin
      _EVAL_1116 <= _EVAL_890;
    end
    if (_EVAL_110) begin
      _EVAL_1120 <= 1'h0;
    end else if (_EVAL_1504) begin
      _EVAL_1120 <= _EVAL_685;
    end
    if (_EVAL_110) begin
      _EVAL_1127 <= 1'h0;
    end else if (_EVAL_834) begin
      _EVAL_1127 <= _EVAL_1890;
    end
    if (_EVAL_244) begin
      _EVAL_1134 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_1138 <= 1'h0;
    end else if (_EVAL_3610) begin
      _EVAL_1138 <= _EVAL_973;
    end
    if (_EVAL_110) begin
      _EVAL_1147 <= 1'h0;
    end else if (_EVAL_1853) begin
      _EVAL_1147 <= _EVAL_641;
    end
    if (_EVAL_110) begin
      _EVAL_1175 <= 1'h0;
    end else if (_EVAL_2896) begin
      _EVAL_1175 <= _EVAL_3316;
    end
    if (_EVAL_2318) begin
      _EVAL_1199 <= _EVAL_810;
    end
    if (_EVAL_2846) begin
      _EVAL_1252 <= _EVAL_810;
    end
    if (_EVAL_2658) begin
      _EVAL_1268 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_1270 <= 1'h0;
    end else if (_EVAL_2043) begin
      _EVAL_1270 <= _EVAL_2399;
    end
    if (_EVAL_2142) begin
      _EVAL_1283 <= _EVAL_810;
    end
    if (_EVAL_223) begin
      _EVAL_1293 <= _EVAL_810;
    end
    if (_EVAL_510) begin
      _EVAL_1340 <= _EVAL_3245;
    end
    if (_EVAL_1905) begin
      _EVAL_1341 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_1347 <= 1'h0;
    end else if (_EVAL_2556) begin
      _EVAL_1347 <= _EVAL_1954;
    end
    if (_EVAL_2734) begin
      _EVAL_1358 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_1365 <= 1'h0;
    end else if (_EVAL_247) begin
      _EVAL_1365 <= _EVAL_3642;
    end
    if (_EVAL_110) begin
      _EVAL_1368 <= 1'h0;
    end else if (_EVAL_1624) begin
      _EVAL_1368 <= _EVAL_1447;
    end
    if (_EVAL_110) begin
      _EVAL_1369 <= 1'h0;
    end else if (_EVAL_2770) begin
      _EVAL_1369 <= _EVAL_889;
    end
    if (_EVAL_1539) begin
      _EVAL_1380 <= _EVAL_2379;
    end
    if (_EVAL_110) begin
      _EVAL_1392 <= 1'h0;
    end else if (_EVAL_490) begin
      _EVAL_1392 <= _EVAL_1010;
    end
    if (_EVAL_2362) begin
      _EVAL_1407 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_1417 <= 1'h0;
    end else if (_EVAL_2700) begin
      _EVAL_1417 <= _EVAL_3183;
    end
    if (_EVAL_110) begin
      _EVAL_1434 <= 1'h0;
    end else if (_EVAL_1520) begin
      _EVAL_1434 <= _EVAL_630;
    end
    if (_EVAL_2661) begin
      _EVAL_1459 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_1467 <= 1'h0;
    end else if (_EVAL_933) begin
      _EVAL_1467 <= _EVAL_848;
    end
    if (_EVAL_772) begin
      _EVAL_1471 <= _EVAL_3245;
    end
    if (_EVAL_110) begin
      _EVAL_1507 <= 1'h0;
    end else if (_EVAL_3632) begin
      _EVAL_1507 <= _EVAL_1907;
    end
    if (_EVAL_1426) begin
      _EVAL_1517 <= _EVAL_2745;
    end
    if (_EVAL_110) begin
      _EVAL_1524 <= 1'h0;
    end else if (_EVAL_343) begin
      _EVAL_1524 <= _EVAL_3639;
    end
    if (_EVAL_1328) begin
      _EVAL_1527 <= _EVAL_810;
    end
    if (_EVAL_2097) begin
      _EVAL_1528 <= _EVAL_810;
    end
    if (_EVAL_1769) begin
      _EVAL_1548 <= _EVAL_2379;
    end
    if (_EVAL_110) begin
      _EVAL_1565 <= 1'h0;
    end else if (_EVAL_2148) begin
      _EVAL_1565 <= _EVAL_3324;
    end
    if (_EVAL_2990) begin
      _EVAL_1569 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_1576 <= 1'h0;
    end else if (_EVAL_2348) begin
      _EVAL_1576 <= _EVAL_1422;
    end
    if (_EVAL_862) begin
      _EVAL_1621 <= _EVAL_810;
    end
    if (_EVAL_1972) begin
      _EVAL_1634 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_1638 <= 1'h0;
    end else if (_EVAL_721) begin
      _EVAL_1638 <= _EVAL_719;
    end
    if (_EVAL_652) begin
      _EVAL_1647 <= _EVAL_810;
    end
    if (_EVAL_1535) begin
      _EVAL_1655 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_1673 <= 1'h0;
    end else if (_EVAL_280) begin
      _EVAL_1673 <= _EVAL_3626;
    end
    if (_EVAL_3068) begin
      _EVAL_1687 <= _EVAL_810;
    end
    if (_EVAL_1164) begin
      _EVAL_1692 <= _EVAL_810;
    end
    if (_EVAL_3179) begin
      _EVAL_1695 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_1710 <= 1'h0;
    end else if (_EVAL_2392) begin
      _EVAL_1710 <= _EVAL_3793;
    end
    if (_EVAL_3097) begin
      _EVAL_1745 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_1749 <= 1'h0;
    end else if (_EVAL_219) begin
      _EVAL_1749 <= _EVAL_3595;
    end
    if (_EVAL_1250) begin
      _EVAL_1758 <= _EVAL_810;
    end
    if (_EVAL_2651) begin
      _EVAL_1771 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_1774 <= 1'h0;
    end else if (_EVAL_3593) begin
      _EVAL_1774 <= _EVAL_603;
    end
    if (_EVAL_917) begin
      _EVAL_1789 <= _EVAL_810;
    end
    if (_EVAL_2270) begin
      _EVAL_1796 <= _EVAL_810;
    end
    if (_EVAL_1320) begin
      _EVAL_1805 <= _EVAL_810;
    end
    if (_EVAL_2054) begin
      _EVAL_1843 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_1847 <= 1'h0;
    end else if (_EVAL_2453) begin
      _EVAL_1847 <= _EVAL_918;
    end
    if (_EVAL_110) begin
      _EVAL_1872 <= 1'h0;
    end else if (_EVAL_2064) begin
      _EVAL_1872 <= _EVAL_3035;
    end
    if (_EVAL_533) begin
      _EVAL_1876 <= _EVAL_810;
    end
    if (_EVAL_765) begin
      _EVAL_1925 <= _EVAL_2697;
    end
    if (_EVAL_110) begin
      _EVAL_1928 <= 1'h0;
    end else if (_EVAL_1359) begin
      _EVAL_1928 <= _EVAL_3844;
    end
    if (_EVAL_110) begin
      _EVAL_1937 <= 1'h0;
    end else if (_EVAL_827) begin
      _EVAL_1937 <= _EVAL_231;
    end
    if (_EVAL_110) begin
      _EVAL_1944 <= 1'h0;
    end else if (_EVAL_2479) begin
      _EVAL_1944 <= _EVAL_1031;
    end
    if (_EVAL_110) begin
      _EVAL_1948 <= 1'h0;
    end else if (_EVAL_3683) begin
      _EVAL_1948 <= _EVAL_567;
    end
    if (_EVAL_2328) begin
      _EVAL_1963 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_1964 <= 1'h0;
    end else if (_EVAL_3777) begin
      _EVAL_1964 <= _EVAL_3376;
    end
    if (_EVAL_3443) begin
      _EVAL_1968 <= _EVAL_810;
    end
    if (_EVAL_2327) begin
      _EVAL_1988 <= _EVAL_810;
    end
    if (_EVAL_3008) begin
      _EVAL_2004 <= _EVAL_810;
    end
    if (_EVAL_1103) begin
      _EVAL_2012 <= _EVAL_810;
    end
    if (_EVAL_3056) begin
      _EVAL_2030 <= _EVAL_810;
    end
    if (_EVAL_1750) begin
      _EVAL_2070 <= _EVAL_2379;
    end
    if (_EVAL_1301) begin
      _EVAL_2079 <= _EVAL_810;
    end
    if (_EVAL_2403) begin
      _EVAL_2121 <= _EVAL_2379;
    end
    if (_EVAL_110) begin
      _EVAL_2143 <= 1'h0;
    end else if (_EVAL_1382) begin
      _EVAL_2143 <= _EVAL_462;
    end
    if (_EVAL_110) begin
      _EVAL_2153 <= 1'h0;
    end else if (_EVAL_1832) begin
      _EVAL_2153 <= _EVAL_1985;
    end
    if (_EVAL_110) begin
      _EVAL_2160 <= 1'h0;
    end else if (_EVAL_3483) begin
      _EVAL_2160 <= _EVAL_2369;
    end
    if (_EVAL_110) begin
      _EVAL_2165 <= 1'h0;
    end else if (_EVAL_3317) begin
      _EVAL_2165 <= _EVAL_783;
    end
    if (_EVAL_110) begin
      _EVAL_2167 <= 1'h0;
    end else if (_EVAL_1773) begin
      _EVAL_2167 <= _EVAL_3791;
    end
    if (_EVAL_110) begin
      _EVAL_2174 <= 1'h0;
    end else if (_EVAL_855) begin
      _EVAL_2174 <= _EVAL_937;
    end
    if (_EVAL_110) begin
      _EVAL_2178 <= 1'h0;
    end else if (_EVAL_2888) begin
      _EVAL_2178 <= _EVAL_1855;
    end
    if (_EVAL_1521) begin
      _EVAL_2182 <= _EVAL_810;
    end
    if (_EVAL_1051) begin
      _EVAL_2186 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_2193 <= 1'h0;
    end else if (_EVAL_899) begin
      _EVAL_2193 <= _EVAL_1783;
    end
    if (_EVAL_110) begin
      _EVAL_2197 <= 1'h0;
    end else if (_EVAL_3531) begin
      _EVAL_2197 <= _EVAL_1222;
    end
    if (_EVAL_259) begin
      _EVAL_2211 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_2221 <= 1'h0;
    end else if (_EVAL_3576) begin
      _EVAL_2221 <= _EVAL_755;
    end
    if (_EVAL_1591) begin
      _EVAL_2262 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_2268 <= 1'h0;
    end else if (_EVAL_2629) begin
      _EVAL_2268 <= _EVAL_3685;
    end
    if (_EVAL_908) begin
      _EVAL_2281 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_2297 <= 1'h0;
    end else if (_EVAL_3851) begin
      _EVAL_2297 <= _EVAL_2460;
    end
    if (_EVAL_575) begin
      _EVAL_2306 <= _EVAL_810;
    end
    if (_EVAL_1720) begin
      _EVAL_2309 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_2344 <= 1'h0;
    end else if (_EVAL_534) begin
      _EVAL_2344 <= _EVAL_1366;
    end
    if (_EVAL_110) begin
      _EVAL_2370 <= 1'h0;
    end else if (_EVAL_2910) begin
      _EVAL_2370 <= _EVAL_3304;
    end
    if (_EVAL_2015) begin
      _EVAL_2384 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_2396 <= 1'h0;
    end else if (_EVAL_787) begin
      _EVAL_2396 <= _EVAL_1957;
    end
    if (_EVAL_3809) begin
      _EVAL_2418 <= _EVAL_3265;
    end
    if (_EVAL_110) begin
      _EVAL_2427 <= 1'h0;
    end else if (_EVAL_1698) begin
      _EVAL_2427 <= _EVAL_228;
    end
    if (_EVAL_2499) begin
      _EVAL_2466 <= _EVAL_810;
    end
    if (_EVAL_2425) begin
      _EVAL_2477 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_2488 <= 1'h0;
    end else if (_EVAL_2833) begin
      _EVAL_2488 <= _EVAL_995;
    end
    if (_EVAL_110) begin
      _EVAL_2502 <= 1'h0;
    end else if (_EVAL_2315) begin
      _EVAL_2502 <= _EVAL_2966;
    end
    if (_EVAL_110) begin
      _EVAL_2509 <= 1'h0;
    end else if (_EVAL_254) begin
      _EVAL_2509 <= _EVAL_2253;
    end
    if (_EVAL_2577) begin
      _EVAL_2518 <= _EVAL_810;
    end
    if (_EVAL_2454) begin
      _EVAL_2531 <= _EVAL_810;
    end
    if (_EVAL_613) begin
      _EVAL_2575 <= _EVAL_810;
    end
    if (_EVAL_3720) begin
      _EVAL_2580 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_2618 <= 1'h0;
    end else if (_EVAL_2289) begin
      _EVAL_2618 <= _EVAL_992;
    end
    if (_EVAL_3662) begin
      _EVAL_2621 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_2627 <= 1'h0;
    end else if (_EVAL_653) begin
      _EVAL_2627 <= _EVAL_3027;
    end
    if (_EVAL_868) begin
      _EVAL_2637 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_2655 <= 1'h0;
    end else if (_EVAL_967) begin
      _EVAL_2655 <= _EVAL_762;
    end
    if (_EVAL_110) begin
      _EVAL_2668 <= 1'h0;
    end else if (_EVAL_3486) begin
      _EVAL_2668 <= _EVAL_1969;
    end
    if (_EVAL_110) begin
      _EVAL_2682 <= 1'h0;
    end else if (_EVAL_3354) begin
      _EVAL_2682 <= _EVAL_505;
    end
    if (_EVAL_110) begin
      _EVAL_2685 <= 1'h0;
    end else if (_EVAL_2439) begin
      _EVAL_2685 <= _EVAL_3353;
    end
    if (_EVAL_110) begin
      _EVAL_2698 <= 1'h0;
    end else if (_EVAL_466) begin
      _EVAL_2698 <= _EVAL_1903;
    end
    if (_EVAL_2756) begin
      _EVAL_2711 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_2719 <= 1'h0;
    end else if (_EVAL_253) begin
      _EVAL_2719 <= _EVAL_2431;
    end
    if (_EVAL_110) begin
      _EVAL_2737 <= 1'h0;
    end else if (_EVAL_1785) begin
      _EVAL_2737 <= _EVAL_2701;
    end
    if (_EVAL_335) begin
      _EVAL_2753 <= _EVAL_810;
    end
    _EVAL_2757 <= fanin__EVAL_86;
    if (_EVAL_110) begin
      _EVAL_2793 <= 1'h0;
    end else if (_EVAL_458) begin
      _EVAL_2793 <= _EVAL_2276;
    end
    if (_EVAL_110) begin
      _EVAL_2799 <= 1'h0;
    end else if (_EVAL_907) begin
      _EVAL_2799 <= _EVAL_1555;
    end
    if (_EVAL_1263) begin
      _EVAL_2828 <= _EVAL_810;
    end
    if (_EVAL_1218) begin
      _EVAL_2845 <= _EVAL_810;
    end
    if (_EVAL_723) begin
      _EVAL_2853 <= _EVAL_810;
    end
    if (_EVAL_2329) begin
      _EVAL_2873 <= _EVAL_810;
    end
    if (_EVAL_1146) begin
      _EVAL_2877 <= _EVAL_2745;
    end
    if (_EVAL_632) begin
      _EVAL_2878 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_2900 <= 1'h0;
    end else if (_EVAL_1733) begin
      _EVAL_2900 <= _EVAL_371;
    end
    if (_EVAL_1953) begin
      _EVAL_2921 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_2944 <= 1'h0;
    end else if (_EVAL_148) begin
      _EVAL_2944 <= _EVAL_2444;
    end
    if (_EVAL_110) begin
      _EVAL_2951 <= 1'h0;
    end else if (_EVAL_3264) begin
      _EVAL_2951 <= _EVAL_2083;
    end
    if (_EVAL_110) begin
      _EVAL_2961 <= 1'h0;
    end else if (_EVAL_383) begin
      _EVAL_2961 <= _EVAL_2130;
    end
    if (_EVAL_1715) begin
      _EVAL_2981 <= _EVAL_810;
    end
    if (_EVAL_851) begin
      _EVAL_2982 <= _EVAL_810;
    end
    if (_EVAL_275) begin
      _EVAL_2986 <= _EVAL_810;
    end
    if (_EVAL_3715) begin
      _EVAL_2988 <= _EVAL_810;
    end
    if (_EVAL_1613) begin
      _EVAL_2996 <= _EVAL_810;
    end
    if (_EVAL_604) begin
      _EVAL_3005 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_3011 <= 1'h0;
    end else if (_EVAL_2913) begin
      _EVAL_3011 <= _EVAL_710;
    end
    if (_EVAL_3410) begin
      _EVAL_3013 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_3014 <= 1'h0;
    end else if (_EVAL_2911) begin
      _EVAL_3014 <= _EVAL_1020;
    end
    if (_EVAL_110) begin
      _EVAL_3043 <= 1'h0;
    end else if (_EVAL_1658) begin
      _EVAL_3043 <= _EVAL_944;
    end
    if (_EVAL_3286) begin
      _EVAL_3055 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_3059 <= 1'h0;
    end else if (_EVAL_1024) begin
      _EVAL_3059 <= _EVAL_585;
    end
    if (_EVAL_590) begin
      _EVAL_3063 <= _EVAL_810;
    end
    if (_EVAL_2198) begin
      _EVAL_3072 <= _EVAL_810;
    end
    if (_EVAL_3787) begin
      _EVAL_3080 <= _EVAL_810;
    end
    if (_EVAL_1401) begin
      _EVAL_3096 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_3107 <= 1'h0;
    end else if (_EVAL_1364) begin
      _EVAL_3107 <= _EVAL_1674;
    end
    if (_EVAL_110) begin
      _EVAL_3112 <= 1'h0;
    end else if (_EVAL_2345) begin
      _EVAL_3112 <= _EVAL_2028;
    end
    if (_EVAL_110) begin
      _EVAL_3129 <= 1'h0;
    end else if (_EVAL_2337) begin
      _EVAL_3129 <= _EVAL_2106;
    end
    if (_EVAL_110) begin
      _EVAL_3140 <= 1'h0;
    end else if (_EVAL_3807) begin
      _EVAL_3140 <= _EVAL_1314;
    end
    if (_EVAL_110) begin
      _EVAL_3145 <= 1'h0;
    end else if (_EVAL_1153) begin
      _EVAL_3145 <= _EVAL_3210;
    end
    if (_EVAL_110) begin
      _EVAL_3150 <= 1'h0;
    end else if (_EVAL_2649) begin
      _EVAL_3150 <= _EVAL_679;
    end
    if (_EVAL_110) begin
      _EVAL_3151 <= 1'h0;
    end else if (_EVAL_2122) begin
      _EVAL_3151 <= _EVAL_3061;
    end
    if (_EVAL_320) begin
      _EVAL_3156 <= _EVAL_810;
    end
    if (_EVAL_485) begin
      _EVAL_3191 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_3199 <= 1'h0;
    end else if (_EVAL_156) begin
      _EVAL_3199 <= _EVAL_2805;
    end
    if (_EVAL_110) begin
      _EVAL_3200 <= 1'h0;
    end else if (_EVAL_1023) begin
      _EVAL_3200 <= _EVAL_1549;
    end
    if (_EVAL_110) begin
      _EVAL_3213 <= 1'h0;
    end else if (_EVAL_3002) begin
      _EVAL_3213 <= _EVAL_3106;
    end
    if (_EVAL_1267) begin
      _EVAL_3216 <= _EVAL_810;
    end
    if (_EVAL_2689) begin
      _EVAL_3218 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_3242 <= 1'h0;
    end else if (_EVAL_331) begin
      _EVAL_3242 <= _EVAL_2483;
    end
    if (_EVAL_110) begin
      _EVAL_3268 <= 1'h0;
    end else if (_EVAL_2380) begin
      _EVAL_3268 <= _EVAL_2787;
    end
    if (_EVAL_2963) begin
      _EVAL_3284 <= _EVAL_810;
    end
    if (_EVAL_1896) begin
      _EVAL_3290 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_3305 <= 1'h0;
    end else if (_EVAL_270) begin
      _EVAL_3305 <= _EVAL_495;
    end
    if (_EVAL_3719) begin
      _EVAL_3315 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_3331 <= 1'h0;
    end else if (_EVAL_1752) begin
      _EVAL_3331 <= _EVAL_688;
    end
    if (_EVAL_1202) begin
      _EVAL_3342 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_3346 <= 1'h0;
    end else if (_EVAL_607) begin
      _EVAL_3346 <= _EVAL_1536;
    end
    if (_EVAL_3494) begin
      _EVAL_3357 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_3366 <= 1'h0;
    end else if (_EVAL_2915) begin
      _EVAL_3366 <= _EVAL_3436;
    end
    if (_EVAL_110) begin
      _EVAL_3387 <= 1'h0;
    end else if (_EVAL_1684) begin
      _EVAL_3387 <= _EVAL_2231;
    end
    if (_EVAL_110) begin
      _EVAL_3395 <= 1'h0;
    end else if (_EVAL_2667) begin
      _EVAL_3395 <= _EVAL_759;
    end
    if (_EVAL_110) begin
      _EVAL_3420 <= 1'h0;
    end else if (_EVAL_3521) begin
      _EVAL_3420 <= _EVAL_712;
    end
    if (_EVAL_3064) begin
      _EVAL_3437 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_3440 <= 1'h0;
    end else if (_EVAL_177) begin
      _EVAL_3440 <= _EVAL_2294;
    end
    if (_EVAL_2113) begin
      _EVAL_3446 <= _EVAL_810;
    end
    if (_EVAL_2410) begin
      _EVAL_3469 <= _EVAL_810;
    end
    if (_EVAL_2190) begin
      _EVAL_3505 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_3508 <= 1'h0;
    end else if (_EVAL_1473) begin
      _EVAL_3508 <= _EVAL_1286;
    end
    if (_EVAL_799) begin
      _EVAL_3513 <= _EVAL_810;
    end
    if (_EVAL_777) begin
      _EVAL_3516 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_3527 <= 1'h0;
    end else if (_EVAL_480) begin
      _EVAL_3527 <= _EVAL_771;
    end
    if (_EVAL_3321) begin
      _EVAL_3559 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_3589 <= 1'h0;
    end else if (_EVAL_3530) begin
      _EVAL_3589 <= _EVAL_1257;
    end
    if (_EVAL_180) begin
      _EVAL_3590 <= _EVAL_810;
    end
    if (_EVAL_3840) begin
      _EVAL_3624 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_3627 <= 1'h0;
    end else if (_EVAL_1339) begin
      _EVAL_3627 <= _EVAL_296;
    end
    if (_EVAL_1664) begin
      _EVAL_3635 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_3643 <= 1'h0;
    end else if (_EVAL_3155) begin
      _EVAL_3643 <= _EVAL_2145;
    end
    if (_EVAL_2011) begin
      _EVAL_3653 <= _EVAL_810;
    end
    if (_EVAL_3359) begin
      _EVAL_3654 <= _EVAL_2745;
    end
    if (_EVAL_110) begin
      _EVAL_3656 <= 1'h0;
    end else if (_EVAL_610) begin
      _EVAL_3656 <= _EVAL_2498;
    end
    if (_EVAL_1596) begin
      _EVAL_3657 <= _EVAL_810;
    end
    if (_EVAL_1904) begin
      _EVAL_3711 <= _EVAL_810;
    end
    if (_EVAL_333) begin
      _EVAL_3734 <= _EVAL_810;
    end
    if (_EVAL_1797) begin
      _EVAL_3737 <= _EVAL_810;
    end
    if (_EVAL_509) begin
      _EVAL_3744 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_3770 <= 1'h0;
    end else if (_EVAL_1255) begin
      _EVAL_3770 <= _EVAL_1792;
    end
    if (_EVAL_796) begin
      _EVAL_3798 <= _EVAL_810;
    end
    if (_EVAL_110) begin
      _EVAL_3803 <= 1'h0;
    end else if (_EVAL_979) begin
      _EVAL_3803 <= _EVAL_1065;
    end
    if (_EVAL_110) begin
      _EVAL_3824 <= 1'h0;
    end else if (_EVAL_3375) begin
      _EVAL_3824 <= _EVAL_1683;
    end
    if (_EVAL_2087) begin
      _EVAL_3825 <= _EVAL_810;
    end
    if (_EVAL_3722) begin
      _EVAL_3835 <= _EVAL_810;
    end
    if (_EVAL_3347) begin
      _EVAL_3850 <= _EVAL_3265;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_167 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_168 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_172 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_189 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_193 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_202 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_222 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_240 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_276 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_284 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_289 = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_302 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_325 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_350 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_355 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_394 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_414 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _EVAL_415 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _EVAL_423 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  _EVAL_445 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  _EVAL_456 = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  _EVAL_461 = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  _EVAL_498 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  _EVAL_513 = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  _EVAL_517 = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  _EVAL_526 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  _EVAL_552 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  _EVAL_570 = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  _EVAL_594 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  _EVAL_612 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  _EVAL_628 = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  _EVAL_642 = _RAND_31[2:0];
  _RAND_32 = {1{`RANDOM}};
  _EVAL_668 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  _EVAL_677 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  _EVAL_692 = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  _EVAL_700 = _RAND_35[2:0];
  _RAND_36 = {1{`RANDOM}};
  _EVAL_707 = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  _EVAL_727 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  _EVAL_744 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  _EVAL_770 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  _EVAL_778 = _RAND_40[2:0];
  _RAND_41 = {1{`RANDOM}};
  _EVAL_779 = _RAND_41[2:0];
  _RAND_42 = {1{`RANDOM}};
  _EVAL_780 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  _EVAL_797 = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  _EVAL_809 = _RAND_44[2:0];
  _RAND_45 = {1{`RANDOM}};
  _EVAL_811 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  _EVAL_813 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  _EVAL_819 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  _EVAL_853 = _RAND_48[2:0];
  _RAND_49 = {1{`RANDOM}};
  _EVAL_854 = _RAND_49[2:0];
  _RAND_50 = {1{`RANDOM}};
  _EVAL_865 = _RAND_50[2:0];
  _RAND_51 = {1{`RANDOM}};
  _EVAL_872 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  _EVAL_902 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  _EVAL_911 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  _EVAL_930 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  _EVAL_936 = _RAND_55[2:0];
  _RAND_56 = {1{`RANDOM}};
  _EVAL_953 = _RAND_56[2:0];
  _RAND_57 = {1{`RANDOM}};
  _EVAL_965 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  _EVAL_966 = _RAND_58[2:0];
  _RAND_59 = {1{`RANDOM}};
  _EVAL_1005 = _RAND_59[2:0];
  _RAND_60 = {1{`RANDOM}};
  _EVAL_1030 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  _EVAL_1085 = _RAND_61[2:0];
  _RAND_62 = {1{`RANDOM}};
  _EVAL_1099 = _RAND_62[2:0];
  _RAND_63 = {1{`RANDOM}};
  _EVAL_1116 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  _EVAL_1120 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  _EVAL_1127 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  _EVAL_1134 = _RAND_66[2:0];
  _RAND_67 = {1{`RANDOM}};
  _EVAL_1138 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  _EVAL_1147 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  _EVAL_1175 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  _EVAL_1199 = _RAND_70[2:0];
  _RAND_71 = {1{`RANDOM}};
  _EVAL_1252 = _RAND_71[2:0];
  _RAND_72 = {1{`RANDOM}};
  _EVAL_1268 = _RAND_72[2:0];
  _RAND_73 = {1{`RANDOM}};
  _EVAL_1270 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  _EVAL_1283 = _RAND_74[2:0];
  _RAND_75 = {1{`RANDOM}};
  _EVAL_1293 = _RAND_75[2:0];
  _RAND_76 = {1{`RANDOM}};
  _EVAL_1340 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  _EVAL_1341 = _RAND_77[2:0];
  _RAND_78 = {1{`RANDOM}};
  _EVAL_1347 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  _EVAL_1358 = _RAND_79[2:0];
  _RAND_80 = {1{`RANDOM}};
  _EVAL_1365 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  _EVAL_1368 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  _EVAL_1369 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  _EVAL_1380 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  _EVAL_1392 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  _EVAL_1407 = _RAND_85[2:0];
  _RAND_86 = {1{`RANDOM}};
  _EVAL_1417 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  _EVAL_1434 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  _EVAL_1459 = _RAND_88[2:0];
  _RAND_89 = {1{`RANDOM}};
  _EVAL_1467 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  _EVAL_1471 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  _EVAL_1507 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  _EVAL_1517 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  _EVAL_1524 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  _EVAL_1527 = _RAND_94[2:0];
  _RAND_95 = {1{`RANDOM}};
  _EVAL_1528 = _RAND_95[2:0];
  _RAND_96 = {1{`RANDOM}};
  _EVAL_1548 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  _EVAL_1565 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  _EVAL_1569 = _RAND_98[2:0];
  _RAND_99 = {1{`RANDOM}};
  _EVAL_1576 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  _EVAL_1621 = _RAND_100[2:0];
  _RAND_101 = {1{`RANDOM}};
  _EVAL_1634 = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  _EVAL_1638 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  _EVAL_1647 = _RAND_103[2:0];
  _RAND_104 = {1{`RANDOM}};
  _EVAL_1655 = _RAND_104[2:0];
  _RAND_105 = {1{`RANDOM}};
  _EVAL_1673 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  _EVAL_1687 = _RAND_106[2:0];
  _RAND_107 = {1{`RANDOM}};
  _EVAL_1692 = _RAND_107[2:0];
  _RAND_108 = {1{`RANDOM}};
  _EVAL_1695 = _RAND_108[2:0];
  _RAND_109 = {1{`RANDOM}};
  _EVAL_1710 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  _EVAL_1745 = _RAND_110[2:0];
  _RAND_111 = {1{`RANDOM}};
  _EVAL_1749 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  _EVAL_1758 = _RAND_112[2:0];
  _RAND_113 = {1{`RANDOM}};
  _EVAL_1771 = _RAND_113[2:0];
  _RAND_114 = {1{`RANDOM}};
  _EVAL_1774 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  _EVAL_1789 = _RAND_115[2:0];
  _RAND_116 = {1{`RANDOM}};
  _EVAL_1796 = _RAND_116[2:0];
  _RAND_117 = {1{`RANDOM}};
  _EVAL_1805 = _RAND_117[2:0];
  _RAND_118 = {1{`RANDOM}};
  _EVAL_1843 = _RAND_118[2:0];
  _RAND_119 = {1{`RANDOM}};
  _EVAL_1847 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  _EVAL_1872 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  _EVAL_1876 = _RAND_121[2:0];
  _RAND_122 = {1{`RANDOM}};
  _EVAL_1925 = _RAND_122[6:0];
  _RAND_123 = {1{`RANDOM}};
  _EVAL_1928 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  _EVAL_1937 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  _EVAL_1944 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  _EVAL_1948 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  _EVAL_1963 = _RAND_127[2:0];
  _RAND_128 = {1{`RANDOM}};
  _EVAL_1964 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  _EVAL_1968 = _RAND_129[2:0];
  _RAND_130 = {1{`RANDOM}};
  _EVAL_1988 = _RAND_130[2:0];
  _RAND_131 = {1{`RANDOM}};
  _EVAL_2004 = _RAND_131[2:0];
  _RAND_132 = {1{`RANDOM}};
  _EVAL_2012 = _RAND_132[2:0];
  _RAND_133 = {1{`RANDOM}};
  _EVAL_2030 = _RAND_133[2:0];
  _RAND_134 = {1{`RANDOM}};
  _EVAL_2070 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  _EVAL_2079 = _RAND_135[2:0];
  _RAND_136 = {1{`RANDOM}};
  _EVAL_2121 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  _EVAL_2143 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  _EVAL_2153 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  _EVAL_2160 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  _EVAL_2165 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  _EVAL_2167 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  _EVAL_2174 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  _EVAL_2178 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  _EVAL_2182 = _RAND_144[2:0];
  _RAND_145 = {1{`RANDOM}};
  _EVAL_2186 = _RAND_145[2:0];
  _RAND_146 = {1{`RANDOM}};
  _EVAL_2193 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  _EVAL_2197 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  _EVAL_2211 = _RAND_148[2:0];
  _RAND_149 = {1{`RANDOM}};
  _EVAL_2221 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  _EVAL_2262 = _RAND_150[2:0];
  _RAND_151 = {1{`RANDOM}};
  _EVAL_2268 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  _EVAL_2281 = _RAND_152[2:0];
  _RAND_153 = {1{`RANDOM}};
  _EVAL_2297 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  _EVAL_2306 = _RAND_154[2:0];
  _RAND_155 = {1{`RANDOM}};
  _EVAL_2309 = _RAND_155[2:0];
  _RAND_156 = {1{`RANDOM}};
  _EVAL_2344 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  _EVAL_2370 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  _EVAL_2384 = _RAND_158[2:0];
  _RAND_159 = {1{`RANDOM}};
  _EVAL_2396 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  _EVAL_2418 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  _EVAL_2427 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  _EVAL_2466 = _RAND_162[2:0];
  _RAND_163 = {1{`RANDOM}};
  _EVAL_2477 = _RAND_163[2:0];
  _RAND_164 = {1{`RANDOM}};
  _EVAL_2488 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  _EVAL_2502 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  _EVAL_2509 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  _EVAL_2518 = _RAND_167[2:0];
  _RAND_168 = {1{`RANDOM}};
  _EVAL_2531 = _RAND_168[2:0];
  _RAND_169 = {1{`RANDOM}};
  _EVAL_2575 = _RAND_169[2:0];
  _RAND_170 = {1{`RANDOM}};
  _EVAL_2580 = _RAND_170[2:0];
  _RAND_171 = {1{`RANDOM}};
  _EVAL_2618 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  _EVAL_2621 = _RAND_172[2:0];
  _RAND_173 = {1{`RANDOM}};
  _EVAL_2627 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  _EVAL_2637 = _RAND_174[2:0];
  _RAND_175 = {1{`RANDOM}};
  _EVAL_2655 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  _EVAL_2668 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  _EVAL_2682 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  _EVAL_2685 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  _EVAL_2698 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  _EVAL_2711 = _RAND_180[2:0];
  _RAND_181 = {1{`RANDOM}};
  _EVAL_2719 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  _EVAL_2737 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  _EVAL_2753 = _RAND_183[2:0];
  _RAND_184 = {1{`RANDOM}};
  _EVAL_2757 = _RAND_184[6:0];
  _RAND_185 = {1{`RANDOM}};
  _EVAL_2793 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  _EVAL_2799 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  _EVAL_2828 = _RAND_187[2:0];
  _RAND_188 = {1{`RANDOM}};
  _EVAL_2845 = _RAND_188[2:0];
  _RAND_189 = {1{`RANDOM}};
  _EVAL_2853 = _RAND_189[2:0];
  _RAND_190 = {1{`RANDOM}};
  _EVAL_2873 = _RAND_190[2:0];
  _RAND_191 = {1{`RANDOM}};
  _EVAL_2877 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  _EVAL_2878 = _RAND_192[2:0];
  _RAND_193 = {1{`RANDOM}};
  _EVAL_2900 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  _EVAL_2921 = _RAND_194[2:0];
  _RAND_195 = {1{`RANDOM}};
  _EVAL_2944 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  _EVAL_2951 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  _EVAL_2961 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  _EVAL_2981 = _RAND_198[2:0];
  _RAND_199 = {1{`RANDOM}};
  _EVAL_2982 = _RAND_199[2:0];
  _RAND_200 = {1{`RANDOM}};
  _EVAL_2986 = _RAND_200[2:0];
  _RAND_201 = {1{`RANDOM}};
  _EVAL_2988 = _RAND_201[2:0];
  _RAND_202 = {1{`RANDOM}};
  _EVAL_2996 = _RAND_202[2:0];
  _RAND_203 = {1{`RANDOM}};
  _EVAL_3005 = _RAND_203[2:0];
  _RAND_204 = {1{`RANDOM}};
  _EVAL_3011 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  _EVAL_3013 = _RAND_205[2:0];
  _RAND_206 = {1{`RANDOM}};
  _EVAL_3014 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  _EVAL_3043 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  _EVAL_3055 = _RAND_208[2:0];
  _RAND_209 = {1{`RANDOM}};
  _EVAL_3059 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  _EVAL_3063 = _RAND_210[2:0];
  _RAND_211 = {1{`RANDOM}};
  _EVAL_3072 = _RAND_211[2:0];
  _RAND_212 = {1{`RANDOM}};
  _EVAL_3080 = _RAND_212[2:0];
  _RAND_213 = {1{`RANDOM}};
  _EVAL_3096 = _RAND_213[2:0];
  _RAND_214 = {1{`RANDOM}};
  _EVAL_3107 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  _EVAL_3112 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  _EVAL_3129 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  _EVAL_3140 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  _EVAL_3145 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  _EVAL_3150 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  _EVAL_3151 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  _EVAL_3156 = _RAND_221[2:0];
  _RAND_222 = {1{`RANDOM}};
  _EVAL_3191 = _RAND_222[2:0];
  _RAND_223 = {1{`RANDOM}};
  _EVAL_3199 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  _EVAL_3200 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  _EVAL_3213 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  _EVAL_3216 = _RAND_226[2:0];
  _RAND_227 = {1{`RANDOM}};
  _EVAL_3218 = _RAND_227[2:0];
  _RAND_228 = {1{`RANDOM}};
  _EVAL_3242 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  _EVAL_3268 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  _EVAL_3284 = _RAND_230[2:0];
  _RAND_231 = {1{`RANDOM}};
  _EVAL_3290 = _RAND_231[2:0];
  _RAND_232 = {1{`RANDOM}};
  _EVAL_3305 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  _EVAL_3315 = _RAND_233[2:0];
  _RAND_234 = {1{`RANDOM}};
  _EVAL_3331 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  _EVAL_3342 = _RAND_235[2:0];
  _RAND_236 = {1{`RANDOM}};
  _EVAL_3346 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  _EVAL_3357 = _RAND_237[2:0];
  _RAND_238 = {1{`RANDOM}};
  _EVAL_3366 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  _EVAL_3387 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  _EVAL_3395 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  _EVAL_3420 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  _EVAL_3437 = _RAND_242[2:0];
  _RAND_243 = {1{`RANDOM}};
  _EVAL_3440 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  _EVAL_3446 = _RAND_244[2:0];
  _RAND_245 = {1{`RANDOM}};
  _EVAL_3469 = _RAND_245[2:0];
  _RAND_246 = {1{`RANDOM}};
  _EVAL_3505 = _RAND_246[2:0];
  _RAND_247 = {1{`RANDOM}};
  _EVAL_3508 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  _EVAL_3513 = _RAND_248[2:0];
  _RAND_249 = {1{`RANDOM}};
  _EVAL_3516 = _RAND_249[2:0];
  _RAND_250 = {1{`RANDOM}};
  _EVAL_3527 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  _EVAL_3559 = _RAND_251[2:0];
  _RAND_252 = {1{`RANDOM}};
  _EVAL_3589 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  _EVAL_3590 = _RAND_253[2:0];
  _RAND_254 = {1{`RANDOM}};
  _EVAL_3624 = _RAND_254[2:0];
  _RAND_255 = {1{`RANDOM}};
  _EVAL_3627 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  _EVAL_3635 = _RAND_256[2:0];
  _RAND_257 = {1{`RANDOM}};
  _EVAL_3643 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  _EVAL_3653 = _RAND_258[2:0];
  _RAND_259 = {1{`RANDOM}};
  _EVAL_3654 = _RAND_259[7:0];
  _RAND_260 = {1{`RANDOM}};
  _EVAL_3656 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  _EVAL_3657 = _RAND_261[2:0];
  _RAND_262 = {1{`RANDOM}};
  _EVAL_3711 = _RAND_262[2:0];
  _RAND_263 = {1{`RANDOM}};
  _EVAL_3734 = _RAND_263[2:0];
  _RAND_264 = {1{`RANDOM}};
  _EVAL_3737 = _RAND_264[2:0];
  _RAND_265 = {1{`RANDOM}};
  _EVAL_3744 = _RAND_265[2:0];
  _RAND_266 = {1{`RANDOM}};
  _EVAL_3770 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  _EVAL_3798 = _RAND_267[2:0];
  _RAND_268 = {1{`RANDOM}};
  _EVAL_3803 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  _EVAL_3824 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  _EVAL_3825 = _RAND_270[2:0];
  _RAND_271 = {1{`RANDOM}};
  _EVAL_3835 = _RAND_271[2:0];
  _RAND_272 = {1{`RANDOM}};
  _EVAL_3850 = _RAND_272[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
