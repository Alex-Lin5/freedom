//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_39(
  output        _EVAL,
  output        _EVAL_0,
  input         _EVAL_1,
  input  [2:0]  _EVAL_2,
  output [31:0] _EVAL_3,
  output [31:0] _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  output        _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  output [31:0] _EVAL_10,
  output        _EVAL_11,
  output [3:0]  _EVAL_12,
  input  [1:0]  _EVAL_13,
  output        _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input  [3:0]  _EVAL_17,
  output [2:0]  _EVAL_18,
  input         _EVAL_19,
  output [2:0]  _EVAL_20,
  input  [31:0] _EVAL_21,
  input  [3:0]  _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  input  [31:0] _EVAL_25,
  output [3:0]  _EVAL_26,
  input  [31:0] _EVAL_27,
  output        _EVAL_28,
  output        _EVAL_29,
  input  [1:0]  _EVAL_30,
  output        _EVAL_31,
  output        _EVAL_32,
  output        _EVAL_33,
  input         _EVAL_34,
  input  [2:0]  _EVAL_35
);
  wire [2:0] fixer__EVAL;
  wire  fixer__EVAL_0;
  wire [2:0] fixer__EVAL_1;
  wire  fixer__EVAL_2;
  wire  fixer__EVAL_3;
  wire  fixer__EVAL_4;
  wire [3:0] fixer__EVAL_5;
  wire [1:0] fixer__EVAL_6;
  wire [3:0] fixer__EVAL_7;
  wire  fixer__EVAL_8;
  wire [3:0] fixer__EVAL_9;
  wire [31:0] fixer__EVAL_10;
  wire  fixer__EVAL_11;
  wire [2:0] fixer__EVAL_12;
  wire  fixer__EVAL_13;
  wire  fixer__EVAL_14;
  wire  fixer__EVAL_15;
  wire [31:0] fixer__EVAL_16;
  wire [3:0] fixer__EVAL_17;
  wire  fixer__EVAL_18;
  wire  fixer__EVAL_19;
  wire  fixer__EVAL_20;
  wire  fixer__EVAL_21;
  wire  fixer__EVAL_22;
  wire [31:0] fixer__EVAL_23;
  wire  fixer__EVAL_24;
  wire [31:0] fixer__EVAL_25;
  wire [31:0] fixer__EVAL_26;
  wire  fixer__EVAL_27;
  wire  fixer__EVAL_28;
  wire  fixer__EVAL_29;
  wire  fixer__EVAL_30;
  wire  fixer__EVAL_31;
  wire  fixer__EVAL_32;
  wire [31:0] fixer__EVAL_33;
  wire  fixer__EVAL_34;
  wire [3:0] fixer__EVAL_35;
  wire  fixer__EVAL_36;
  wire  fixer__EVAL_37;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire [31:0] _EVAL_38;
  wire [3:0] _EVAL_39;
  wire  _EVAL_40;
  wire [3:0] _EVAL_41;
  wire [31:0] _EVAL_42;
  wire [3:0] _EVAL_43;
  wire  _EVAL_44;
  wire [31:0] _EVAL_45;
  wire  _EVAL_46;
  wire [2:0] _EVAL_47;
  wire  _EVAL_48;
  wire [31:0] _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire [31:0] _EVAL_52;
  wire  buffer__EVAL;
  wire [2:0] buffer__EVAL_0;
  wire  buffer__EVAL_1;
  wire  buffer__EVAL_2;
  wire  buffer__EVAL_3;
  wire [2:0] buffer__EVAL_4;
  wire  buffer__EVAL_5;
  wire [31:0] buffer__EVAL_6;
  wire [3:0] buffer__EVAL_7;
  wire  buffer__EVAL_8;
  wire  buffer__EVAL_9;
  wire  buffer__EVAL_10;
  wire  buffer__EVAL_11;
  wire  buffer__EVAL_12;
  wire  buffer__EVAL_13;
  wire  buffer__EVAL_14;
  wire [31:0] buffer__EVAL_15;
  wire [3:0] buffer__EVAL_16;
  wire [2:0] buffer__EVAL_17;
  wire  buffer__EVAL_18;
  wire  buffer__EVAL_19;
  wire  buffer__EVAL_20;
  wire [31:0] buffer__EVAL_21;
  wire [3:0] buffer__EVAL_22;
  wire [2:0] buffer__EVAL_23;
  wire  buffer__EVAL_24;
  wire  buffer__EVAL_25;
  wire [31:0] buffer__EVAL_26;
  wire [31:0] buffer__EVAL_27;
  wire  buffer__EVAL_28;
  wire  buffer__EVAL_29;
  wire  buffer__EVAL_30;
  wire  buffer__EVAL_31;
  wire [1:0] buffer__EVAL_32;
  wire [3:0] buffer__EVAL_33;
  wire [3:0] buffer__EVAL_34;
  wire  buffer__EVAL_35;
  wire  buffer__EVAL_36;
  wire  buffer__EVAL_37;
  wire  buffer__EVAL_38;
  wire  buffer__EVAL_39;
  wire [2:0] buffer__EVAL_40;
  wire [3:0] buffer__EVAL_41;
  wire  buffer__EVAL_42;
  wire [1:0] buffer__EVAL_43;
  wire [31:0] buffer__EVAL_44;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  ahb2tl__EVAL;
  wire [2:0] ahb2tl__EVAL_0;
  wire  ahb2tl__EVAL_1;
  wire  ahb2tl__EVAL_2;
  wire [31:0] ahb2tl__EVAL_3;
  wire [31:0] ahb2tl__EVAL_4;
  wire  ahb2tl__EVAL_5;
  wire  ahb2tl__EVAL_6;
  wire  ahb2tl__EVAL_7;
  wire  ahb2tl__EVAL_8;
  wire  ahb2tl__EVAL_9;
  wire [31:0] ahb2tl__EVAL_10;
  wire  ahb2tl__EVAL_11;
  wire [31:0] ahb2tl__EVAL_12;
  wire [2:0] ahb2tl__EVAL_13;
  wire  ahb2tl__EVAL_14;
  wire [31:0] ahb2tl__EVAL_15;
  wire [3:0] ahb2tl__EVAL_16;
  wire  ahb2tl__EVAL_17;
  wire [3:0] ahb2tl__EVAL_18;
  wire  ahb2tl__EVAL_19;
  wire  ahb2tl__EVAL_20;
  wire  ahb2tl__EVAL_21;
  wire [31:0] ahb2tl__EVAL_22;
  wire [1:0] ahb2tl__EVAL_23;
  wire  ahb2tl__EVAL_24;
  wire  ahb2tl__EVAL_25;
  wire [3:0] ahb2tl__EVAL_26;
  wire  ahb2tl__EVAL_27;
  wire [2:0] ahb2tl__EVAL_28;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire [31:0] _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire [2:0] _EVAL_64;
  wire [3:0] _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  _EVAL_37 fixer (
    ._EVAL(fixer__EVAL),
    ._EVAL_0(fixer__EVAL_0),
    ._EVAL_1(fixer__EVAL_1),
    ._EVAL_2(fixer__EVAL_2),
    ._EVAL_3(fixer__EVAL_3),
    ._EVAL_4(fixer__EVAL_4),
    ._EVAL_5(fixer__EVAL_5),
    ._EVAL_6(fixer__EVAL_6),
    ._EVAL_7(fixer__EVAL_7),
    ._EVAL_8(fixer__EVAL_8),
    ._EVAL_9(fixer__EVAL_9),
    ._EVAL_10(fixer__EVAL_10),
    ._EVAL_11(fixer__EVAL_11),
    ._EVAL_12(fixer__EVAL_12),
    ._EVAL_13(fixer__EVAL_13),
    ._EVAL_14(fixer__EVAL_14),
    ._EVAL_15(fixer__EVAL_15),
    ._EVAL_16(fixer__EVAL_16),
    ._EVAL_17(fixer__EVAL_17),
    ._EVAL_18(fixer__EVAL_18),
    ._EVAL_19(fixer__EVAL_19),
    ._EVAL_20(fixer__EVAL_20),
    ._EVAL_21(fixer__EVAL_21),
    ._EVAL_22(fixer__EVAL_22),
    ._EVAL_23(fixer__EVAL_23),
    ._EVAL_24(fixer__EVAL_24),
    ._EVAL_25(fixer__EVAL_25),
    ._EVAL_26(fixer__EVAL_26),
    ._EVAL_27(fixer__EVAL_27),
    ._EVAL_28(fixer__EVAL_28),
    ._EVAL_29(fixer__EVAL_29),
    ._EVAL_30(fixer__EVAL_30),
    ._EVAL_31(fixer__EVAL_31),
    ._EVAL_32(fixer__EVAL_32),
    ._EVAL_33(fixer__EVAL_33),
    ._EVAL_34(fixer__EVAL_34),
    ._EVAL_35(fixer__EVAL_35),
    ._EVAL_36(fixer__EVAL_36),
    ._EVAL_37(fixer__EVAL_37)
  );
  _EVAL_35 buffer (
    ._EVAL(buffer__EVAL),
    ._EVAL_0(buffer__EVAL_0),
    ._EVAL_1(buffer__EVAL_1),
    ._EVAL_2(buffer__EVAL_2),
    ._EVAL_3(buffer__EVAL_3),
    ._EVAL_4(buffer__EVAL_4),
    ._EVAL_5(buffer__EVAL_5),
    ._EVAL_6(buffer__EVAL_6),
    ._EVAL_7(buffer__EVAL_7),
    ._EVAL_8(buffer__EVAL_8),
    ._EVAL_9(buffer__EVAL_9),
    ._EVAL_10(buffer__EVAL_10),
    ._EVAL_11(buffer__EVAL_11),
    ._EVAL_12(buffer__EVAL_12),
    ._EVAL_13(buffer__EVAL_13),
    ._EVAL_14(buffer__EVAL_14),
    ._EVAL_15(buffer__EVAL_15),
    ._EVAL_16(buffer__EVAL_16),
    ._EVAL_17(buffer__EVAL_17),
    ._EVAL_18(buffer__EVAL_18),
    ._EVAL_19(buffer__EVAL_19),
    ._EVAL_20(buffer__EVAL_20),
    ._EVAL_21(buffer__EVAL_21),
    ._EVAL_22(buffer__EVAL_22),
    ._EVAL_23(buffer__EVAL_23),
    ._EVAL_24(buffer__EVAL_24),
    ._EVAL_25(buffer__EVAL_25),
    ._EVAL_26(buffer__EVAL_26),
    ._EVAL_27(buffer__EVAL_27),
    ._EVAL_28(buffer__EVAL_28),
    ._EVAL_29(buffer__EVAL_29),
    ._EVAL_30(buffer__EVAL_30),
    ._EVAL_31(buffer__EVAL_31),
    ._EVAL_32(buffer__EVAL_32),
    ._EVAL_33(buffer__EVAL_33),
    ._EVAL_34(buffer__EVAL_34),
    ._EVAL_35(buffer__EVAL_35),
    ._EVAL_36(buffer__EVAL_36),
    ._EVAL_37(buffer__EVAL_37),
    ._EVAL_38(buffer__EVAL_38),
    ._EVAL_39(buffer__EVAL_39),
    ._EVAL_40(buffer__EVAL_40),
    ._EVAL_41(buffer__EVAL_41),
    ._EVAL_42(buffer__EVAL_42),
    ._EVAL_43(buffer__EVAL_43),
    ._EVAL_44(buffer__EVAL_44)
  );
  _EVAL_38 ahb2tl (
    ._EVAL(ahb2tl__EVAL),
    ._EVAL_0(ahb2tl__EVAL_0),
    ._EVAL_1(ahb2tl__EVAL_1),
    ._EVAL_2(ahb2tl__EVAL_2),
    ._EVAL_3(ahb2tl__EVAL_3),
    ._EVAL_4(ahb2tl__EVAL_4),
    ._EVAL_5(ahb2tl__EVAL_5),
    ._EVAL_6(ahb2tl__EVAL_6),
    ._EVAL_7(ahb2tl__EVAL_7),
    ._EVAL_8(ahb2tl__EVAL_8),
    ._EVAL_9(ahb2tl__EVAL_9),
    ._EVAL_10(ahb2tl__EVAL_10),
    ._EVAL_11(ahb2tl__EVAL_11),
    ._EVAL_12(ahb2tl__EVAL_12),
    ._EVAL_13(ahb2tl__EVAL_13),
    ._EVAL_14(ahb2tl__EVAL_14),
    ._EVAL_15(ahb2tl__EVAL_15),
    ._EVAL_16(ahb2tl__EVAL_16),
    ._EVAL_17(ahb2tl__EVAL_17),
    ._EVAL_18(ahb2tl__EVAL_18),
    ._EVAL_19(ahb2tl__EVAL_19),
    ._EVAL_20(ahb2tl__EVAL_20),
    ._EVAL_21(ahb2tl__EVAL_21),
    ._EVAL_22(ahb2tl__EVAL_22),
    ._EVAL_23(ahb2tl__EVAL_23),
    ._EVAL_24(ahb2tl__EVAL_24),
    ._EVAL_25(ahb2tl__EVAL_25),
    ._EVAL_26(ahb2tl__EVAL_26),
    ._EVAL_27(ahb2tl__EVAL_27),
    ._EVAL_28(ahb2tl__EVAL_28)
  );
  assign _EVAL_49 = ahb2tl__EVAL_3;
  assign _EVAL_66 = _EVAL_56;
  assign buffer__EVAL_9 = _EVAL_15;
  assign _EVAL_7 = buffer__EVAL_13;
  assign ahb2tl__EVAL_11 = _EVAL_24;
  assign fixer__EVAL_22 = buffer__EVAL_42;
  assign fixer__EVAL_30 = _EVAL_67;
  assign ahb2tl__EVAL_4 = _EVAL_45;
  assign ahb2tl__EVAL_13 = _EVAL_35;
  assign fixer__EVAL_24 = _EVAL_50;
  assign _EVAL_36 = ahb2tl__EVAL_7;
  assign _EVAL_18 = buffer__EVAL_23;
  assign ahb2tl__EVAL_20 = _EVAL_66;
  assign _EVAL_10 = ahb2tl__EVAL_12;
  assign fixer__EVAL_28 = _EVAL_61;
  assign fixer__EVAL_25 = _EVAL_52;
  assign _EVAL_26 = buffer__EVAL_7;
  assign _EVAL_3 = buffer__EVAL_15;
  assign fixer__EVAL_23 = buffer__EVAL_21;
  assign _EVAL_43 = ahb2tl__EVAL_26;
  assign _EVAL_62 = _EVAL_58;
  assign buffer__EVAL_27 = fixer__EVAL_10;
  assign _EVAL_37 = _EVAL_54;
  assign buffer__EVAL_44 = fixer__EVAL_26;
  assign fixer__EVAL_20 = _EVAL_62;
  assign buffer__EVAL_0 = fixer__EVAL;
  assign buffer__EVAL_20 = _EVAL_19;
  assign ahb2tl__EVAL_1 = _EVAL_9;
  assign _EVAL_12 = buffer__EVAL_22;
  assign buffer__EVAL_35 = fixer__EVAL_3;
  assign _EVAL_55 = _EVAL_51;
  assign _EVAL_40 = _EVAL_36;
  assign _EVAL_48 = fixer__EVAL_21;
  assign ahb2tl__EVAL_15 = _EVAL_21;
  assign _EVAL_52 = _EVAL_42;
  assign _EVAL_53 = _EVAL_46;
  assign fixer__EVAL_17 = _EVAL_41;
  assign _EVAL_64 = _EVAL_47;
  assign buffer__EVAL_34 = _EVAL_22;
  assign buffer__EVAL_32 = _EVAL_30;
  assign ahb2tl__EVAL_23 = _EVAL_13;
  assign ahb2tl__EVAL_2 = _EVAL_55;
  assign ahb2tl__EVAL_16 = _EVAL_17;
  assign _EVAL_59 = _EVAL_49;
  assign buffer__EVAL_41 = fixer__EVAL_35;
  assign _EVAL_11 = buffer__EVAL_18;
  assign buffer__EVAL_39 = _EVAL_6;
  assign _EVAL_41 = _EVAL_39;
  assign fixer__EVAL_5 = buffer__EVAL_33;
  assign fixer__EVAL_33 = _EVAL_59;
  assign buffer__EVAL_3 = _EVAL_23;
  assign fixer__EVAL_14 = buffer__EVAL_31;
  assign _EVAL_28 = buffer__EVAL_30;
  assign _EVAL_42 = ahb2tl__EVAL_10;
  assign _EVAL_47 = ahb2tl__EVAL_0;
  assign _EVAL_14 = buffer__EVAL_8;
  assign _EVAL_39 = ahb2tl__EVAL_18;
  assign _EVAL_56 = fixer__EVAL_13;
  assign fixer__EVAL_29 = _EVAL_40;
  assign ahb2tl__EVAL_24 = _EVAL_16;
  assign _EVAL_31 = buffer__EVAL_12;
  assign fixer__EVAL_2 = buffer__EVAL_25;
  assign _EVAL_50 = _EVAL_63;
  assign fixer__EVAL_15 = _EVAL_34;
  assign fixer__EVAL_0 = _EVAL_9;
  assign buffer__EVAL_1 = fixer__EVAL_34;
  assign _EVAL_29 = ahb2tl__EVAL;
  assign fixer__EVAL_11 = buffer__EVAL_2;
  assign _EVAL_58 = ahb2tl__EVAL_27;
  assign buffer__EVAL = _EVAL_9;
  assign fixer__EVAL_19 = buffer__EVAL_36;
  assign _EVAL_44 = ahb2tl__EVAL_6;
  assign ahb2tl__EVAL_28 = _EVAL_2;
  assign buffer__EVAL_29 = fixer__EVAL_8;
  assign ahb2tl__EVAL_14 = _EVAL_34;
  assign _EVAL_46 = ahb2tl__EVAL_9;
  assign _EVAL_54 = fixer__EVAL_18;
  assign ahb2tl__EVAL_25 = _EVAL_8;
  assign buffer__EVAL_5 = _EVAL_34;
  assign _EVAL_60 = _EVAL_48;
  assign _EVAL_32 = ahb2tl__EVAL_5;
  assign fixer__EVAL_36 = buffer__EVAL_10;
  assign buffer__EVAL_38 = fixer__EVAL_27;
  assign _EVAL_63 = ahb2tl__EVAL_21;
  assign buffer__EVAL_16 = fixer__EVAL_7;
  assign _EVAL_67 = _EVAL_44;
  assign buffer__EVAL_6 = _EVAL_27;
  assign fixer__EVAL_31 = _EVAL_53;
  assign _EVAL_61 = _EVAL_57;
  assign buffer__EVAL_11 = fixer__EVAL_32;
  assign _EVAL_51 = fixer__EVAL_4;
  assign ahb2tl__EVAL_17 = _EVAL_37;
  assign _EVAL = buffer__EVAL_19;
  assign _EVAL_57 = ahb2tl__EVAL_19;
  assign _EVAL_38 = fixer__EVAL_16;
  assign _EVAL_4 = buffer__EVAL_26;
  assign fixer__EVAL_6 = buffer__EVAL_43;
  assign fixer__EVAL_1 = _EVAL_64;
  assign _EVAL_20 = buffer__EVAL_4;
  assign buffer__EVAL_28 = fixer__EVAL_37;
  assign fixer__EVAL_12 = buffer__EVAL_17;
  assign ahb2tl__EVAL_22 = _EVAL_25;
  assign ahb2tl__EVAL_8 = _EVAL_60;
  assign _EVAL_33 = buffer__EVAL_24;
  assign _EVAL_65 = _EVAL_43;
  assign buffer__EVAL_37 = _EVAL_1;
  assign _EVAL_0 = buffer__EVAL_14;
  assign buffer__EVAL_40 = _EVAL_5;
  assign _EVAL_45 = _EVAL_38;
  assign fixer__EVAL_9 = _EVAL_65;
endmodule
