//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_41(
  output        _EVAL,
  output [7:0]  _EVAL_0,
  input         _EVAL_1,
  output        _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  output        _EVAL_6,
  input  [3:0]  _EVAL_7,
  output        _EVAL_8,
  output        _EVAL_9,
  output        _EVAL_10,
  input  [31:0] _EVAL_11,
  output        _EVAL_12,
  input  [31:0] _EVAL_13,
  input         _EVAL_14,
  output        _EVAL_15,
  output [3:0]  _EVAL_16,
  input  [2:0]  _EVAL_17,
  output        _EVAL_18,
  output [2:0]  _EVAL_19,
  input  [2:0]  _EVAL_20,
  input  [3:0]  _EVAL_21,
  output        _EVAL_22,
  input         _EVAL_23,
  input  [7:0]  _EVAL_24,
  input         _EVAL_25,
  output        _EVAL_26,
  input  [3:0]  _EVAL_27,
  input  [1:0]  _EVAL_28,
  input         _EVAL_29,
  input         _EVAL_30,
  input         _EVAL_31,
  input  [31:0] _EVAL_32,
  input         _EVAL_33,
  output        _EVAL_34,
  output [31:0] _EVAL_35,
  input         _EVAL_36,
  output [2:0]  _EVAL_37,
  input  [1:0]  _EVAL_38,
  output [31:0] _EVAL_39,
  input  [31:0] _EVAL_40,
  output        _EVAL_41,
  input  [2:0]  _EVAL_42,
  input         _EVAL_43,
  output [3:0]  _EVAL_44,
  input         _EVAL_45,
  output [31:0] _EVAL_46,
  output        _EVAL_47
);
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  coupler_from_port_named_ahb_front_port__EVAL;
  wire  coupler_from_port_named_ahb_front_port__EVAL_0;
  wire  coupler_from_port_named_ahb_front_port__EVAL_1;
  wire  coupler_from_port_named_ahb_front_port__EVAL_2;
  wire  coupler_from_port_named_ahb_front_port__EVAL_3;
  wire  coupler_from_port_named_ahb_front_port__EVAL_4;
  wire [1:0] coupler_from_port_named_ahb_front_port__EVAL_5;
  wire [2:0] coupler_from_port_named_ahb_front_port__EVAL_6;
  wire  coupler_from_port_named_ahb_front_port__EVAL_7;
  wire  coupler_from_port_named_ahb_front_port__EVAL_8;
  wire  coupler_from_port_named_ahb_front_port__EVAL_9;
  wire  coupler_from_port_named_ahb_front_port__EVAL_10;
  wire [3:0] coupler_from_port_named_ahb_front_port__EVAL_11;
  wire [2:0] coupler_from_port_named_ahb_front_port__EVAL_12;
  wire [1:0] coupler_from_port_named_ahb_front_port__EVAL_13;
  wire  coupler_from_port_named_ahb_front_port__EVAL_14;
  wire [3:0] coupler_from_port_named_ahb_front_port__EVAL_15;
  wire  coupler_from_port_named_ahb_front_port__EVAL_16;
  wire  coupler_from_port_named_ahb_front_port__EVAL_17;
  wire  coupler_from_port_named_ahb_front_port__EVAL_18;
  wire [2:0] coupler_from_port_named_ahb_front_port__EVAL_19;
  wire [31:0] coupler_from_port_named_ahb_front_port__EVAL_20;
  wire [31:0] coupler_from_port_named_ahb_front_port__EVAL_21;
  wire  coupler_from_port_named_ahb_front_port__EVAL_22;
  wire [3:0] coupler_from_port_named_ahb_front_port__EVAL_23;
  wire  coupler_from_port_named_ahb_front_port__EVAL_24;
  wire [31:0] coupler_from_port_named_ahb_front_port__EVAL_25;
  wire [3:0] coupler_from_port_named_ahb_front_port__EVAL_26;
  wire [31:0] coupler_from_port_named_ahb_front_port__EVAL_27;
  wire [2:0] coupler_from_port_named_ahb_front_port__EVAL_28;
  wire [31:0] coupler_from_port_named_ahb_front_port__EVAL_29;
  wire  coupler_from_port_named_ahb_front_port__EVAL_30;
  wire  coupler_from_port_named_ahb_front_port__EVAL_31;
  wire [31:0] coupler_from_port_named_ahb_front_port__EVAL_32;
  wire  coupler_from_port_named_ahb_front_port__EVAL_33;
  wire [2:0] coupler_from_port_named_ahb_front_port__EVAL_34;
  wire  coupler_from_port_named_ahb_front_port__EVAL_35;
  wire  _EVAL_51;
  wire [31:0] subsystem_fbus_xbar__EVAL;
  wire  subsystem_fbus_xbar__EVAL_0;
  wire [3:0] subsystem_fbus_xbar__EVAL_1;
  wire [31:0] subsystem_fbus_xbar__EVAL_2;
  wire  subsystem_fbus_xbar__EVAL_3;
  wire [31:0] subsystem_fbus_xbar__EVAL_4;
  wire  subsystem_fbus_xbar__EVAL_5;
  wire  subsystem_fbus_xbar__EVAL_6;
  wire  subsystem_fbus_xbar__EVAL_7;
  wire  subsystem_fbus_xbar__EVAL_8;
  wire [3:0] subsystem_fbus_xbar__EVAL_9;
  wire [2:0] subsystem_fbus_xbar__EVAL_10;
  wire [1:0] subsystem_fbus_xbar__EVAL_11;
  wire [3:0] subsystem_fbus_xbar__EVAL_12;
  wire [2:0] subsystem_fbus_xbar__EVAL_13;
  wire  subsystem_fbus_xbar__EVAL_14;
  wire  subsystem_fbus_xbar__EVAL_15;
  wire [3:0] subsystem_fbus_xbar__EVAL_16;
  wire [2:0] subsystem_fbus_xbar__EVAL_17;
  wire [31:0] subsystem_fbus_xbar__EVAL_18;
  wire  subsystem_fbus_xbar__EVAL_19;
  wire  subsystem_fbus_xbar__EVAL_20;
  wire  subsystem_fbus_xbar__EVAL_21;
  wire [31:0] subsystem_fbus_xbar__EVAL_22;
  wire  subsystem_fbus_xbar__EVAL_23;
  wire  subsystem_fbus_xbar__EVAL_24;
  wire  subsystem_fbus_xbar__EVAL_25;
  wire  subsystem_fbus_xbar__EVAL_26;
  wire  subsystem_fbus_xbar__EVAL_27;
  wire [2:0] subsystem_fbus_xbar__EVAL_28;
  wire [1:0] subsystem_fbus_xbar__EVAL_29;
  wire  subsystem_fbus_xbar__EVAL_30;
  wire  subsystem_fbus_xbar__EVAL_31;
  wire  subsystem_fbus_xbar__EVAL_32;
  wire  subsystem_fbus_xbar__EVAL_33;
  wire [2:0] subsystem_fbus_xbar__EVAL_34;
  wire  subsystem_fbus_xbar__EVAL_35;
  wire  subsystem_fbus_xbar__EVAL_36;
  wire  subsystem_fbus_xbar__EVAL_37;
  wire [3:0] subsystem_fbus_xbar__EVAL_38;
  wire  subsystem_fbus_xbar__EVAL_39;
  wire  subsystem_fbus_xbar__EVAL_40;
  wire  subsystem_fbus_xbar__EVAL_41;
  wire [31:0] subsystem_fbus_xbar__EVAL_42;
  wire [3:0] subsystem_fbus_xbar__EVAL_43;
  wire  subsystem_fbus_xbar__EVAL_44;
  wire [2:0] subsystem_fbus_xbar__EVAL_45;
  wire [3:0] subsystem_fbus_xbar__EVAL_46;
  wire  subsystem_fbus_xbar__EVAL_47;
  wire  subsystem_fbus_xbar__EVAL_48;
  wire [3:0] subsystem_fbus_xbar__EVAL_49;
  wire  subsystem_fbus_xbar__EVAL_50;
  wire [2:0] subsystem_fbus_xbar__EVAL_51;
  wire [31:0] subsystem_fbus_xbar__EVAL_52;
  wire  subsystem_fbus_xbar__EVAL_53;
  wire  subsystem_fbus_xbar__EVAL_54;
  wire  subsystem_fbus_xbar__EVAL_55;
  wire  subsystem_fbus_xbar__EVAL_56;
  wire [31:0] subsystem_fbus_xbar__EVAL_57;
  wire [1:0] subsystem_fbus_xbar__EVAL_58;
  wire  subsystem_fbus_xbar__EVAL_59;
  wire [3:0] subsystem_fbus_xbar__EVAL_60;
  wire  subsystem_fbus_xbar__EVAL_61;
  wire [2:0] subsystem_fbus_xbar__EVAL_62;
  wire [31:0] subsystem_fbus_xbar__EVAL_63;
  wire  buffer__EVAL;
  wire  buffer__EVAL_0;
  wire  buffer__EVAL_1;
  wire  buffer__EVAL_2;
  wire [31:0] buffer__EVAL_3;
  wire  buffer__EVAL_4;
  wire  buffer__EVAL_5;
  wire  buffer__EVAL_6;
  wire [31:0] buffer__EVAL_7;
  wire  buffer__EVAL_8;
  wire  buffer__EVAL_9;
  wire [3:0] buffer__EVAL_10;
  wire  buffer__EVAL_11;
  wire  buffer__EVAL_12;
  wire  buffer__EVAL_13;
  wire [2:0] buffer__EVAL_14;
  wire  buffer__EVAL_15;
  wire  buffer__EVAL_16;
  wire [31:0] buffer__EVAL_17;
  wire [31:0] buffer__EVAL_18;
  wire [3:0] buffer__EVAL_19;
  wire  buffer__EVAL_20;
  wire [2:0] buffer__EVAL_21;
  wire  buffer__EVAL_22;
  wire [2:0] buffer__EVAL_23;
  wire  buffer__EVAL_24;
  wire [3:0] buffer__EVAL_25;
  wire  buffer__EVAL_26;
  wire [2:0] buffer__EVAL_27;
  wire  buffer__EVAL_28;
  wire [31:0] buffer__EVAL_29;
  wire  buffer__EVAL_30;
  wire  buffer__EVAL_31;
  wire [2:0] buffer__EVAL_32;
  wire [2:0] buffer__EVAL_33;
  wire  buffer__EVAL_34;
  wire [31:0] buffer__EVAL_35;
  wire  buffer__EVAL_36;
  wire [1:0] buffer__EVAL_37;
  wire  buffer__EVAL_38;
  wire  buffer__EVAL_39;
  wire [3:0] buffer__EVAL_40;
  wire [1:0] buffer__EVAL_41;
  wire  buffer__EVAL_42;
  wire [3:0] buffer__EVAL_43;
  wire  buffer__EVAL_44;
  wire  buffer__EVAL_45;
  wire  buffer__EVAL_46;
  wire  buffer__EVAL_47;
  wire [3:0] buffer__EVAL_48;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire [7:0] coupler_from_debug_sb__EVAL;
  wire  coupler_from_debug_sb__EVAL_0;
  wire [2:0] coupler_from_debug_sb__EVAL_1;
  wire  coupler_from_debug_sb__EVAL_2;
  wire [3:0] coupler_from_debug_sb__EVAL_3;
  wire [3:0] coupler_from_debug_sb__EVAL_4;
  wire  coupler_from_debug_sb__EVAL_5;
  wire  coupler_from_debug_sb__EVAL_6;
  wire  coupler_from_debug_sb__EVAL_7;
  wire  coupler_from_debug_sb__EVAL_8;
  wire [31:0] coupler_from_debug_sb__EVAL_9;
  wire  coupler_from_debug_sb__EVAL_10;
  wire [3:0] coupler_from_debug_sb__EVAL_11;
  wire [2:0] coupler_from_debug_sb__EVAL_12;
  wire  coupler_from_debug_sb__EVAL_13;
  wire  coupler_from_debug_sb__EVAL_14;
  wire  coupler_from_debug_sb__EVAL_15;
  wire [31:0] coupler_from_debug_sb__EVAL_16;
  wire  coupler_from_debug_sb__EVAL_17;
  wire  coupler_from_debug_sb__EVAL_18;
  wire  coupler_from_debug_sb__EVAL_19;
  wire [7:0] coupler_from_debug_sb__EVAL_20;
  wire  coupler_from_debug_sb__EVAL_21;
  wire [3:0] coupler_from_debug_sb__EVAL_22;
  wire [2:0] coupler_from_debug_sb__EVAL_23;
  wire [31:0] coupler_from_debug_sb__EVAL_24;
  wire [31:0] coupler_from_debug_sb__EVAL_25;
  wire  coupler_from_debug_sb__EVAL_26;
  wire [1:0] coupler_from_debug_sb__EVAL_27;
  _EVAL_40 coupler_from_port_named_ahb_front_port (
    ._EVAL(coupler_from_port_named_ahb_front_port__EVAL),
    ._EVAL_0(coupler_from_port_named_ahb_front_port__EVAL_0),
    ._EVAL_1(coupler_from_port_named_ahb_front_port__EVAL_1),
    ._EVAL_2(coupler_from_port_named_ahb_front_port__EVAL_2),
    ._EVAL_3(coupler_from_port_named_ahb_front_port__EVAL_3),
    ._EVAL_4(coupler_from_port_named_ahb_front_port__EVAL_4),
    ._EVAL_5(coupler_from_port_named_ahb_front_port__EVAL_5),
    ._EVAL_6(coupler_from_port_named_ahb_front_port__EVAL_6),
    ._EVAL_7(coupler_from_port_named_ahb_front_port__EVAL_7),
    ._EVAL_8(coupler_from_port_named_ahb_front_port__EVAL_8),
    ._EVAL_9(coupler_from_port_named_ahb_front_port__EVAL_9),
    ._EVAL_10(coupler_from_port_named_ahb_front_port__EVAL_10),
    ._EVAL_11(coupler_from_port_named_ahb_front_port__EVAL_11),
    ._EVAL_12(coupler_from_port_named_ahb_front_port__EVAL_12),
    ._EVAL_13(coupler_from_port_named_ahb_front_port__EVAL_13),
    ._EVAL_14(coupler_from_port_named_ahb_front_port__EVAL_14),
    ._EVAL_15(coupler_from_port_named_ahb_front_port__EVAL_15),
    ._EVAL_16(coupler_from_port_named_ahb_front_port__EVAL_16),
    ._EVAL_17(coupler_from_port_named_ahb_front_port__EVAL_17),
    ._EVAL_18(coupler_from_port_named_ahb_front_port__EVAL_18),
    ._EVAL_19(coupler_from_port_named_ahb_front_port__EVAL_19),
    ._EVAL_20(coupler_from_port_named_ahb_front_port__EVAL_20),
    ._EVAL_21(coupler_from_port_named_ahb_front_port__EVAL_21),
    ._EVAL_22(coupler_from_port_named_ahb_front_port__EVAL_22),
    ._EVAL_23(coupler_from_port_named_ahb_front_port__EVAL_23),
    ._EVAL_24(coupler_from_port_named_ahb_front_port__EVAL_24),
    ._EVAL_25(coupler_from_port_named_ahb_front_port__EVAL_25),
    ._EVAL_26(coupler_from_port_named_ahb_front_port__EVAL_26),
    ._EVAL_27(coupler_from_port_named_ahb_front_port__EVAL_27),
    ._EVAL_28(coupler_from_port_named_ahb_front_port__EVAL_28),
    ._EVAL_29(coupler_from_port_named_ahb_front_port__EVAL_29),
    ._EVAL_30(coupler_from_port_named_ahb_front_port__EVAL_30),
    ._EVAL_31(coupler_from_port_named_ahb_front_port__EVAL_31),
    ._EVAL_32(coupler_from_port_named_ahb_front_port__EVAL_32),
    ._EVAL_33(coupler_from_port_named_ahb_front_port__EVAL_33),
    ._EVAL_34(coupler_from_port_named_ahb_front_port__EVAL_34),
    ._EVAL_35(coupler_from_port_named_ahb_front_port__EVAL_35)
  );
  _EVAL_25 subsystem_fbus_xbar (
    ._EVAL(subsystem_fbus_xbar__EVAL),
    ._EVAL_0(subsystem_fbus_xbar__EVAL_0),
    ._EVAL_1(subsystem_fbus_xbar__EVAL_1),
    ._EVAL_2(subsystem_fbus_xbar__EVAL_2),
    ._EVAL_3(subsystem_fbus_xbar__EVAL_3),
    ._EVAL_4(subsystem_fbus_xbar__EVAL_4),
    ._EVAL_5(subsystem_fbus_xbar__EVAL_5),
    ._EVAL_6(subsystem_fbus_xbar__EVAL_6),
    ._EVAL_7(subsystem_fbus_xbar__EVAL_7),
    ._EVAL_8(subsystem_fbus_xbar__EVAL_8),
    ._EVAL_9(subsystem_fbus_xbar__EVAL_9),
    ._EVAL_10(subsystem_fbus_xbar__EVAL_10),
    ._EVAL_11(subsystem_fbus_xbar__EVAL_11),
    ._EVAL_12(subsystem_fbus_xbar__EVAL_12),
    ._EVAL_13(subsystem_fbus_xbar__EVAL_13),
    ._EVAL_14(subsystem_fbus_xbar__EVAL_14),
    ._EVAL_15(subsystem_fbus_xbar__EVAL_15),
    ._EVAL_16(subsystem_fbus_xbar__EVAL_16),
    ._EVAL_17(subsystem_fbus_xbar__EVAL_17),
    ._EVAL_18(subsystem_fbus_xbar__EVAL_18),
    ._EVAL_19(subsystem_fbus_xbar__EVAL_19),
    ._EVAL_20(subsystem_fbus_xbar__EVAL_20),
    ._EVAL_21(subsystem_fbus_xbar__EVAL_21),
    ._EVAL_22(subsystem_fbus_xbar__EVAL_22),
    ._EVAL_23(subsystem_fbus_xbar__EVAL_23),
    ._EVAL_24(subsystem_fbus_xbar__EVAL_24),
    ._EVAL_25(subsystem_fbus_xbar__EVAL_25),
    ._EVAL_26(subsystem_fbus_xbar__EVAL_26),
    ._EVAL_27(subsystem_fbus_xbar__EVAL_27),
    ._EVAL_28(subsystem_fbus_xbar__EVAL_28),
    ._EVAL_29(subsystem_fbus_xbar__EVAL_29),
    ._EVAL_30(subsystem_fbus_xbar__EVAL_30),
    ._EVAL_31(subsystem_fbus_xbar__EVAL_31),
    ._EVAL_32(subsystem_fbus_xbar__EVAL_32),
    ._EVAL_33(subsystem_fbus_xbar__EVAL_33),
    ._EVAL_34(subsystem_fbus_xbar__EVAL_34),
    ._EVAL_35(subsystem_fbus_xbar__EVAL_35),
    ._EVAL_36(subsystem_fbus_xbar__EVAL_36),
    ._EVAL_37(subsystem_fbus_xbar__EVAL_37),
    ._EVAL_38(subsystem_fbus_xbar__EVAL_38),
    ._EVAL_39(subsystem_fbus_xbar__EVAL_39),
    ._EVAL_40(subsystem_fbus_xbar__EVAL_40),
    ._EVAL_41(subsystem_fbus_xbar__EVAL_41),
    ._EVAL_42(subsystem_fbus_xbar__EVAL_42),
    ._EVAL_43(subsystem_fbus_xbar__EVAL_43),
    ._EVAL_44(subsystem_fbus_xbar__EVAL_44),
    ._EVAL_45(subsystem_fbus_xbar__EVAL_45),
    ._EVAL_46(subsystem_fbus_xbar__EVAL_46),
    ._EVAL_47(subsystem_fbus_xbar__EVAL_47),
    ._EVAL_48(subsystem_fbus_xbar__EVAL_48),
    ._EVAL_49(subsystem_fbus_xbar__EVAL_49),
    ._EVAL_50(subsystem_fbus_xbar__EVAL_50),
    ._EVAL_51(subsystem_fbus_xbar__EVAL_51),
    ._EVAL_52(subsystem_fbus_xbar__EVAL_52),
    ._EVAL_53(subsystem_fbus_xbar__EVAL_53),
    ._EVAL_54(subsystem_fbus_xbar__EVAL_54),
    ._EVAL_55(subsystem_fbus_xbar__EVAL_55),
    ._EVAL_56(subsystem_fbus_xbar__EVAL_56),
    ._EVAL_57(subsystem_fbus_xbar__EVAL_57),
    ._EVAL_58(subsystem_fbus_xbar__EVAL_58),
    ._EVAL_59(subsystem_fbus_xbar__EVAL_59),
    ._EVAL_60(subsystem_fbus_xbar__EVAL_60),
    ._EVAL_61(subsystem_fbus_xbar__EVAL_61),
    ._EVAL_62(subsystem_fbus_xbar__EVAL_62),
    ._EVAL_63(subsystem_fbus_xbar__EVAL_63)
  );
  _EVAL_29 buffer (
    ._EVAL(buffer__EVAL),
    ._EVAL_0(buffer__EVAL_0),
    ._EVAL_1(buffer__EVAL_1),
    ._EVAL_2(buffer__EVAL_2),
    ._EVAL_3(buffer__EVAL_3),
    ._EVAL_4(buffer__EVAL_4),
    ._EVAL_5(buffer__EVAL_5),
    ._EVAL_6(buffer__EVAL_6),
    ._EVAL_7(buffer__EVAL_7),
    ._EVAL_8(buffer__EVAL_8),
    ._EVAL_9(buffer__EVAL_9),
    ._EVAL_10(buffer__EVAL_10),
    ._EVAL_11(buffer__EVAL_11),
    ._EVAL_12(buffer__EVAL_12),
    ._EVAL_13(buffer__EVAL_13),
    ._EVAL_14(buffer__EVAL_14),
    ._EVAL_15(buffer__EVAL_15),
    ._EVAL_16(buffer__EVAL_16),
    ._EVAL_17(buffer__EVAL_17),
    ._EVAL_18(buffer__EVAL_18),
    ._EVAL_19(buffer__EVAL_19),
    ._EVAL_20(buffer__EVAL_20),
    ._EVAL_21(buffer__EVAL_21),
    ._EVAL_22(buffer__EVAL_22),
    ._EVAL_23(buffer__EVAL_23),
    ._EVAL_24(buffer__EVAL_24),
    ._EVAL_25(buffer__EVAL_25),
    ._EVAL_26(buffer__EVAL_26),
    ._EVAL_27(buffer__EVAL_27),
    ._EVAL_28(buffer__EVAL_28),
    ._EVAL_29(buffer__EVAL_29),
    ._EVAL_30(buffer__EVAL_30),
    ._EVAL_31(buffer__EVAL_31),
    ._EVAL_32(buffer__EVAL_32),
    ._EVAL_33(buffer__EVAL_33),
    ._EVAL_34(buffer__EVAL_34),
    ._EVAL_35(buffer__EVAL_35),
    ._EVAL_36(buffer__EVAL_36),
    ._EVAL_37(buffer__EVAL_37),
    ._EVAL_38(buffer__EVAL_38),
    ._EVAL_39(buffer__EVAL_39),
    ._EVAL_40(buffer__EVAL_40),
    ._EVAL_41(buffer__EVAL_41),
    ._EVAL_42(buffer__EVAL_42),
    ._EVAL_43(buffer__EVAL_43),
    ._EVAL_44(buffer__EVAL_44),
    ._EVAL_45(buffer__EVAL_45),
    ._EVAL_46(buffer__EVAL_46),
    ._EVAL_47(buffer__EVAL_47),
    ._EVAL_48(buffer__EVAL_48)
  );
  _EVAL_33 coupler_from_debug_sb (
    ._EVAL(coupler_from_debug_sb__EVAL),
    ._EVAL_0(coupler_from_debug_sb__EVAL_0),
    ._EVAL_1(coupler_from_debug_sb__EVAL_1),
    ._EVAL_2(coupler_from_debug_sb__EVAL_2),
    ._EVAL_3(coupler_from_debug_sb__EVAL_3),
    ._EVAL_4(coupler_from_debug_sb__EVAL_4),
    ._EVAL_5(coupler_from_debug_sb__EVAL_5),
    ._EVAL_6(coupler_from_debug_sb__EVAL_6),
    ._EVAL_7(coupler_from_debug_sb__EVAL_7),
    ._EVAL_8(coupler_from_debug_sb__EVAL_8),
    ._EVAL_9(coupler_from_debug_sb__EVAL_9),
    ._EVAL_10(coupler_from_debug_sb__EVAL_10),
    ._EVAL_11(coupler_from_debug_sb__EVAL_11),
    ._EVAL_12(coupler_from_debug_sb__EVAL_12),
    ._EVAL_13(coupler_from_debug_sb__EVAL_13),
    ._EVAL_14(coupler_from_debug_sb__EVAL_14),
    ._EVAL_15(coupler_from_debug_sb__EVAL_15),
    ._EVAL_16(coupler_from_debug_sb__EVAL_16),
    ._EVAL_17(coupler_from_debug_sb__EVAL_17),
    ._EVAL_18(coupler_from_debug_sb__EVAL_18),
    ._EVAL_19(coupler_from_debug_sb__EVAL_19),
    ._EVAL_20(coupler_from_debug_sb__EVAL_20),
    ._EVAL_21(coupler_from_debug_sb__EVAL_21),
    ._EVAL_22(coupler_from_debug_sb__EVAL_22),
    ._EVAL_23(coupler_from_debug_sb__EVAL_23),
    ._EVAL_24(coupler_from_debug_sb__EVAL_24),
    ._EVAL_25(coupler_from_debug_sb__EVAL_25),
    ._EVAL_26(coupler_from_debug_sb__EVAL_26),
    ._EVAL_27(coupler_from_debug_sb__EVAL_27)
  );
  assign buffer__EVAL_16 = subsystem_fbus_xbar__EVAL_31;
  assign buffer__EVAL_30 = _EVAL_3;
  assign _EVAL_12 = buffer__EVAL_34;
  assign _EVAL_2 = coupler_from_port_named_ahb_front_port__EVAL_2;
  assign subsystem_fbus_xbar__EVAL_40 = buffer__EVAL_46;
  assign buffer__EVAL_14 = _EVAL_5;
  assign subsystem_fbus_xbar__EVAL = coupler_from_debug_sb__EVAL_16;
  assign buffer__EVAL_15 = _EVAL_52;
  assign subsystem_fbus_xbar__EVAL_22 = coupler_from_debug_sb__EVAL_24;
  assign subsystem_fbus_xbar__EVAL_61 = coupler_from_port_named_ahb_front_port__EVAL_0;
  assign subsystem_fbus_xbar__EVAL_2 = coupler_from_port_named_ahb_front_port__EVAL_32;
  assign coupler_from_debug_sb__EVAL_25 = subsystem_fbus_xbar__EVAL_52;
  assign buffer__EVAL_0 = _EVAL_23;
  assign coupler_from_port_named_ahb_front_port__EVAL_17 = subsystem_fbus_xbar__EVAL_3;
  assign subsystem_fbus_xbar__EVAL_6 = buffer__EVAL_5;
  assign _EVAL_46 = buffer__EVAL_7;
  assign coupler_from_port_named_ahb_front_port__EVAL_13 = _EVAL_38;
  assign subsystem_fbus_xbar__EVAL_18 = buffer__EVAL_3;
  assign _EVAL_0 = coupler_from_debug_sb__EVAL;
  assign coupler_from_debug_sb__EVAL_20 = _EVAL_24;
  assign buffer__EVAL_10 = subsystem_fbus_xbar__EVAL_46;
  assign coupler_from_debug_sb__EVAL_5 = subsystem_fbus_xbar__EVAL_25;
  assign coupler_from_port_named_ahb_front_port__EVAL_10 = _EVAL_45;
  assign subsystem_fbus_xbar__EVAL_32 = coupler_from_debug_sb__EVAL_8;
  assign buffer__EVAL_20 = subsystem_fbus_xbar__EVAL_20;
  assign subsystem_fbus_xbar__EVAL_51 = coupler_from_port_named_ahb_front_port__EVAL_34;
  assign coupler_from_port_named_ahb_front_port__EVAL_1 = _EVAL_52;
  assign subsystem_fbus_xbar__EVAL_49 = coupler_from_port_named_ahb_front_port__EVAL_26;
  assign coupler_from_debug_sb__EVAL_26 = subsystem_fbus_xbar__EVAL_53;
  assign _EVAL_34 = coupler_from_port_named_ahb_front_port__EVAL_30;
  assign coupler_from_port_named_ahb_front_port__EVAL_19 = _EVAL_42;
  assign _EVAL_48 = _EVAL_56;
  assign subsystem_fbus_xbar__EVAL_58 = buffer__EVAL_41;
  assign _EVAL_59 = _EVAL_54;
  assign buffer__EVAL_35 = subsystem_fbus_xbar__EVAL_4;
  assign _EVAL = coupler_from_debug_sb__EVAL_10;
  assign _EVAL_56 = _EVAL_31;
  assign _EVAL_50 = _EVAL_36;
  assign subsystem_fbus_xbar__EVAL_13 = coupler_from_debug_sb__EVAL_1;
  assign coupler_from_debug_sb__EVAL_3 = subsystem_fbus_xbar__EVAL_38;
  assign _EVAL_6 = buffer__EVAL_44;
  assign subsystem_fbus_xbar__EVAL_36 = buffer__EVAL_38;
  assign _EVAL_49 = _EVAL_55;
  assign subsystem_fbus_xbar__EVAL_44 = coupler_from_port_named_ahb_front_port__EVAL_7;
  assign coupler_from_debug_sb__EVAL_27 = subsystem_fbus_xbar__EVAL_29;
  assign coupler_from_port_named_ahb_front_port__EVAL_21 = _EVAL_32;
  assign _EVAL_35 = buffer__EVAL_17;
  assign _EVAL_8 = coupler_from_debug_sb__EVAL_7;
  assign buffer__EVAL_39 = subsystem_fbus_xbar__EVAL_8;
  assign subsystem_fbus_xbar__EVAL_41 = coupler_from_debug_sb__EVAL_0;
  assign coupler_from_port_named_ahb_front_port__EVAL_8 = _EVAL_51;
  assign _EVAL_26 = buffer__EVAL;
  assign subsystem_fbus_xbar__EVAL_1 = coupler_from_debug_sb__EVAL_22;
  assign coupler_from_debug_sb__EVAL_12 = _EVAL_20;
  assign _EVAL_53 = _EVAL_59;
  assign coupler_from_port_named_ahb_front_port__EVAL_16 = subsystem_fbus_xbar__EVAL_26;
  assign coupler_from_port_named_ahb_front_port__EVAL_3 = subsystem_fbus_xbar__EVAL_24;
  assign _EVAL_54 = _EVAL_48;
  assign buffer__EVAL_11 = _EVAL_25;
  assign subsystem_fbus_xbar__EVAL_14 = coupler_from_port_named_ahb_front_port__EVAL;
  assign subsystem_fbus_xbar__EVAL_42 = coupler_from_port_named_ahb_front_port__EVAL_25;
  assign _EVAL_22 = buffer__EVAL_12;
  assign _EVAL_51 = _EVAL_49;
  assign _EVAL_52 = _EVAL_53;
  assign coupler_from_port_named_ahb_front_port__EVAL_11 = _EVAL_21;
  assign subsystem_fbus_xbar__EVAL_5 = buffer__EVAL_8;
  assign coupler_from_debug_sb__EVAL_14 = _EVAL_51;
  assign _EVAL_41 = buffer__EVAL_26;
  assign subsystem_fbus_xbar__EVAL_28 = coupler_from_port_named_ahb_front_port__EVAL_28;
  assign _EVAL_39 = coupler_from_port_named_ahb_front_port__EVAL_27;
  assign _EVAL_47 = buffer__EVAL_42;
  assign coupler_from_port_named_ahb_front_port__EVAL_5 = subsystem_fbus_xbar__EVAL_11;
  assign subsystem_fbus_xbar__EVAL_12 = coupler_from_debug_sb__EVAL_4;
  assign coupler_from_port_named_ahb_front_port__EVAL_24 = _EVAL_43;
  assign subsystem_fbus_xbar__EVAL_16 = coupler_from_port_named_ahb_front_port__EVAL_15;
  assign buffer__EVAL_22 = subsystem_fbus_xbar__EVAL_39;
  assign _EVAL_16 = buffer__EVAL_48;
  assign subsystem_fbus_xbar__EVAL_15 = coupler_from_port_named_ahb_front_port__EVAL_35;
  assign _EVAL_58 = _EVAL_57;
  assign buffer__EVAL_18 = subsystem_fbus_xbar__EVAL_57;
  assign subsystem_fbus_xbar__EVAL_54 = _EVAL_52;
  assign _EVAL_44 = buffer__EVAL_43;
  assign coupler_from_debug_sb__EVAL_6 = subsystem_fbus_xbar__EVAL_59;
  assign subsystem_fbus_xbar__EVAL_56 = coupler_from_port_named_ahb_front_port__EVAL_18;
  assign subsystem_fbus_xbar__EVAL_60 = buffer__EVAL_40;
  assign buffer__EVAL_29 = _EVAL_13;
  assign _EVAL_19 = buffer__EVAL_21;
  assign buffer__EVAL_1 = subsystem_fbus_xbar__EVAL_50;
  assign subsystem_fbus_xbar__EVAL_7 = _EVAL_51;
  assign coupler_from_debug_sb__EVAL_19 = subsystem_fbus_xbar__EVAL_48;
  assign coupler_from_debug_sb__EVAL_15 = _EVAL_30;
  assign _EVAL_10 = buffer__EVAL_28;
  assign coupler_from_debug_sb__EVAL_11 = _EVAL_27;
  assign coupler_from_port_named_ahb_front_port__EVAL_33 = subsystem_fbus_xbar__EVAL_27;
  assign _EVAL_57 = _EVAL_50;
  assign buffer__EVAL_36 = subsystem_fbus_xbar__EVAL_21;
  assign coupler_from_port_named_ahb_front_port__EVAL_6 = _EVAL_17;
  assign coupler_from_port_named_ahb_front_port__EVAL_23 = subsystem_fbus_xbar__EVAL_43;
  assign buffer__EVAL_25 = _EVAL_7;
  assign subsystem_fbus_xbar__EVAL_55 = coupler_from_port_named_ahb_front_port__EVAL_22;
  assign buffer__EVAL_24 = _EVAL_14;
  assign buffer__EVAL_9 = _EVAL_33;
  assign subsystem_fbus_xbar__EVAL_37 = buffer__EVAL_31;
  assign coupler_from_debug_sb__EVAL_9 = _EVAL_11;
  assign buffer__EVAL_37 = _EVAL_28;
  assign subsystem_fbus_xbar__EVAL_23 = coupler_from_port_named_ahb_front_port__EVAL_14;
  assign coupler_from_debug_sb__EVAL_2 = subsystem_fbus_xbar__EVAL_19;
  assign coupler_from_debug_sb__EVAL_17 = _EVAL_52;
  assign _EVAL_15 = coupler_from_debug_sb__EVAL_18;
  assign coupler_from_port_named_ahb_front_port__EVAL_31 = _EVAL_1;
  assign _EVAL_18 = buffer__EVAL_47;
  assign coupler_from_port_named_ahb_front_port__EVAL_4 = subsystem_fbus_xbar__EVAL_35;
  assign coupler_from_debug_sb__EVAL_23 = subsystem_fbus_xbar__EVAL_34;
  assign buffer__EVAL_4 = subsystem_fbus_xbar__EVAL_47;
  assign buffer__EVAL_13 = _EVAL_29;
  assign _EVAL_9 = coupler_from_debug_sb__EVAL_13;
  assign _EVAL_55 = _EVAL_58;
  assign buffer__EVAL_19 = subsystem_fbus_xbar__EVAL_9;
  assign buffer__EVAL_33 = subsystem_fbus_xbar__EVAL_45;
  assign coupler_from_port_named_ahb_front_port__EVAL_12 = subsystem_fbus_xbar__EVAL_10;
  assign _EVAL_37 = buffer__EVAL_32;
  assign buffer__EVAL_45 = _EVAL_51;
  assign subsystem_fbus_xbar__EVAL_0 = coupler_from_port_named_ahb_front_port__EVAL_9;
  assign coupler_from_port_named_ahb_front_port__EVAL_29 = _EVAL_40;
  assign coupler_from_port_named_ahb_front_port__EVAL_20 = subsystem_fbus_xbar__EVAL_63;
  assign subsystem_fbus_xbar__EVAL_62 = buffer__EVAL_23;
  assign buffer__EVAL_27 = subsystem_fbus_xbar__EVAL_17;
  assign buffer__EVAL_2 = subsystem_fbus_xbar__EVAL_33;
  assign coupler_from_debug_sb__EVAL_21 = _EVAL_4;
  assign subsystem_fbus_xbar__EVAL_30 = buffer__EVAL_6;
endmodule
