//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_105(
  output        _EVAL,
  input  [31:0] _EVAL_0,
  input  [29:0] _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input  [29:0] _EVAL_5,
  input         _EVAL_6,
  input  [1:0]  _EVAL_7,
  input         _EVAL_8,
  output        _EVAL_9,
  input  [1:0]  _EVAL_10,
  input  [1:0]  _EVAL_11,
  input  [1:0]  _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input  [1:0]  _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18,
  input         _EVAL_19,
  input  [29:0] _EVAL_20,
  input         _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23,
  input  [31:0] _EVAL_24,
  input         _EVAL_25,
  input         _EVAL_26,
  input  [31:0] _EVAL_27,
  input  [31:0] _EVAL_28,
  input  [31:0] _EVAL_29,
  input         _EVAL_30,
  input  [1:0]  _EVAL_31,
  input  [1:0]  _EVAL_32,
  input  [29:0] _EVAL_33,
  input  [31:0] _EVAL_34,
  input         _EVAL_35,
  input         _EVAL_36,
  input         _EVAL_37,
  input  [31:0] _EVAL_38,
  input  [31:0] _EVAL_39,
  input  [1:0]  _EVAL_40,
  input  [29:0] _EVAL_41,
  input  [29:0] _EVAL_42,
  input         _EVAL_43,
  input         _EVAL_44,
  input  [29:0] _EVAL_45,
  input  [31:0] _EVAL_46,
  input  [1:0]  _EVAL_47,
  input         _EVAL_48,
  input         _EVAL_49,
  input         _EVAL_50,
  input         _EVAL_51,
  input         _EVAL_52,
  input  [29:0] _EVAL_53,
  output        _EVAL_54,
  input         _EVAL_55,
  input         _EVAL_56,
  input         _EVAL_57,
  input         _EVAL_58,
  input         _EVAL_59,
  input         _EVAL_60,
  input         _EVAL_61
);
  wire  _EVAL_63;
  wire [31:0] _EVAL_64;
  wire  _EVAL_67;
  wire [31:0] _EVAL_68;
  wire  _EVAL_70;
  wire  _EVAL_72;
  wire  _EVAL_74;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire [31:0] _EVAL_80;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire [31:0] _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_94;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_103;
  wire [31:0] _EVAL_105;
  wire  _EVAL_111;
  wire  _EVAL_113;
  wire [31:0] _EVAL_115;
  wire  _EVAL_116;
  wire [31:0] _EVAL_117;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_122;
  wire  _EVAL_125;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire [31:0] _EVAL_130;
  wire [31:0] _EVAL_132;
  wire  _EVAL_134;
  wire [31:0] _EVAL_135;
  wire [31:0] _EVAL_137;
  wire [31:0] _EVAL_139;
  wire [31:0] _EVAL_140;
  wire  _EVAL_143;
  wire [31:0] _EVAL_144;
  wire  _EVAL_145;
  wire [31:0] _EVAL_146;
  wire  _EVAL_147;
  wire [31:0] _EVAL_148;
  wire [31:0] _EVAL_150;
  wire [31:0] _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire [31:0] _EVAL_162;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_177;
  wire [31:0] _EVAL_179;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire [31:0] _EVAL_183;
  wire  _EVAL_185;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire [31:0] _EVAL_196;
  wire  _EVAL_198;
  wire [31:0] _EVAL_202;
  wire [31:0] _EVAL_203;
  wire  _EVAL_204;
  wire [31:0] _EVAL_205;
  wire [31:0] _EVAL_207;
  wire [31:0] _EVAL_208;
  wire [31:0] _EVAL_209;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire [31:0] _EVAL_218;
  wire  _EVAL_223;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire [31:0] _EVAL_228;
  wire  _EVAL_231;
  wire [31:0] _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire [31:0] _EVAL_236;
  wire [31:0] _EVAL_239;
  wire [31:0] _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_244;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_251;
  wire [31:0] _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_259;
  wire  _EVAL_261;
  wire  _EVAL_263;
  wire [31:0] _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire [31:0] _EVAL_267;
  wire [31:0] _EVAL_268;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_277;
  wire [31:0] _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_283;
  wire  _EVAL_285;
  wire [31:0] _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire [31:0] _EVAL_291;
  wire [31:0] _EVAL_292;
  wire  _EVAL_294;
  wire [31:0] _EVAL_297;
  wire  _EVAL_302;
  wire [31:0] _EVAL_303;
  wire [31:0] _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_308;
  wire [31:0] _EVAL_314;
  wire  _EVAL_317;
  wire  _EVAL_320;
  wire  _EVAL_321;
  wire [31:0] _EVAL_322;
  wire [31:0] _EVAL_323;
  wire  _EVAL_324;
  wire [31:0] _EVAL_325;
  wire  _EVAL_327;
  wire  _EVAL_328;
  wire  _EVAL_330;
  wire [31:0] _EVAL_331;
  wire  _EVAL_332;
  wire  _EVAL_334;
  wire  _EVAL_336;
  wire  _EVAL_344;
  wire  _EVAL_345;
  wire  _EVAL_348;
  wire [31:0] _EVAL_354;
  wire  _EVAL_357;
  wire  _EVAL_361;
  wire  _EVAL_364;
  wire [31:0] _EVAL_366;
  wire [31:0] _EVAL_367;
  wire  _EVAL_370;
  wire [31:0] _EVAL_374;
  wire  _EVAL_376;
  wire [31:0] _EVAL_377;
  wire  _EVAL_378;
  wire  _EVAL_379;
  wire [31:0] _EVAL_381;
  wire  _EVAL_386;
  wire  _EVAL_389;
  wire  _EVAL_392;
  wire  _EVAL_396;
  wire  _EVAL_397;
  wire  _EVAL_400;
  wire  _EVAL_401;
  assign _EVAL_103 = _EVAL_32[0];
  assign _EVAL_364 = _EVAL_308 ? _EVAL_246 : _EVAL_190;
  assign _EVAL_361 = _EVAL_308 ? _EVAL_100 : _EVAL_227;
  assign _EVAL_325 = ~_EVAL_130;
  assign _EVAL_345 = _EVAL_94 & _EVAL_86;
  assign _EVAL_161 = _EVAL_321 & _EVAL_70;
  assign _EVAL_113 = _EVAL_327 & _EVAL_116;
  assign _EVAL_287 = _EVAL_16[1];
  assign _EVAL_265 = _EVAL_202 == 32'h0;
  assign _EVAL_357 = _EVAL_103 & _EVAL_397;
  assign _EVAL_152 = _EVAL_10[0];
  assign _EVAL_366 = _EVAL_322 | 32'h3;
  assign _EVAL_244 = ~_EVAL_43;
  assign _EVAL_209 = ~_EVAL_305;
  assign _EVAL_193 = _EVAL_83 & _EVAL_122;
  assign _EVAL_332 = _EVAL_327 & _EVAL_324;
  assign _EVAL_272 = _EVAL_31[0];
  assign _EVAL_277 = _EVAL_251 & _EVAL_345;
  assign _EVAL_305 = {_EVAL_53, 2'h0};
  assign _EVAL_181 = _EVAL_223 ? _EVAL_401 : _EVAL_334;
  assign _EVAL_344 = _EVAL_80 == 32'h0;
  assign _EVAL_179 = _EVAL_38 ^ _EVAL_236;
  assign _EVAL_247 = _EVAL_242 & _EVAL_166;
  assign _EVAL_155 = ~_EVAL_61;
  assign _EVAL_146 = _EVAL_209 | 32'h3;
  assign _EVAL_9 = _EVAL_119 ? _EVAL_283 : _EVAL_235;
  assign _EVAL_207 = _EVAL_140 | 32'h3;
  assign _EVAL_367 = _EVAL_38 ^ _EVAL_68;
  assign _EVAL_83 = ~_EVAL_70;
  assign _EVAL_292 = ~_EVAL_233;
  assign _EVAL_236 = ~_EVAL_366;
  assign _EVAL_115 = ~_EVAL_377;
  assign _EVAL_137 = ~_EVAL_150;
  assign _EVAL_290 = _EVAL_151 == 32'h0;
  assign _EVAL_314 = _EVAL_264 & _EVAL_381;
  assign _EVAL_203 = ~_EVAL_253;
  assign _EVAL_242 = _EVAL_40[0];
  assign _EVAL_162 = {_EVAL_20, 2'h0};
  assign _EVAL_100 = _EVAL_49 | _EVAL_332;
  assign _EVAL_271 = _EVAL_23 | _EVAL_173;
  assign _EVAL_72 = _EVAL_57 | _EVAL_113;
  assign _EVAL_168 = ~_EVAL_88;
  assign _EVAL_323 = {_EVAL_41, 2'h0};
  assign _EVAL_150 = _EVAL_292 | 32'h3;
  assign _EVAL_119 = _EVAL_189 ? _EVAL_344 : _EVAL_255;
  assign _EVAL_261 = _EVAL_55 | _EVAL_84;
  assign _EVAL_320 = _EVAL_127 & _EVAL_234;
  assign _EVAL_370 = _EVAL_11[0];
  assign _EVAL_233 = {_EVAL_5, 2'h0};
  assign _EVAL_143 = _EVAL_32[1];
  assign _EVAL_68 = ~_EVAL_218;
  assign _EVAL_160 = _EVAL_308 ? _EVAL_134 : _EVAL_182;
  assign _EVAL_85 = ~_EVAL_24;
  assign _EVAL_289 = _EVAL_60 | _EVAL_173;
  assign _EVAL_169 = _EVAL_48 | _EVAL_113;
  assign _EVAL_223 = _EVAL_11[1];
  assign _EVAL_74 = _EVAL_58 | _EVAL_248;
  assign _EVAL_78 = _EVAL_22 | _EVAL_328;
  assign _EVAL_187 = _EVAL_44 | _EVAL_378;
  assign _EVAL_322 = ~_EVAL_323;
  assign _EVAL_183 = _EVAL_38 ^ _EVAL_135;
  assign _EVAL_185 = _EVAL_132 == 32'h0;
  assign _EVAL_63 = _EVAL_36 | _EVAL_173;
  assign _EVAL_396 = _EVAL_143 ? _EVAL_265 : _EVAL_357;
  assign _EVAL_381 = ~_EVAL_29;
  assign _EVAL_215 = _EVAL_254 ? _EVAL_289 : _EVAL_156;
  assign _EVAL_234 = _EVAL_38 < _EVAL_139;
  assign _EVAL_84 = _EVAL_327 & _EVAL_256;
  assign _EVAL_172 = _EVAL_21 | _EVAL_113;
  assign _EVAL_334 = _EVAL_370 & _EVAL_161;
  assign _EVAL_145 = _EVAL_3 | _EVAL_378;
  assign _EVAL_392 = _EVAL_17 | _EVAL_84;
  assign _EVAL_266 = _EVAL_31[1];
  assign _EVAL_191 = _EVAL_254 ? _EVAL_63 : _EVAL_120;
  assign _EVAL_190 = _EVAL_204 ? _EVAL_169 : _EVAL_191;
  assign _EVAL_182 = _EVAL_204 ? _EVAL_72 : _EVAL_215;
  assign _EVAL_294 = ~_EVAL_35;
  assign _EVAL_89 = _EVAL_18 | _EVAL_159;
  assign _EVAL_99 = _EVAL_10[1];
  assign _EVAL_267 = ~_EVAL_162;
  assign _EVAL_196 = ~_EVAL_39;
  assign _EVAL_286 = {_EVAL_1, 2'h0};
  assign _EVAL_120 = _EVAL_285 ? _EVAL_145 : _EVAL_336;
  assign _EVAL_331 = ~_EVAL_34;
  assign _EVAL_202 = _EVAL_367 & _EVAL_331;
  assign _EVAL_148 = ~_EVAL_144;
  assign _EVAL_144 = {_EVAL_42, 2'h0};
  assign _EVAL_274 = _EVAL_297 == 32'h0;
  assign _EVAL_140 = ~_EVAL_286;
  assign _EVAL_400 = ~_EVAL_51;
  assign _EVAL_227 = _EVAL_204 ? _EVAL_172 : _EVAL_67;
  assign _EVAL_198 = ~_EVAL_167;
  assign _EVAL_275 = _EVAL_26 | _EVAL_159;
  assign _EVAL_132 = _EVAL_183 & _EVAL_196;
  assign _EVAL_139 = ~_EVAL_291;
  assign _EVAL_122 = _EVAL_38 < _EVAL_115;
  assign _EVAL_90 = _EVAL_152 & _EVAL_111;
  assign _EVAL_328 = _EVAL_327 & _EVAL_400;
  assign _EVAL_240 = {_EVAL_33, 2'h0};
  assign _EVAL_389 = _EVAL_125 ? _EVAL_171 : _EVAL_327;
  assign _EVAL_156 = _EVAL_285 ? _EVAL_187 : _EVAL_241;
  assign _EVAL_324 = ~_EVAL_6;
  assign _EVAL_64 = ~_EVAL_0;
  assign _EVAL_354 = ~_EVAL_146;
  assign _EVAL_151 = _EVAL_117 & _EVAL_239;
  assign _EVAL_253 = {_EVAL_45, 2'h0};
  assign _EVAL_116 = ~_EVAL_19;
  assign _EVAL_94 = ~_EVAL_288;
  assign _EVAL_302 = ~_EVAL_234;
  assign _EVAL_256 = ~_EVAL_13;
  assign _EVAL_268 = ~_EVAL_28;
  assign _EVAL_321 = ~_EVAL_86;
  assign _EVAL_86 = _EVAL_38 < _EVAL_236;
  assign _EVAL_248 = _EVAL_327 & _EVAL_294;
  assign _EVAL_135 = ~_EVAL_207;
  assign _EVAL_192 = _EVAL_8 | _EVAL_378;
  assign _EVAL_303 = _EVAL_38 ^ _EVAL_354;
  assign _EVAL_79 = _EVAL_285 ? _EVAL_192 : _EVAL_379;
  assign _EVAL_214 = ~_EVAL_2;
  assign _EVAL_188 = _EVAL_15 | _EVAL_248;
  assign _EVAL_134 = _EVAL_4 | _EVAL_332;
  assign _EVAL_288 = _EVAL_38 < _EVAL_137;
  assign _EVAL_241 = _EVAL_181 ? _EVAL_392 : _EVAL_330;
  assign _EVAL_255 = _EVAL_157 & _EVAL_167;
  assign _EVAL = _EVAL_119 ? _EVAL_78 : _EVAL_231;
  assign _EVAL_235 = _EVAL_396 ? _EVAL_275 : _EVAL_364;
  assign _EVAL_226 = _EVAL_16[0];
  assign _EVAL_204 = _EVAL_99 ? _EVAL_185 : _EVAL_90;
  assign _EVAL_205 = ~_EVAL_240;
  assign _EVAL_283 = _EVAL_25 | _EVAL_328;
  assign _EVAL_264 = _EVAL_38 ^ _EVAL_139;
  assign _EVAL_159 = _EVAL_327 & _EVAL_155;
  assign _EVAL_377 = _EVAL_148 | 32'h3;
  assign _EVAL_386 = _EVAL_396 ? _EVAL_348 : _EVAL_160;
  assign _EVAL_228 = ~_EVAL_27;
  assign _EVAL_67 = _EVAL_254 ? _EVAL_271 : _EVAL_79;
  assign _EVAL_166 = _EVAL_168 & _EVAL_288;
  assign _EVAL_111 = _EVAL_302 & _EVAL_88;
  assign _EVAL_263 = _EVAL_56 | _EVAL_84;
  assign _EVAL_231 = _EVAL_396 ? _EVAL_89 : _EVAL_361;
  assign _EVAL_279 = _EVAL_179 & _EVAL_228;
  assign _EVAL_308 = _EVAL_287 ? _EVAL_376 : _EVAL_306;
  assign _EVAL_285 = _EVAL_177 ? _EVAL_158 : _EVAL_277;
  assign _EVAL_125 = _EVAL_266 ? _EVAL_274 : _EVAL_280;
  assign _EVAL_70 = _EVAL_38 < _EVAL_354;
  assign _EVAL_297 = _EVAL_374 & _EVAL_64;
  assign _EVAL_117 = _EVAL_38 ^ _EVAL_137;
  assign _EVAL_306 = _EVAL_226 & _EVAL_320;
  assign _EVAL_401 = _EVAL_105 == 32'h0;
  assign _EVAL_376 = _EVAL_314 == 32'h0;
  assign _EVAL_127 = ~_EVAL_317;
  assign _EVAL_54 = _EVAL_119 ? _EVAL_147 : _EVAL_386;
  assign _EVAL_379 = _EVAL_181 ? _EVAL_261 : _EVAL_259;
  assign _EVAL_171 = _EVAL_52 | _EVAL_248;
  assign _EVAL_374 = _EVAL_38 ^ _EVAL_115;
  assign _EVAL_280 = _EVAL_272 & _EVAL_193;
  assign _EVAL_348 = _EVAL_50 | _EVAL_159;
  assign _EVAL_246 = _EVAL_14 | _EVAL_332;
  assign _EVAL_189 = _EVAL_12[1];
  assign _EVAL_336 = _EVAL_181 ? _EVAL_263 : _EVAL_389;
  assign _EVAL_317 = _EVAL_38 < _EVAL_68;
  assign _EVAL_128 = _EVAL_40[1];
  assign _EVAL_254 = _EVAL_128 ? _EVAL_290 : _EVAL_247;
  assign _EVAL_173 = _EVAL_327 & _EVAL_244;
  assign _EVAL_147 = _EVAL_59 | _EVAL_328;
  assign _EVAL_259 = _EVAL_125 ? _EVAL_74 : _EVAL_327;
  assign _EVAL_130 = _EVAL_203 | 32'h3;
  assign _EVAL_158 = _EVAL_279 == 32'h0;
  assign _EVAL_80 = _EVAL_208 & _EVAL_268;
  assign _EVAL_88 = _EVAL_38 < _EVAL_135;
  assign _EVAL_105 = _EVAL_303 & _EVAL_85;
  assign _EVAL_167 = _EVAL_38 < _EVAL_325;
  assign _EVAL_251 = _EVAL_7[0];
  assign _EVAL_378 = _EVAL_327 & _EVAL_214;
  assign _EVAL_397 = _EVAL_198 & _EVAL_317;
  assign _EVAL_327 = _EVAL_47 > 2'h1;
  assign _EVAL_291 = _EVAL_267 | 32'h3;
  assign _EVAL_218 = _EVAL_205 | 32'h3;
  assign _EVAL_330 = _EVAL_125 ? _EVAL_188 : _EVAL_327;
  assign _EVAL_157 = _EVAL_12[0];
  assign _EVAL_208 = _EVAL_38 ^ _EVAL_325;
  assign _EVAL_239 = ~_EVAL_46;
  assign _EVAL_177 = _EVAL_7[1];
endmodule
