//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_194_assert(
  input  [9:0]  _EVAL,
  input  [14:0] _EVAL_0,
  input         _EVAL_1,
  input  [2:0]  _EVAL_2,
  input  [3:0]  _EVAL_3,
  input  [1:0]  _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input  [1:0]  _EVAL_8,
  input         _EVAL_9,
  input  [2:0]  _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input  [9:0]  _EVAL_13
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [575:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_14;
  wire  _EVAL_15;
  wire  _EVAL_16;
  reg [1:0] _EVAL_17;
  reg [9:0] _EVAL_18;
  wire [1:0] _EVAL_19;
  wire  _EVAL_20;
  wire [1:0] _EVAL_21;
  wire [1:0] _EVAL_22;
  wire [1:0] _EVAL_23;
  wire [14:0] _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  reg [14:0] _EVAL_28;
  wire [3:0] _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_32;
  wire  _EVAL_33;
  reg [31:0] _EVAL_34;
  wire [575:0] _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  reg [2:0] _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire [1023:0] _EVAL_41;
  wire [1:0] _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire [1023:0] _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire [4:0] _EVAL_55;
  wire  _EVAL_56;
  reg  _EVAL_57;
  wire  _EVAL_58;
  wire [15:0] _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  reg [1:0] _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  reg  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  reg [575:0] _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  reg [2:0] _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire [1:0] _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  reg [2:0] _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire [15:0] _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  reg  _EVAL_95;
  wire [14:0] _EVAL_96;
  wire [3:0] _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  reg  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire [1023:0] _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire [32:0] _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire [575:0] _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire [1023:0] _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire [3:0] _EVAL_136;
  wire  _EVAL_137;
  wire [14:0] _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire [575:0] _EVAL_143;
  wire [1:0] _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  reg [9:0] _EVAL_149;
  wire [31:0] _EVAL_150;
  wire  _EVAL_151;
  wire [575:0] _EVAL_152;
  wire [3:0] _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire [15:0] _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire [1:0] _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire [575:0] _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire [575:0] _EVAL_182;
  wire  _EVAL_183;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire [575:0] _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_112 = _EVAL_49 & _EVAL_204;
  assign _EVAL_83 = 2'h1 << _EVAL_192;
  assign _EVAL_14 = _EVAL_9 & _EVAL_66;
  assign _EVAL_155 = _EVAL_5 == 3'h7;
  assign _EVAL_52 = _EVAL_47 ? _EVAL_41 : 1024'h0;
  assign _EVAL_144 = _EVAL_104 - 1'h1;
  assign _EVAL_168 = _EVAL_6 & _EVAL_50;
  assign _EVAL_157 = _EVAL_22[1];
  assign _EVAL_101 = _EVAL_34 < plusarg_reader_out;
  assign _EVAL_56 = _EVAL_9 & _EVAL_125;
  assign _EVAL_51 = _EVAL_127 | _EVAL_48;
  assign _EVAL_42 = _EVAL_55[1:0];
  assign _EVAL_77 = ~_EVAL_54;
  assign _EVAL_143 = _EVAL_188 | _EVAL_71;
  assign _EVAL_102 = _EVAL_24 == 15'h0;
  assign _EVAL_73 = _EVAL_6 & _EVAL_139;
  assign _EVAL_160 = ~_EVAL_102;
  assign _EVAL_63 = _EVAL_176 & _EVAL_142;
  assign _EVAL_195 = _EVAL_6 & _EVAL_32;
  assign _EVAL_36 = ~_EVAL_81;
  assign _EVAL_154 = |_EVAL_71;
  assign _EVAL_185 = _EVAL_2 <= 3'h2;
  assign _EVAL_190 = _EVAL_188 != _EVAL_35;
  assign _EVAL_163 = _EVAL_0[1];
  assign _EVAL_182 = _EVAL_71 | _EVAL_188;
  assign _EVAL_180 = _EVAL_81 & _EVAL_63;
  assign _EVAL_199 = _EVAL_5 == 3'h0;
  assign _EVAL_15 = ~_EVAL_170;
  assign _EVAL_198 = ~_EVAL_163;
  assign _EVAL_107 = ~_EVAL_126;
  assign _EVAL_53 = _EVAL_137 & _EVAL_135;
  assign _EVAL_178 = _EVAL_71 >> _EVAL_13;
  assign _EVAL_125 = _EVAL_10 == 3'h1;
  assign _EVAL_197 = ~_EVAL_167;
  assign _EVAL_177 = _EVAL_5 == 3'h6;
  assign _EVAL_90 = ~_EVAL_66;
  assign _EVAL_84 = _EVAL_9 & _EVAL_158;
  assign _EVAL_156 = ~_EVAL_33;
  assign _EVAL_202 = _EVAL_6 & _EVAL_116;
  assign _EVAL_184 = _EVAL_10 == 3'h4;
  assign _EVAL_67 = ~_EVAL_118;
  assign _EVAL_35 = _EVAL_52[575:0];
  assign _EVAL_108 = _EVAL_6 & _EVAL_109;
  assign _EVAL_147 = ~_EVAL_185;
  assign _EVAL_193 = ~_EVAL_154;
  assign _EVAL_131 = _EVAL_198 & _EVAL_100;
  assign _EVAL_58 = _EVAL_2 == _EVAL_87;
  assign _EVAL_123 = ~_EVAL_159;
  assign _EVAL_54 = _EVAL_29 == 4'h0;
  assign _EVAL_133 = ~_EVAL_122;
  assign _EVAL_61 = ~_EVAL_180;
  assign _EVAL_37 = ~_EVAL_204;
  assign _EVAL_81 = _EVAL_13 <= 10'h23f;
  assign _EVAL_192 = _EVAL_8[0];
  assign _EVAL_129 = _EVAL_3 == _EVAL_136;
  assign _EVAL_92 = _EVAL_44 | _EVAL_43;
  assign _EVAL_74 = _EVAL_9 & _EVAL_62;
  assign _EVAL_109 = _EVAL_5 == 3'h5;
  assign _EVAL_175 = ~_EVAL_42;
  assign _EVAL_103 = ~_EVAL_57;
  assign _EVAL_170 = _EVAL_4 == _EVAL_65;
  assign _EVAL_164 = _EVAL_10 == 3'h0;
  assign _EVAL_116 = _EVAL_5 == 3'h3;
  assign _EVAL_117 = ~_EVAL_80;
  assign _EVAL_165 = ~_EVAL_20;
  assign _EVAL_40 = ~_EVAL_191;
  assign _EVAL_111 = _EVAL_9 & _EVAL_184;
  assign _EVAL_76 = ~_EVAL_30;
  assign _EVAL_69 = _EVAL_198 & _EVAL_75;
  assign _EVAL_128 = _EVAL_143 >> _EVAL;
  assign _EVAL_162 = _EVAL_127 | _EVAL_25;
  assign _EVAL_55 = 5'h3 << _EVAL_8;
  assign _EVAL_188 = _EVAL_132[575:0];
  assign _EVAL_91 = $signed(_EVAL_171) & -16'sh1000;
  assign _EVAL_159 = _EVAL_2 <= 3'h3;
  assign _EVAL_89 = ~_EVAL_194;
  assign _EVAL_189 = _EVAL_153 == 4'h0;
  assign _EVAL_49 = _EVAL_1 & _EVAL_6;
  assign _EVAL_66 = _EVAL_10 == 3'h6;
  assign _EVAL_142 = $signed(_EVAL_59) == 16'sh0;
  assign _EVAL_203 = _EVAL_21[0];
  assign _EVAL_80 = _EVAL_190 | _EVAL_186;
  assign _EVAL_110 = _EVAL_23[0];
  assign _EVAL_127 = _EVAL_183 | _EVAL_169;
  assign _EVAL_32 = _EVAL_5 == 3'h1;
  assign _EVAL_139 = _EVAL_5 == 3'h2;
  assign _EVAL_113 = _EVAL_178[0];
  assign _EVAL_146 = _EVAL_9 & _EVAL_173;
  assign _EVAL_82 = _EVAL_12 & _EVAL_9;
  assign _EVAL_50 = _EVAL_5 == 3'h4;
  assign _EVAL_145 = ~_EVAL_46;
  assign _EVAL_126 = _EVAL_201 | _EVAL_101;
  assign _EVAL_179 = ~_EVAL_119;
  assign _EVAL_141 = ~_EVAL_104;
  assign _EVAL_173 = _EVAL_10 == 3'h2;
  assign _EVAL_205 = ~_EVAL_95;
  assign _EVAL_59 = _EVAL_91;
  assign _EVAL_140 = _EVAL_9 & _EVAL_164;
  assign _EVAL_176 = _EVAL_8 <= 2'h2;
  assign _EVAL_21 = _EVAL_95 - 1'h1;
  assign _EVAL_166 = ~_EVAL_129;
  assign _EVAL_44 = _EVAL_183 | _EVAL_72;
  assign _EVAL_45 = _EVAL_6 & _EVAL_155;
  assign _EVAL_124 = |_EVAL_188;
  assign _EVAL_137 = _EVAL_22[0];
  assign _EVAL_204 = ~_EVAL_68;
  assign _EVAL_153 = ~_EVAL_3;
  assign _EVAL_132 = _EVAL_93 ? _EVAL_115 : 1024'h0;
  assign _EVAL_99 = ~_EVAL_187;
  assign _EVAL_201 = _EVAL_193 | _EVAL_200;
  assign _EVAL_136 = {_EVAL_92,_EVAL_181,_EVAL_51,_EVAL_162};
  assign _EVAL_24 = _EVAL_0 & _EVAL_96;
  assign _EVAL_183 = _EVAL_8 >= 2'h2;
  assign _EVAL_120 = _EVAL_34 + 32'h1;
  assign _EVAL_169 = _EVAL_157 & _EVAL_198;
  assign _EVAL_151 = ~_EVAL_130;
  assign _EVAL_20 = _EVAL <= 10'h23f;
  assign _EVAL_119 = ~_EVAL_113;
  assign _EVAL_85 = ~_EVAL_58;
  assign _EVAL_171 = {1'b0,$signed(_EVAL_138)};
  assign _EVAL_100 = _EVAL_0[0];
  assign _EVAL_194 = _EVAL_0 == _EVAL_28;
  assign _EVAL_167 = _EVAL_2 <= 3'h1;
  assign _EVAL_39 = _EVAL_6 & _EVAL_177;
  assign _EVAL_94 = ~_EVAL_189;
  assign _EVAL_64 = _EVAL_82 & _EVAL_141;
  assign _EVAL_46 = _EVAL_5 == _EVAL_38;
  assign _EVAL_75 = ~_EVAL_100;
  assign _EVAL_19 = _EVAL_57 - 1'h1;
  assign _EVAL_98 = ~_EVAL_183;
  assign _EVAL_118 = _EVAL_10 <= 3'h6;
  assign _EVAL_134 = ~_EVAL_148;
  assign _EVAL_122 = _EVAL_13 == _EVAL_18;
  assign _EVAL_135 = _EVAL_163 & _EVAL_75;
  assign _EVAL_174 = ~_EVAL_105;
  assign _EVAL_70 = ~_EVAL_206;
  assign _EVAL_206 = _EVAL_10 == _EVAL_79;
  assign _EVAL_93 = _EVAL_49 & _EVAL_103;
  assign _EVAL_105 = _EVAL_2 == 3'h0;
  assign _EVAL_30 = _EVAL_128[0];
  assign _EVAL_130 = ~_EVAL_7;
  assign _EVAL_186 = ~_EVAL_124;
  assign _EVAL_47 = _EVAL_26 & _EVAL_90;
  assign _EVAL_78 = ~_EVAL_86;
  assign _EVAL_26 = _EVAL_82 & _EVAL_205;
  assign _EVAL_200 = plusarg_reader_out == 32'h0;
  assign _EVAL_23 = _EVAL_68 - 1'h1;
  assign _EVAL_72 = _EVAL_157 & _EVAL_163;
  assign _EVAL_148 = _EVAL == _EVAL_149;
  assign _EVAL_48 = _EVAL_137 & _EVAL_131;
  assign _EVAL_106 = _EVAL_144[0];
  assign _EVAL_62 = ~_EVAL_141;
  assign _EVAL_191 = _EVAL_4 >= 2'h2;
  assign _EVAL_121 = _EVAL_6 & _EVAL_37;
  assign _EVAL_115 = 1024'h1 << _EVAL_13;
  assign _EVAL_187 = _EVAL_2 <= 3'h4;
  assign _EVAL_22 = _EVAL_83 | 2'h1;
  assign _EVAL_181 = _EVAL_44 | _EVAL_53;
  assign _EVAL_25 = _EVAL_137 & _EVAL_69;
  assign _EVAL_96 = {{13'd0}, _EVAL_175};
  assign _EVAL_60 = _EVAL_6 & _EVAL_199;
  assign _EVAL_43 = _EVAL_137 & _EVAL_27;
  assign _EVAL_158 = _EVAL_10 == 3'h5;
  assign _EVAL_29 = _EVAL_3 & _EVAL_97;
  assign _EVAL_27 = _EVAL_163 & _EVAL_100;
  assign _EVAL_150 = _EVAL_120[31:0];
  assign _EVAL_172 = _EVAL_49 | _EVAL_82;
  assign _EVAL_97 = ~_EVAL_136;
  assign _EVAL_16 = ~_EVAL_63;
  assign _EVAL_138 = _EVAL_0 ^ 15'h4000;
  assign _EVAL_86 = _EVAL_8 == _EVAL_17;
  assign _EVAL_33 = _EVAL_2 != 3'h0;
  assign _EVAL_88 = _EVAL_19[0];
  assign _EVAL_152 = ~_EVAL_35;
  assign _EVAL_41 = 1024'h1 << _EVAL;
  always @(posedge _EVAL_11) begin
    if (_EVAL_112) begin
      _EVAL_17 <= _EVAL_8;
    end
    if (_EVAL_112) begin
      _EVAL_18 <= _EVAL_13;
    end
    if (_EVAL_112) begin
      _EVAL_28 <= _EVAL_0;
    end
    if (_EVAL_172) begin
      _EVAL_34 <= 32'h0;
    end else begin
      _EVAL_34 <= _EVAL_150;
    end
    if (_EVAL_112) begin
      _EVAL_38 <= _EVAL_5;
    end
    if (_EVAL_49) begin
      if (_EVAL_103) begin
        _EVAL_57 <= 1'h0;
      end else begin
        _EVAL_57 <= _EVAL_88;
      end
    end
    if (_EVAL_64) begin
      _EVAL_65 <= _EVAL_4;
    end
    if (_EVAL_49) begin
      if (_EVAL_204) begin
        _EVAL_68 <= 1'h0;
      end else begin
        _EVAL_68 <= _EVAL_110;
      end
    end
    _EVAL_71 <= _EVAL_182 & _EVAL_152;
    if (_EVAL_64) begin
      _EVAL_79 <= _EVAL_10;
    end
    if (_EVAL_112) begin
      _EVAL_87 <= _EVAL_2;
    end
    if (_EVAL_82) begin
      if (_EVAL_205) begin
        _EVAL_95 <= 1'h0;
      end else begin
        _EVAL_95 <= _EVAL_203;
      end
    end
    if (_EVAL_82) begin
      if (_EVAL_141) begin
        _EVAL_104 <= 1'h0;
      end else begin
        _EVAL_104 <= _EVAL_106;
      end
    end
    if (_EVAL_64) begin
      _EVAL_149 <= _EVAL;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4992fcb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68f0de8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1250331e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42f05e0d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_99) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14285234)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea440944)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8aef1f6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_16) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8508ba8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4348a3fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb0c3d03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db8f96c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77b29a67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce4b5d78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a70f4cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d04add6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c80fd8f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6373ad32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_16) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5dd82052)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b65461b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86a00167)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7378147a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(381f55cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3bbb0705)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(752f86b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_16) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14a349e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94684e51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_99) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32740455)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_145) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0da4c94)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51e5801d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99c4c67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7e50901)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f7d8cce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12926f9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b07bcf4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(372ae319)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63adc1c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b1263b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15b9a388)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1291e9ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28dce979)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4964a82a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6aaf914)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17f2b3d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ad35b23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_146 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed335ed1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e57fedec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_15) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(854cc06f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52145d5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e680afb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3c1e484)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c80fd8f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7db77e7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c779ea9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(677b0de5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c471ac1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e83633c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(633501dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60e7472f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23ed9480)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf3e54df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_16) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(608d9cdc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17cd8959)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f46c9e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_15) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(277764ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70da14fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86e0b1b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48ada1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1024b89f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7e25c49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_9 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e7837df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de9cea5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5faaf7c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb6a23e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_60 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f66f5756)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a80178a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7439c9d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_17 = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_18 = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_28 = _RAND_2[14:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_34 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_38 = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_57 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_65 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_68 = _RAND_7[0:0];
  _RAND_8 = {18{`RANDOM}};
  _EVAL_71 = _RAND_8[575:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_79 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_87 = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_95 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_104 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_149 = _RAND_13[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
