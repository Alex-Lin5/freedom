//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_34_assert(
  input         _EVAL,
  input  [3:0]  _EVAL_0,
  input  [1:0]  _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input  [31:0] _EVAL_10,
  input         _EVAL_11,
  input  [3:0]  _EVAL_12,
  input         _EVAL_13,
  input  [3:0]  _EVAL_14,
  input         _EVAL_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire [32:0] _EVAL_19;
  wire  _EVAL_20;
  wire [32:0] _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire [32:0] _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire [32:0] _EVAL_31;
  wire [6:0] _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire [1:0] _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire [1:0] _EVAL_56;
  wire [32:0] _EVAL_57;
  wire  _EVAL_58;
  wire [32:0] _EVAL_59;
  wire [5:0] _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire [32:0] _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire [32:0] _EVAL_69;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  reg [2:0] _EVAL_76;
  wire  _EVAL_77;
  wire [5:0] _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire [32:0] _EVAL_87;
  wire [3:0] _EVAL_88;
  wire [6:0] _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire [22:0] _EVAL_94;
  wire  _EVAL_95;
  wire [31:0] _EVAL_96;
  wire [5:0] _EVAL_97;
  wire  _EVAL_98;
  wire [32:0] _EVAL_99;
  wire  _EVAL_100;
  wire [6:0] _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire [7:0] _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire [32:0] _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire [32:0] _EVAL_124;
  wire  _EVAL_125;
  reg [3:0] _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire [7:0] _EVAL_134;
  wire  _EVAL_135;
  wire [32:0] _EVAL_136;
  wire [31:0] _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire [3:0] _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire [5:0] _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  reg [5:0] _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  reg [5:0] _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire [1:0] _EVAL_162;
  wire  _EVAL_164;
  wire [31:0] _EVAL_165;
  wire [7:0] _EVAL_166;
  wire [1:0] _EVAL_167;
  reg  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire [32:0] _EVAL_174;
  wire [5:0] _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  reg  _EVAL_182;
  reg [31:0] _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire [31:0] _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire [31:0] _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire [32:0] _EVAL_194;
  wire [7:0] _EVAL_195;
  wire  _EVAL_196;
  reg [5:0] _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire [32:0] _EVAL_200;
  wire  _EVAL_201;
  reg [1:0] _EVAL_202;
  wire  _EVAL_203;
  wire [32:0] _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire [32:0] _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire [31:0] _EVAL_219;
  wire  _EVAL_220;
  reg  _EVAL_221;
  wire  _EVAL_222;
  wire [5:0] _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire [6:0] _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_232;
  reg [3:0] _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire [32:0] _EVAL_238;
  reg  _EVAL_239;
  wire  _EVAL_241;
  wire [32:0] _EVAL_242;
  reg [2:0] _EVAL_243;
  wire  _EVAL_244;
  wire [22:0] _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire [32:0] _EVAL_254;
  wire [32:0] _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  reg [31:0] _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire [32:0] _EVAL_264;
  wire [3:0] _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire [1:0] _EVAL_272;
  wire [31:0] _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire [31:0] _EVAL_277;
  wire [32:0] _EVAL_278;
  wire  _EVAL_279;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_284;
  reg [5:0] _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_292;
  wire  _EVAL_293;
  wire [31:0] _EVAL_294;
  wire  _EVAL_295;
  wire  _EVAL_296;
  wire [31:0] _EVAL_297;
  wire  _EVAL_298;
  wire [32:0] _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire [3:0] _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_304;
  wire  _EVAL_305;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_18 = _EVAL_52 | _EVAL_9;
  assign _EVAL_208 = _EVAL_10 == _EVAL_258;
  assign _EVAL_234 = $signed(_EVAL_19) == 33'sh0;
  assign _EVAL_128 = _EVAL_274 | _EVAL_224;
  assign _EVAL_255 = $signed(_EVAL_21) & -33'sh4000;
  assign _EVAL_194 = $signed(_EVAL_25) & -33'sh1000;
  assign _EVAL_253 = ~_EVAL_267;
  assign _EVAL_20 = _EVAL_269 & _EVAL_259;
  assign _EVAL_92 = _EVAL_269 & _EVAL_284;
  assign _EVAL_122 = _EVAL_15 & _EVAL_72;
  assign _EVAL_293 = _EVAL_277 == 32'h0;
  assign _EVAL_157 = $signed(_EVAL_209) == 33'sh0;
  assign _EVAL_152 = $signed(_EVAL_278) == 33'sh0;
  assign _EVAL_217 = _EVAL_1 != 2'h2;
  assign _EVAL_187 = _EVAL_260 | _EVAL_289;
  assign _EVAL_297 = _EVAL_10 ^ 32'h40000000;
  assign _EVAL_279 = _EVAL_53 & _EVAL_259;
  assign _EVAL_63 = {1'b0,$signed(_EVAL_297)};
  assign _EVAL_186 = _EVAL_71 | _EVAL_170;
  assign _EVAL_74 = _EVAL_260 | _EVAL_151;
  assign _EVAL_68 = $signed(_EVAL_299) == 33'sh0;
  assign _EVAL_86 = ~_EVAL_304;
  assign _EVAL_19 = _EVAL_57;
  assign _EVAL_165 = _EVAL_10 ^ 32'h3000;
  assign _EVAL_96 = _EVAL_10 ^ 32'h20000000;
  assign _EVAL_238 = $signed(_EVAL_69) & -33'sh4000;
  assign _EVAL_78 = _EVAL_89[5:0];
  assign _EVAL_302 = ~_EVAL_265;
  assign _EVAL_90 = _EVAL_0 <= 4'h8;
  assign _EVAL_282 = _EVAL_3 <= 3'h6;
  assign _EVAL_121 = _EVAL_38 | _EVAL_9;
  assign _EVAL_191 = {{24'd0}, _EVAL_166};
  assign _EVAL_35 = _EVAL_181 & _EVAL_154;
  assign _EVAL_61 = ~_EVAL_225;
  assign _EVAL_147 = ~_EVAL_30;
  assign _EVAL_290 = _EVAL_214 | _EVAL_9;
  assign _EVAL_33 = _EVAL_234 | _EVAL_22;
  assign _EVAL_283 = _EVAL_6 == 3'h1;
  assign _EVAL_263 = ~_EVAL_189;
  assign _EVAL_296 = _EVAL_260 | _EVAL_44;
  assign _EVAL_259 = _EVAL_10[0];
  assign _EVAL_300 = _EVAL_0 <= 4'hb;
  assign _EVAL_131 = _EVAL_272[0];
  assign _EVAL_174 = {1'b0,$signed(_EVAL_294)};
  assign _EVAL_16 = ~_EVAL_145;
  assign _EVAL_82 = ~_EVAL_37;
  assign _EVAL_287 = _EVAL_2 & _EVAL_15;
  assign _EVAL_251 = ~_EVAL_305;
  assign _EVAL_249 = _EVAL_139 | _EVAL_9;
  assign _EVAL_44 = _EVAL_123 & _EVAL_275;
  assign _EVAL_203 = _EVAL_15 & _EVAL_58;
  assign _EVAL_28 = ~_EVAL_182;
  assign _EVAL_228 = _EVAL_287 & _EVAL_303;
  assign _EVAL_160 = _EVAL_182 | _EVAL_104;
  assign _EVAL_114 = _EVAL_131 & _EVAL_20;
  assign _EVAL_151 = _EVAL_123 & _EVAL_48;
  assign _EVAL_84 = _EVAL_131 & _EVAL_279;
  assign _EVAL_212 = _EVAL_274 | _EVAL_157;
  assign _EVAL_49 = _EVAL_159 == 6'h0;
  assign _EVAL_142 = _EVAL_244 | _EVAL_9;
  assign _EVAL_37 = _EVAL_206 | _EVAL_9;
  assign _EVAL_303 = _EVAL_285 == 6'h0;
  assign _EVAL_87 = {1'b0,$signed(_EVAL_96)};
  assign _EVAL_104 = _EVAL_56[0];
  assign _EVAL_26 = ~_EVAL_129;
  assign _EVAL_71 = _EVAL_246 | _EVAL_158;
  assign _EVAL_62 = _EVAL_153 == 6'h0;
  assign _EVAL_219 = _EVAL_10 ^ 32'hc000000;
  assign _EVAL_94 = 23'hff << _EVAL_12;
  assign _EVAL_248 = _EVAL_53 & _EVAL_284;
  assign _EVAL_273 = _EVAL_10 ^ 32'h80000000;
  assign _EVAL_272 = _EVAL_45 | 2'h1;
  assign _EVAL_214 = _EVAL == _EVAL_221;
  assign _EVAL_230 = _EVAL_217 | _EVAL_9;
  assign _EVAL_32 = _EVAL_153 - 6'h1;
  assign _EVAL_45 = 2'h1 << _EVAL_150;
  assign _EVAL_124 = _EVAL_183 + 32'h1;
  assign _EVAL_116 = ~_EVAL_34;
  assign _EVAL_173 = ~_EVAL_270;
  assign _EVAL_220 = ~_EVAL_250;
  assign _EVAL_222 = _EVAL_3[0];
  assign _EVAL_31 = $signed(_EVAL_174) & -33'sh10000;
  assign _EVAL_289 = _EVAL_123 & _EVAL_128;
  assign _EVAL_54 = ~_EVAL_142;
  assign _EVAL_79 = _EVAL_71 | _EVAL_114;
  assign _EVAL_39 = _EVAL_8 & _EVAL_80;
  assign _EVAL_64 = _EVAL_199 | _EVAL_9;
  assign _EVAL_55 = _EVAL_8 & _EVAL_81;
  assign _EVAL_278 = _EVAL_264;
  assign _EVAL_295 = _EVAL_15 & _EVAL_262;
  assign _EVAL_129 = _EVAL_28 | _EVAL_9;
  assign _EVAL_42 = ~_EVAL_73;
  assign _EVAL_41 = ~_EVAL_9;
  assign _EVAL_274 = _EVAL_216 | _EVAL_152;
  assign _EVAL_29 = _EVAL_15 & _EVAL_301;
  assign _EVAL_181 = _EVAL_127 & _EVAL_49;
  assign _EVAL_178 = ~_EVAL_193;
  assign _EVAL_51 = _EVAL_6 == 3'h5;
  assign _EVAL_193 = _EVAL_95 | _EVAL_9;
  assign _EVAL_246 = _EVAL_0 >= 4'h2;
  assign _EVAL_72 = ~_EVAL_62;
  assign _EVAL_275 = _EVAL_257 | _EVAL_224;
  assign _EVAL_83 = _EVAL_23 | _EVAL_9;
  assign _EVAL_46 = _EVAL_210 >> _EVAL;
  assign _EVAL_271 = ~_EVAL;
  assign _EVAL_244 = _EVAL_3 == _EVAL_243;
  assign _EVAL_134 = _EVAL_245[7:0];
  assign _EVAL_73 = _EVAL_300 | _EVAL_9;
  assign _EVAL_22 = $signed(_EVAL_118) == 33'sh0;
  assign _EVAL_288 = ~_EVAL_149;
  assign _EVAL_245 = 23'hff << _EVAL_0;
  assign _EVAL_101 = _EVAL_197 - 6'h1;
  assign _EVAL_132 = ~_EVAL_227;
  assign _EVAL_148 = _EVAL_226[5:0];
  assign _EVAL_211 = _EVAL_162[0];
  assign _EVAL_209 = _EVAL_136;
  assign _EVAL_195 = _EVAL_94[7:0];
  assign _EVAL_223 = _EVAL_101[5:0];
  assign _EVAL_185 = _EVAL_1 == _EVAL_202;
  assign _EVAL_117 = _EVAL_272[1];
  assign _EVAL_150 = _EVAL_0[0];
  assign _EVAL_136 = $signed(_EVAL_87) & -33'sh2000;
  assign _EVAL_141 = _EVAL_1 == 2'h0;
  assign _EVAL_48 = _EVAL_157 | _EVAL_115;
  assign _EVAL_250 = _EVAL_17 | _EVAL_9;
  assign _EVAL_77 = _EVAL_0 == _EVAL_233;
  assign _EVAL_267 = _EVAL_247 | _EVAL_9;
  assign _EVAL_91 = _EVAL_199 | _EVAL_7;
  assign _EVAL_88 = _EVAL_14 & _EVAL_302;
  assign _EVAL_266 = _EVAL_141 | _EVAL_9;
  assign _EVAL_89 = _EVAL_285 - 6'h1;
  assign _EVAL_130 = ~_EVAL_211;
  assign _EVAL_57 = $signed(_EVAL_254) & -33'sh5000;
  assign _EVAL_265 = {_EVAL_110,_EVAL_27,_EVAL_79,_EVAL_186};
  assign _EVAL_107 = ~_EVAL_195;
  assign _EVAL_167 = 2'h1 << _EVAL;
  assign _EVAL_115 = $signed(_EVAL_204) == 33'sh0;
  assign _EVAL_127 = _EVAL_5 & _EVAL_8;
  assign _EVAL_286 = _EVAL_169 | _EVAL_9;
  assign _EVAL_25 = {1'b0,$signed(_EVAL_165)};
  assign _EVAL_102 = _EVAL_15 & _EVAL_105;
  assign _EVAL_260 = _EVAL_90 & _EVAL_68;
  assign _EVAL_149 = _EVAL_185 | _EVAL_9;
  assign _EVAL_65 = ~_EVAL_111;
  assign _EVAL_305 = _EVAL_46 | _EVAL_9;
  assign _EVAL_111 = |_EVAL_104;
  assign _EVAL_162 = _EVAL_35 ? _EVAL_167 : 2'h0;
  assign _EVAL_67 = _EVAL_74 | _EVAL_9;
  assign _EVAL_81 = _EVAL_3 == 3'h6;
  assign _EVAL_180 = _EVAL_276 | _EVAL_236;
  assign _EVAL_270 = _EVAL_296 | _EVAL_9;
  assign _EVAL_176 = ~_EVAL_249;
  assign _EVAL_207 = |_EVAL_182;
  assign _EVAL_69 = {1'b0,$signed(_EVAL_273)};
  assign _EVAL_23 = _EVAL_138 | _EVAL_65;
  assign _EVAL_171 = _EVAL_15 & _EVAL_283;
  assign _EVAL_256 = _EVAL_3 == 3'h2;
  assign _EVAL_125 = _EVAL_8 & _EVAL_256;
  assign _EVAL_140 = _EVAL_13 == _EVAL_239;
  assign _EVAL_225 = _EVAL_77 | _EVAL_9;
  assign _EVAL_299 = _EVAL_194;
  assign _EVAL_210 = _EVAL_104 | _EVAL_182;
  assign _EVAL_146 = ~_EVAL_172;
  assign _EVAL_192 = _EVAL_131 & _EVAL_248;
  assign _EVAL_105 = _EVAL_6 == 3'h6;
  assign _EVAL_206 = _EVAL_4 == _EVAL_168;
  assign _EVAL_232 = _EVAL_271 | _EVAL_9;
  assign _EVAL_277 = _EVAL_10 & _EVAL_191;
  assign _EVAL_103 = ~_EVAL_286;
  assign _EVAL_80 = _EVAL_3 == 3'h1;
  assign _EVAL_205 = _EVAL_3 == 3'h4;
  assign _EVAL_120 = _EVAL_117 & _EVAL_53;
  assign _EVAL_254 = {1'b0,$signed(_EVAL_10)};
  assign _EVAL_175 = _EVAL_107[7:2];
  assign _EVAL_172 = _EVAL_282 | _EVAL_9;
  assign _EVAL_247 = _EVAL_12 >= 4'h2;
  assign _EVAL_298 = ~_EVAL_67;
  assign _EVAL_196 = ~_EVAL_232;
  assign _EVAL_301 = _EVAL_6 == 3'h2;
  assign _EVAL_200 = $signed(_EVAL_63) & -33'sh2000;
  assign _EVAL_224 = $signed(_EVAL_242) == 33'sh0;
  assign _EVAL_264 = $signed(_EVAL_59) & -33'sh400000;
  assign _EVAL_237 = _EVAL_8 & _EVAL_205;
  assign _EVAL_166 = ~_EVAL_134;
  assign _EVAL_113 = _EVAL_187 | _EVAL_9;
  assign _EVAL_154 = ~_EVAL_81;
  assign _EVAL_179 = $signed(_EVAL_99) == 33'sh0;
  assign _EVAL_268 = _EVAL_8 & _EVAL_184;
  assign _EVAL_294 = _EVAL_10 ^ 32'h2000000;
  assign _EVAL_145 = _EVAL_6[2];
  assign _EVAL_262 = _EVAL_6 == 3'h7;
  assign _EVAL_235 = ~_EVAL_177;
  assign _EVAL_177 = _EVAL_164 | _EVAL_9;
  assign _EVAL_58 = _EVAL_6 == 3'h4;
  assign _EVAL_284 = ~_EVAL_259;
  assign _EVAL_198 = ~_EVAL_229;
  assign _EVAL_269 = ~_EVAL_53;
  assign _EVAL_201 = _EVAL_208 | _EVAL_9;
  assign _EVAL_27 = _EVAL_144 | _EVAL_192;
  assign _EVAL_137 = _EVAL_10 ^ 32'h1800000;
  assign _EVAL_119 = _EVAL_15 & _EVAL_133;
  assign _EVAL_118 = _EVAL_255;
  assign _EVAL_85 = ~_EVAL_230;
  assign _EVAL_170 = _EVAL_131 & _EVAL_92;
  assign _EVAL_226 = _EVAL_159 - 6'h1;
  assign _EVAL_218 = _EVAL_140 | _EVAL_9;
  assign _EVAL_52 = _EVAL_88 == 4'h0;
  assign _EVAL_161 = ~_EVAL_218;
  assign _EVAL_43 = _EVAL_8 & _EVAL_198;
  assign _EVAL_227 = _EVAL_91 | _EVAL_9;
  assign _EVAL_123 = _EVAL_0 <= 4'h6;
  assign _EVAL_215 = _EVAL_8 & _EVAL_156;
  assign _EVAL_138 = _EVAL_104 != _EVAL_211;
  assign _EVAL_276 = _EVAL_112 | _EVAL_155;
  assign _EVAL_133 = _EVAL_6 == 3'h3;
  assign _EVAL_252 = _EVAL_15 & _EVAL_213;
  assign _EVAL_304 = _EVAL_246 | _EVAL_9;
  assign _EVAL_143 = ~_EVAL_14;
  assign _EVAL_135 = _EVAL_127 & _EVAL_229;
  assign _EVAL_47 = ~_EVAL_113;
  assign _EVAL_53 = _EVAL_10[1];
  assign _EVAL_112 = ~_EVAL_207;
  assign _EVAL_241 = ~_EVAL_201;
  assign _EVAL_38 = _EVAL_12 == _EVAL_126;
  assign _EVAL_156 = _EVAL_3 == 3'h0;
  assign _EVAL_21 = {1'b0,$signed(_EVAL_137)};
  assign _EVAL_199 = ~_EVAL_4;
  assign _EVAL_292 = ~_EVAL_7;
  assign _EVAL_95 = _EVAL_6 == _EVAL_76;
  assign _EVAL_56 = _EVAL_228 ? 2'h1 : 2'h0;
  assign _EVAL_30 = _EVAL_293 | _EVAL_9;
  assign _EVAL_17 = _EVAL_1 <= 2'h2;
  assign _EVAL_155 = plusarg_reader_out == 32'h0;
  assign _EVAL_106 = _EVAL_15 & _EVAL_51;
  assign _EVAL_139 = _EVAL_300 & _EVAL_296;
  assign _EVAL_99 = _EVAL_31;
  assign _EVAL_229 = _EVAL_197 == 6'h0;
  assign _EVAL_216 = _EVAL_33 | _EVAL_179;
  assign _EVAL_34 = _EVAL_292 | _EVAL_9;
  assign _EVAL_60 = _EVAL_32[5:0];
  assign _EVAL_24 = ~_EVAL_64;
  assign _EVAL_144 = _EVAL_246 | _EVAL_120;
  assign _EVAL_281 = _EVAL_287 | _EVAL_127;
  assign _EVAL_36 = ~_EVAL_121;
  assign _EVAL_242 = _EVAL_238;
  assign _EVAL_158 = _EVAL_117 & _EVAL_269;
  assign _EVAL_100 = ~_EVAL_83;
  assign _EVAL_109 = ~_EVAL_266;
  assign _EVAL_108 = ~_EVAL_290;
  assign _EVAL_190 = _EVAL_160 & _EVAL_130;
  assign _EVAL_98 = ~_EVAL_18;
  assign _EVAL_257 = _EVAL_212 | _EVAL_115;
  assign _EVAL_169 = _EVAL_143 == 4'h0;
  assign _EVAL_184 = _EVAL_3 == 3'h5;
  assign _EVAL_164 = _EVAL_14 == _EVAL_265;
  assign _EVAL_189 = _EVAL_180 | _EVAL_9;
  assign _EVAL_50 = _EVAL_287 & _EVAL_62;
  assign _EVAL_213 = _EVAL_6 == 3'h0;
  assign _EVAL_236 = _EVAL_183 < plusarg_reader_out;
  assign _EVAL_97 = _EVAL_166[7:2];
  assign _EVAL_110 = _EVAL_144 | _EVAL_84;
  assign _EVAL_188 = _EVAL_124[31:0];
  assign _EVAL_204 = _EVAL_200;
  assign _EVAL_59 = {1'b0,$signed(_EVAL_219)};
  always @(posedge _EVAL_11) begin
    if (_EVAL_50) begin
      _EVAL_76 <= _EVAL_6;
    end
    if (_EVAL_135) begin
      _EVAL_126 <= _EVAL_12;
    end
    if (_EVAL_9) begin
      _EVAL_153 <= 6'h0;
    end else if (_EVAL_287) begin
      if (_EVAL_62) begin
        if (_EVAL_16) begin
          _EVAL_153 <= _EVAL_97;
        end else begin
          _EVAL_153 <= 6'h0;
        end
      end else begin
        _EVAL_153 <= _EVAL_60;
      end
    end
    if (_EVAL_9) begin
      _EVAL_159 <= 6'h0;
    end else if (_EVAL_127) begin
      if (_EVAL_49) begin
        if (_EVAL_222) begin
          _EVAL_159 <= _EVAL_175;
        end else begin
          _EVAL_159 <= 6'h0;
        end
      end else begin
        _EVAL_159 <= _EVAL_148;
      end
    end
    if (_EVAL_135) begin
      _EVAL_168 <= _EVAL_4;
    end
    if (_EVAL_9) begin
      _EVAL_182 <= 1'h0;
    end else begin
      _EVAL_182 <= _EVAL_190;
    end
    if (_EVAL_9) begin
      _EVAL_183 <= 32'h0;
    end else if (_EVAL_281) begin
      _EVAL_183 <= 32'h0;
    end else begin
      _EVAL_183 <= _EVAL_188;
    end
    if (_EVAL_9) begin
      _EVAL_197 <= 6'h0;
    end else if (_EVAL_127) begin
      if (_EVAL_229) begin
        if (_EVAL_222) begin
          _EVAL_197 <= _EVAL_175;
        end else begin
          _EVAL_197 <= 6'h0;
        end
      end else begin
        _EVAL_197 <= _EVAL_223;
      end
    end
    if (_EVAL_135) begin
      _EVAL_202 <= _EVAL_1;
    end
    if (_EVAL_135) begin
      _EVAL_221 <= _EVAL;
    end
    if (_EVAL_50) begin
      _EVAL_233 <= _EVAL_0;
    end
    if (_EVAL_135) begin
      _EVAL_239 <= _EVAL_13;
    end
    if (_EVAL_135) begin
      _EVAL_243 <= _EVAL_3;
    end
    if (_EVAL_50) begin
      _EVAL_258 <= _EVAL_10;
    end
    if (_EVAL_9) begin
      _EVAL_285 <= 6'h0;
    end else if (_EVAL_287) begin
      if (_EVAL_303) begin
        if (_EVAL_16) begin
          _EVAL_285 <= _EVAL_97;
        end else begin
          _EVAL_285 <= 6'h0;
        end
      end else begin
        _EVAL_285 <= _EVAL_78;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(240f3421)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c886522c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae9c2c1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f31dc89a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f228a42a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_176) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a4d40f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(287601d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9cdb0f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c07cb8fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(555b5fa1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_253) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_253) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5829d37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cab1b99a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d33c048d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c977e216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3db4093)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d60a7991)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ca7b265)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_253) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b4fe685)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_8 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_253) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce2c57fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_298) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(342988c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8afa1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb19176f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9069ee19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(981a2cc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80c029a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95a12441)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_8 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7441aad7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de73524a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abff9cb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_253) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b64abe30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8cd9d0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_253) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8429e093)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b188c6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92950ccb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_176) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea45eb62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e48e9e5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d77c196)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67231e2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c6e6c3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80b61aa2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1c46704)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b55a6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa0869c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(146900f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9069ee19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a80ec9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_288) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fe4dbc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11d1c048)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd9fdb1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_298) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30e59343)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a68f00a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dda8dbe9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_132) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4828ef41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7084525a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b60677c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41e90c39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(904f41b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5dba74f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21544bdc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfbe4a9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bbd9ba3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_119 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ae7cbf7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f054a5f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7a1c171)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65012bad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a95ae53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfe2cc2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(828b4291)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77802b01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_237 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_288) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93888f86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd636fca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_39 & _EVAL_132) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af1d0d10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_76 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_126 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_153 = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_159 = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_168 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_182 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_183 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_197 = _RAND_7[5:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_202 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_221 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_233 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_239 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_243 = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_258 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_285 = _RAND_14[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
