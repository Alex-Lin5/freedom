//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_169(
  output        _EVAL,
  input  [31:0] _EVAL_0,
  input         _EVAL_1,
  output [1:0]  _EVAL_2,
  input  [2:0]  _EVAL_3,
  output        _EVAL_4,
  input         _EVAL_5,
  output [8:0]  _EVAL_6,
  output [2:0]  _EVAL_7,
  output        _EVAL_8,
  output        _EVAL_9,
  input         _EVAL_10,
  input  [2:0]  _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  output        _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  output [31:0] _EVAL_17,
  input  [1:0]  _EVAL_18,
  input  [8:0]  _EVAL_19,
  output        _EVAL_20,
  output        _EVAL_21,
  output [1:0]  _EVAL_22,
  output [31:0] _EVAL_23,
  output        _EVAL_24,
  output [2:0]  _EVAL_25,
  input  [31:0] _EVAL_26
);
  wire  bundleIn_0_d_sink__EVAL;
  wire  bundleIn_0_d_sink__EVAL_0;
  wire  bundleIn_0_d_sink__EVAL_1;
  wire  bundleIn_0_d_sink__EVAL_2;
  wire [1:0] bundleIn_0_d_sink__EVAL_3;
  wire  bundleIn_0_d_sink__EVAL_4;
  wire [31:0] bundleIn_0_d_sink__EVAL_5;
  wire [2:0] bundleIn_0_d_sink__EVAL_6;
  wire  bundleIn_0_d_sink__EVAL_7;
  wire  bundleIn_0_d_sink__EVAL_8;
  wire  bundleIn_0_d_sink__EVAL_9;
  wire [1:0] bundleIn_0_d_sink__EVAL_10;
  wire  bundleIn_0_d_sink__EVAL_11;
  wire [1:0] bundleIn_0_d_sink__EVAL_12;
  wire [31:0] bundleIn_0_d_sink__EVAL_13;
  wire  bundleIn_0_d_sink__EVAL_14;
  wire [2:0] bundleIn_0_d_sink__EVAL_15;
  wire  bundleIn_0_d_sink__EVAL_16;
  wire [2:0] bundleOut_0_a_source__EVAL;
  wire  bundleOut_0_a_source__EVAL_0;
  wire  bundleOut_0_a_source__EVAL_1;
  wire [2:0] bundleOut_0_a_source__EVAL_2;
  wire  bundleOut_0_a_source__EVAL_3;
  wire [31:0] bundleOut_0_a_source__EVAL_4;
  wire [31:0] bundleOut_0_a_source__EVAL_5;
  wire  bundleOut_0_a_source__EVAL_6;
  wire [8:0] bundleOut_0_a_source__EVAL_7;
  wire [8:0] bundleOut_0_a_source__EVAL_8;
  wire  bundleOut_0_a_source__EVAL_9;
  wire  bundleOut_0_a_source__EVAL_10;
  _EVAL_168 bundleIn_0_d_sink (
    ._EVAL(bundleIn_0_d_sink__EVAL),
    ._EVAL_0(bundleIn_0_d_sink__EVAL_0),
    ._EVAL_1(bundleIn_0_d_sink__EVAL_1),
    ._EVAL_2(bundleIn_0_d_sink__EVAL_2),
    ._EVAL_3(bundleIn_0_d_sink__EVAL_3),
    ._EVAL_4(bundleIn_0_d_sink__EVAL_4),
    ._EVAL_5(bundleIn_0_d_sink__EVAL_5),
    ._EVAL_6(bundleIn_0_d_sink__EVAL_6),
    ._EVAL_7(bundleIn_0_d_sink__EVAL_7),
    ._EVAL_8(bundleIn_0_d_sink__EVAL_8),
    ._EVAL_9(bundleIn_0_d_sink__EVAL_9),
    ._EVAL_10(bundleIn_0_d_sink__EVAL_10),
    ._EVAL_11(bundleIn_0_d_sink__EVAL_11),
    ._EVAL_12(bundleIn_0_d_sink__EVAL_12),
    ._EVAL_13(bundleIn_0_d_sink__EVAL_13),
    ._EVAL_14(bundleIn_0_d_sink__EVAL_14),
    ._EVAL_15(bundleIn_0_d_sink__EVAL_15),
    ._EVAL_16(bundleIn_0_d_sink__EVAL_16)
  );
  _EVAL_166 bundleOut_0_a_source (
    ._EVAL(bundleOut_0_a_source__EVAL),
    ._EVAL_0(bundleOut_0_a_source__EVAL_0),
    ._EVAL_1(bundleOut_0_a_source__EVAL_1),
    ._EVAL_2(bundleOut_0_a_source__EVAL_2),
    ._EVAL_3(bundleOut_0_a_source__EVAL_3),
    ._EVAL_4(bundleOut_0_a_source__EVAL_4),
    ._EVAL_5(bundleOut_0_a_source__EVAL_5),
    ._EVAL_6(bundleOut_0_a_source__EVAL_6),
    ._EVAL_7(bundleOut_0_a_source__EVAL_7),
    ._EVAL_8(bundleOut_0_a_source__EVAL_8),
    ._EVAL_9(bundleOut_0_a_source__EVAL_9),
    ._EVAL_10(bundleOut_0_a_source__EVAL_10)
  );
  assign _EVAL_25 = bundleIn_0_d_sink__EVAL_15;
  assign bundleOut_0_a_source__EVAL_8 = _EVAL_19;
  assign _EVAL_7 = bundleOut_0_a_source__EVAL_2;
  assign bundleOut_0_a_source__EVAL_6 = _EVAL_12;
  assign bundleIn_0_d_sink__EVAL_13 = _EVAL_26;
  assign bundleOut_0_a_source__EVAL_4 = _EVAL_0;
  assign bundleIn_0_d_sink__EVAL_2 = _EVAL_12;
  assign bundleIn_0_d_sink__EVAL_6 = _EVAL_3;
  assign _EVAL_9 = bundleIn_0_d_sink__EVAL_14;
  assign bundleOut_0_a_source__EVAL_3 = _EVAL_10;
  assign bundleIn_0_d_sink__EVAL_16 = _EVAL_16;
  assign bundleOut_0_a_source__EVAL_1 = _EVAL_5;
  assign _EVAL_24 = bundleOut_0_a_source__EVAL_10;
  assign _EVAL_21 = bundleOut_0_a_source__EVAL_0;
  assign bundleIn_0_d_sink__EVAL_3 = _EVAL_18;
  assign _EVAL_20 = bundleIn_0_d_sink__EVAL_11;
  assign _EVAL_14 = bundleIn_0_d_sink__EVAL_9;
  assign _EVAL_22 = bundleIn_0_d_sink__EVAL_12;
  assign _EVAL_6 = bundleOut_0_a_source__EVAL_7;
  assign _EVAL_4 = bundleIn_0_d_sink__EVAL_7;
  assign _EVAL_17 = bundleIn_0_d_sink__EVAL_5;
  assign bundleIn_0_d_sink__EVAL_8 = _EVAL_1;
  assign bundleOut_0_a_source__EVAL = _EVAL_11;
  assign _EVAL_2 = bundleIn_0_d_sink__EVAL_10;
  assign bundleIn_0_d_sink__EVAL_4 = _EVAL_5;
  assign _EVAL_8 = bundleIn_0_d_sink__EVAL;
  assign _EVAL_23 = bundleOut_0_a_source__EVAL_5;
  assign _EVAL = bundleIn_0_d_sink__EVAL_1;
  assign bundleOut_0_a_source__EVAL_9 = _EVAL_15;
  assign bundleIn_0_d_sink__EVAL_0 = _EVAL_13;
endmodule
