//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_160_assert(
  input          _EVAL,
  input          _EVAL_0,
  input  [2:0]   _EVAL_1,
  input  [2:0]   _EVAL_2,
  input          _EVAL_3,
  input          _EVAL_4,
  input  [127:0] _EVAL_5,
  input          _EVAL_6,
  input          _EVAL_7,
  input          _EVAL_8
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_9;
  wire  _EVAL_10;
  wire  _EVAL_11;
  wire  _EVAL_12;
  wire [1:0] _EVAL_13;
  wire  _EVAL_14;
  wire  _EVAL_15;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  reg [2:0] _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  reg  _EVAL_32;
  wire [127:0] _EVAL_33;
  wire  _EVAL_34;
  wire [32:0] _EVAL_35;
  wire  _EVAL_36;
  wire [1:0] _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire [1:0] _EVAL_49;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire [128:0] _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  reg [127:0] _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire [128:0] _EVAL_76;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire [1:0] _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  reg  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire [1:0] _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  reg [31:0] _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire [128:0] _EVAL_96;
  reg  _EVAL_97;
  wire [31:0] _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire [1:0] _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  reg  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  reg  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  reg [2:0] _EVAL_125;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_119 = _EVAL_117 | _EVAL_41;
  assign _EVAL_17 = _EVAL_8 & _EVAL_59;
  assign _EVAL_19 = ~_EVAL_86;
  assign _EVAL_46 = _EVAL_8 & _EVAL_62;
  assign _EVAL_59 = _EVAL_2 == 3'h2;
  assign _EVAL_72 = _EVAL_8 & _EVAL_44;
  assign _EVAL_123 = _EVAL_2 == 3'h5;
  assign _EVAL_63 = _EVAL_1 <= 3'h6;
  assign _EVAL_35 = _EVAL_92 + 32'h1;
  assign _EVAL_47 = _EVAL_7 & _EVAL_112;
  assign _EVAL_107 = |_EVAL_115;
  assign _EVAL_102 = _EVAL_4 & _EVAL_7;
  assign _EVAL_12 = _EVAL_39 & _EVAL_82;
  assign _EVAL_18 = _EVAL_9 & _EVAL_23;
  assign _EVAL_41 = _EVAL_92 < plusarg_reader_out;
  assign _EVAL_90 = _EVAL_8 & _EVAL_21;
  assign _EVAL_24 = _EVAL_58 | _EVAL_61;
  assign _EVAL_94 = _EVAL_49[0];
  assign _EVAL_21 = _EVAL_2 == 3'h0;
  assign _EVAL_56 = _EVAL_2 == _EVAL_125;
  assign _EVAL_13 = _EVAL_32 - 1'h1;
  assign _EVAL_89 = _EVAL_18 ? 2'h1 : 2'h0;
  assign _EVAL_70 = ~_EVAL_87;
  assign _EVAL_44 = _EVAL_2 == 3'h1;
  assign _EVAL_122 = ~_EVAL_116;
  assign _EVAL_112 = _EVAL_1 == 3'h1;
  assign _EVAL_58 = ~_EVAL_115;
  assign _EVAL_50 = ~_EVAL_93;
  assign _EVAL_74 = ~_EVAL_24;
  assign _EVAL_34 = ~_EVAL_109;
  assign _EVAL_111 = _EVAL_1 == _EVAL_20;
  assign _EVAL_88 = _EVAL_8 & _EVAL_113;
  assign _EVAL_121 = _EVAL_7 & _EVAL_54;
  assign _EVAL_57 = ~_EVAL_106;
  assign _EVAL_76 = $signed(_EVAL_96) & 129'sh100000000000000000000000000000000;
  assign _EVAL_51 = _EVAL_8 & _EVAL_100;
  assign _EVAL_99 = plusarg_reader_out == 32'h0;
  assign _EVAL_96 = {1'b0,$signed(_EVAL_5)};
  assign _EVAL_54 = _EVAL_1 == 3'h6;
  assign _EVAL_52 = _EVAL_7 & _EVAL_26;
  assign _EVAL_38 = ~_EVAL_32;
  assign _EVAL_66 = _EVAL_7 & _EVAL_55;
  assign _EVAL_108 = _EVAL_8 & _EVAL_79;
  assign _EVAL_82 = ~_EVAL_97;
  assign _EVAL_62 = _EVAL_2 == 3'h3;
  assign _EVAL_23 = ~_EVAL_54;
  assign _EVAL_100 = _EVAL_2 == 3'h4;
  assign _EVAL_61 = _EVAL_3;
  assign _EVAL_48 = _EVAL_1 == 3'h2;
  assign _EVAL_25 = ~_EVAL_40;
  assign _EVAL_16 = _EVAL_71 | _EVAL_61;
  assign _EVAL_87 = _EVAL_89[0];
  assign _EVAL_40 = _EVAL_111 | _EVAL_61;
  assign _EVAL_69 = _EVAL_8 & _EVAL_91;
  assign _EVAL_98 = _EVAL_35[31:0];
  assign _EVAL_75 = ~_EVAL_107;
  assign _EVAL_28 = _EVAL_63 | _EVAL_61;
  assign _EVAL_109 = _EVAL_95 | _EVAL_61;
  assign _EVAL_39 = _EVAL_6 & _EVAL_8;
  assign _EVAL_117 = _EVAL_75 | _EVAL_99;
  assign _EVAL_37 = _EVAL_86 - 1'h1;
  assign _EVAL_71 = _EVAL_94 | _EVAL_115;
  assign _EVAL_55 = _EVAL_1 == 3'h5;
  assign _EVAL_30 = _EVAL_37[0];
  assign _EVAL_9 = _EVAL_102 & _EVAL_38;
  assign _EVAL_27 = ~_EVAL_61;
  assign _EVAL_110 = _EVAL | _EVAL_61;
  assign _EVAL_104 = _EVAL_7 & _EVAL_45;
  assign _EVAL_120 = _EVAL_39 & _EVAL_19;
  assign _EVAL_79 = ~_EVAL_82;
  assign _EVAL_95 = $signed(_EVAL_64) == 129'sh0;
  assign _EVAL_65 = _EVAL_5 == _EVAL_67;
  assign _EVAL_85 = ~_EVAL;
  assign _EVAL_10 = _EVAL_65 | _EVAL_61;
  assign _EVAL_101 = _EVAL_97 - 1'h1;
  assign _EVAL_105 = _EVAL_102 & _EVAL_57;
  assign _EVAL_29 = _EVAL_13[0];
  assign _EVAL_68 = _EVAL_7 & _EVAL_48;
  assign _EVAL_42 = ~_EVAL_110;
  assign _EVAL_93 = _EVAL_119 | _EVAL_61;
  assign _EVAL_53 = ~_EVAL_28;
  assign _EVAL_83 = ~_EVAL_103;
  assign _EVAL_80 = _EVAL_81[0];
  assign _EVAL_22 = _EVAL_33 == 128'h0;
  assign _EVAL_113 = _EVAL_2 == 3'h7;
  assign _EVAL_84 = ~_EVAL_10;
  assign _EVAL_33 = _EVAL_5 & 128'h3;
  assign _EVAL_103 = _EVAL_22 | _EVAL_61;
  assign _EVAL_78 = ~_EVAL_31;
  assign _EVAL_15 = ~_EVAL_57;
  assign _EVAL_81 = _EVAL_106 - 1'h1;
  assign _EVAL_45 = _EVAL_1 == 3'h0;
  assign _EVAL_118 = _EVAL_7 & _EVAL_15;
  assign _EVAL_14 = _EVAL_115 | _EVAL_94;
  assign _EVAL_26 = _EVAL_1 == 3'h4;
  assign _EVAL_43 = _EVAL_101[0];
  assign _EVAL_49 = _EVAL_120 ? 2'h1 : 2'h0;
  assign _EVAL_64 = _EVAL_76;
  assign _EVAL_91 = _EVAL_2 == 3'h6;
  assign _EVAL_116 = _EVAL_56 | _EVAL_61;
  assign _EVAL_11 = _EVAL_39 | _EVAL_102;
  assign _EVAL_114 = ~_EVAL_16;
  assign _EVAL_31 = _EVAL_85 | _EVAL_61;
  assign _EVAL_36 = _EVAL_8 & _EVAL_123;
  always @(posedge _EVAL_0) begin
    if (_EVAL_105) begin
      _EVAL_20 <= _EVAL_1;
    end
    if (_EVAL_12) begin
      _EVAL_67 <= _EVAL_5;
    end
    if (_EVAL_12) begin
      _EVAL_125 <= _EVAL_2;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(171706e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49b4c639)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4014bd8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2446c6ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6822fb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b874d27c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc3c277f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_7 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37de5313)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bea34253)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9b7235d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_7 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e62b5139)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a0f6728)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d9d2897)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39ecf749)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5081c815)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8f95875)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfb2a0fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(613f9a50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb05e6a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ce4cfad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3db6fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f34dcfb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56103bac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df0181a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24ad9e71)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad8281b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aae5a385)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a99a083)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3debd2c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd848d92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e02748db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8141b196)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de229173)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be233d4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(575caf48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2446c6ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_46 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a54a6580)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge _EVAL_0 or posedge _EVAL_3) begin
    if (_EVAL_3) begin
      _EVAL_32 <= 1'h0;
    end else if (_EVAL_102) begin
      if (_EVAL_38) begin
        _EVAL_32 <= 1'h0;
      end else begin
        _EVAL_32 <= _EVAL_29;
      end
    end
  end
  always @(posedge _EVAL_0 or posedge _EVAL_3) begin
    if (_EVAL_3) begin
      _EVAL_86 <= 1'h0;
    end else if (_EVAL_39) begin
      if (_EVAL_19) begin
        _EVAL_86 <= 1'h0;
      end else begin
        _EVAL_86 <= _EVAL_30;
      end
    end
  end
  always @(posedge _EVAL_0 or posedge _EVAL_3) begin
    if (_EVAL_3) begin
      _EVAL_92 <= 32'h0;
    end else if (_EVAL_11) begin
      _EVAL_92 <= 32'h0;
    end else begin
      _EVAL_92 <= _EVAL_98;
    end
  end
  always @(posedge _EVAL_0 or posedge _EVAL_3) begin
    if (_EVAL_3) begin
      _EVAL_97 <= 1'h0;
    end else if (_EVAL_39) begin
      if (_EVAL_82) begin
        _EVAL_97 <= 1'h0;
      end else begin
        _EVAL_97 <= _EVAL_43;
      end
    end
  end
  always @(posedge _EVAL_0 or posedge _EVAL_3) begin
    if (_EVAL_3) begin
      _EVAL_106 <= 1'h0;
    end else if (_EVAL_102) begin
      if (_EVAL_57) begin
        _EVAL_106 <= 1'h0;
      end else begin
        _EVAL_106 <= _EVAL_80;
      end
    end
  end
  always @(posedge _EVAL_0 or posedge _EVAL_3) begin
    if (_EVAL_3) begin
      _EVAL_115 <= 1'h0;
    end else begin
      _EVAL_115 <= _EVAL_14 & _EVAL_70;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_20 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_32 = _RAND_1[0:0];
  _RAND_2 = {4{`RANDOM}};
  _EVAL_67 = _RAND_2[127:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_86 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_92 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_97 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_106 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_115 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_125 = _RAND_8[2:0];
`endif // RANDOMIZE_REG_INIT
  if (_EVAL_3) begin
    _EVAL_32 = 1'h0;
  end
  if (_EVAL_3) begin
    _EVAL_86 = 1'h0;
  end
  if (_EVAL_3) begin
    _EVAL_92 = 32'h0;
  end
  if (_EVAL_3) begin
    _EVAL_97 = 1'h0;
  end
  if (_EVAL_3) begin
    _EVAL_106 = 1'h0;
  end
  if (_EVAL_3) begin
    _EVAL_115 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
