//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_177(
  input         _EVAL,
  output [2:0]  _EVAL_0,
  input         _EVAL_1,
  output        _EVAL_2,
  input  [2:0]  _EVAL_3,
  input         _EVAL_4,
  output [3:0]  _EVAL_5,
  input  [9:0]  _EVAL_6,
  output [31:0] _EVAL_7,
  input  [7:0]  _EVAL_8,
  input  [2:0]  _EVAL_9,
  output        _EVAL_10,
  input  [9:0]  _EVAL_11,
  output [2:0]  _EVAL_12,
  output [31:0] _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  output        _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18,
  input         _EVAL_19,
  input         _EVAL_20,
  output [1:0]  _EVAL_21,
  output        _EVAL_22,
  output [7:0]  _EVAL_23,
  output        _EVAL_24,
  output [9:0]  _EVAL_25,
  input  [2:0]  _EVAL_26,
  input  [2:0]  _EVAL_27,
  output        _EVAL_28,
  output [31:0] _EVAL_29,
  input         _EVAL_30,
  input         _EVAL_31,
  input  [3:0]  _EVAL_32,
  input  [1:0]  _EVAL_33,
  input         _EVAL_34,
  input         _EVAL_35,
  input         _EVAL_36,
  output        _EVAL_37,
  input         _EVAL_38,
  input  [31:0] _EVAL_39,
  input  [31:0] _EVAL_40,
  output [1:0]  _EVAL_41,
  input  [8:0]  _EVAL_42,
  input  [3:0]  _EVAL_43,
  input         _EVAL_44,
  input         _EVAL_45,
  output        _EVAL_46,
  output [2:0]  _EVAL_47,
  input         _EVAL_48,
  input  [1:0]  _EVAL_49,
  input         _EVAL_50,
  input         _EVAL_51,
  output        _EVAL_52,
  input         _EVAL_53,
  input  [11:0] _EVAL_54
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_60;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire [7:0] _EVAL_68;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire [31:0] _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_76;
  wire [31:0] _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_86;
  wire [8:0] _EVAL_87;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_92;
  wire  _EVAL_94;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire [31:0] _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_112;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_120;
  wire [31:0] _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire [2:0] _EVAL_129;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire [127:0] _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_137;
  wire [31:0] _EVAL_139;
  wire [127:0] _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_144;
  wire  _EVAL_146;
  wire  _EVAL_148;
  wire  _EVAL_150;
  wire  _EVAL_154;
  wire [1023:0] _EVAL_155;
  wire  _EVAL_156;
  reg [7:0] _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire [31:0] _EVAL_173;
  wire [31:0] _EVAL_174;
  wire  _EVAL_177;
  wire [7:0] _EVAL_178;
  wire [31:0] _EVAL_180;
  wire  _EVAL_182;
  wire  _EVAL_184;
  wire [31:0] _EVAL_186;
  wire  _EVAL_187;
  wire [13:0] _EVAL_188;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_195;
  wire [1023:0] _EVAL_196;
  wire  _EVAL_198;
  reg [31:0] _EVAL_199;
  wire [6:0] _EVAL_200;
  wire  _EVAL_202;
  wire [31:0] _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_213;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_219;
  wire  _EVAL_222;
  wire  _EVAL_223;
  reg  _EVAL_225;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire [31:0] _EVAL_231;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_237;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire [127:0] _EVAL_242;
  wire [31:0] _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire [31:0] _EVAL_252;
  wire [7:0] _EVAL_253;
  wire  _EVAL_258;
  wire [15:0] _EVAL_259;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire [31:0] _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  reg  _EVAL_274;
  wire  _EVAL_276;
  wire  _EVAL_278;
  wire  _EVAL_280;
  wire [31:0] _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire [31:0] _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire [127:0] _EVAL_295;
  wire  _EVAL_296;
  wire  _EVAL_297;
  wire  _EVAL_298;
  wire [31:0] _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_302;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire [2:0] _EVAL_307;
  reg [7:0] _EVAL_308;
  wire  _EVAL_309;
  wire  _EVAL_310;
  wire  _EVAL_311;
  wire [9:0] _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_317;
  wire  _EVAL_319;
  wire  _EVAL_321;
  wire  _EVAL_322;
  reg [7:0] _EVAL_325;
  wire  _EVAL_326;
  wire  _EVAL_327;
  wire  _EVAL_328;
  wire  _EVAL_331;
  wire  _EVAL_332;
  reg [7:0] _EVAL_333;
  wire  _EVAL_334;
  wire  _EVAL_335;
  wire  _EVAL_336;
  wire  _EVAL_337;
  wire  _EVAL_339;
  wire  _EVAL_340;
  wire  _EVAL_341;
  wire  _EVAL_342;
  wire [9:0] _EVAL_343;
  wire  _EVAL_344;
  wire  _EVAL_345;
  wire  _EVAL_346;
  wire [31:0] _EVAL_347;
  wire  _EVAL_348;
  wire [8:0] _EVAL_351;
  wire  _EVAL_352;
  wire  _EVAL_353;
  wire  _EVAL_354;
  wire  _EVAL_356;
  wire  _EVAL_358;
  wire  _EVAL_359;
  wire  _EVAL_360;
  wire  _EVAL_361;
  wire  _EVAL_362;
  wire  _EVAL_363;
  wire  _EVAL_364;
  wire  _EVAL_366;
  wire  _EVAL_367;
  wire  _EVAL_369;
  reg [7:0] _EVAL_372;
  wire  _EVAL_373;
  wire  _EVAL_374;
  wire  _EVAL_375;
  reg [7:0] _EVAL_379;
  wire  hartIsInResetSync_0_debug_hartReset_0__EVAL;
  wire  hartIsInResetSync_0_debug_hartReset_0__EVAL_0;
  wire  hartIsInResetSync_0_debug_hartReset_0__EVAL_1;
  wire  hartIsInResetSync_0_debug_hartReset_0__EVAL_2;
  wire  _EVAL_380;
  wire  _EVAL_382;
  wire [7:0] _EVAL_383;
  reg  _EVAL_385;
  wire  _EVAL_386;
  reg  _EVAL_388;
  wire  _EVAL_389;
  wire [31:0] _EVAL_390;
  wire  _EVAL_391;
  wire  _EVAL_392;
  wire  _EVAL_393;
  wire  _EVAL_395;
  reg [7:0] _EVAL_397;
  wire  _EVAL_400;
  wire [31:0] _EVAL_403;
  wire  _EVAL_407;
  wire  _EVAL_408;
  wire  _EVAL_410;
  wire  _EVAL_411;
  wire  _EVAL_412;
  wire  _EVAL_413;
  wire [31:0] _EVAL_415;
  wire  _EVAL_416;
  wire  _EVAL_417;
  wire  _EVAL_418;
  wire  _EVAL_419;
  wire  _EVAL_420;
  wire  _EVAL_421;
  wire  _EVAL_422;
  wire  _EVAL_423;
  wire  _EVAL_425;
  wire  _EVAL_426;
  wire  _EVAL_427;
  wire [31:0] _EVAL_428;
  wire  _EVAL_429;
  wire [7:0] _EVAL_430;
  wire  _EVAL_432;
  wire  _EVAL_434;
  wire [31:0] _EVAL_436;
  wire  _EVAL_437;
  wire  _EVAL_438;
  wire  _EVAL_439;
  wire [31:0] _EVAL_441;
  wire  _EVAL_443;
  wire  _EVAL_444;
  wire [31:0] _EVAL_445;
  wire  _EVAL_446;
  wire  _EVAL_447;
  reg [7:0] _EVAL_448;
  wire  _EVAL_449;
  wire  _EVAL_450;
  reg [7:0] _EVAL_451;
  wire  _EVAL_453;
  wire  _EVAL_454;
  wire  _EVAL_455;
  wire  _EVAL_456;
  reg [7:0] _EVAL_458;
  wire  _EVAL_460;
  wire  _EVAL_462;
  wire [2:0] _EVAL_463;
  wire  _EVAL_464;
  wire  _EVAL_466;
  wire  _EVAL_467;
  wire  _EVAL_470;
  wire  _EVAL_471;
  wire  _EVAL_472;
  wire  _EVAL_473;
  wire  _EVAL_474;
  wire [2:0] _EVAL_475;
  wire [31:0] _EVAL_476;
  wire  _EVAL_479;
  wire  _EVAL_481;
  wire  _EVAL_482;
  wire  _EVAL_484;
  wire [31:0] _EVAL_485;
  wire  _EVAL_486;
  wire  _EVAL_491;
  wire  _EVAL_494;
  wire  _EVAL_496;
  wire  _EVAL_497;
  wire  _EVAL_498;
  wire  _EVAL_500;
  wire [31:0] _EVAL_501;
  wire  _EVAL_502;
  wire  _EVAL_503;
  wire  _EVAL_504;
  wire  _EVAL_505;
  reg [7:0] _EVAL_506;
  wire  _EVAL_507;
  wire  _EVAL_508;
  wire  _EVAL_510;
  wire  _EVAL_511;
  wire  _EVAL_513;
  wire  _EVAL_515;
  wire  _EVAL_516;
  wire [31:0] _EVAL_517;
  wire  _EVAL_519;
  reg [7:0] _EVAL_520;
  wire  _EVAL_521;
  wire  _EVAL_522;
  wire  _EVAL_523;
  wire  _EVAL_525;
  wire  _EVAL_526;
  wire  _EVAL_528;
  reg [7:0] _EVAL_529;
  wire  _EVAL_530;
  wire  _EVAL_532;
  wire  _EVAL_534;
  wire  _EVAL_535;
  wire  _EVAL_536;
  wire  _EVAL_537;
  wire  _EVAL_538;
  wire [31:0] _EVAL_540;
  wire  _EVAL_541;
  wire  _EVAL_543;
  wire  _EVAL_544;
  reg [7:0] _EVAL_545;
  wire [31:0] _EVAL_546;
  wire  _EVAL_548;
  wire  _EVAL_549;
  wire  _EVAL_550;
  wire  _EVAL_552;
  reg [7:0] _EVAL_553;
  wire [7:0] _EVAL_554;
  wire  _EVAL_555;
  wire  _EVAL_556;
  wire  _EVAL_557;
  wire  _EVAL_559;
  wire [7:0] _EVAL_560;
  wire  _EVAL_561;
  wire  _EVAL_562;
  wire  _EVAL_563;
  wire  _EVAL_564;
  wire  _EVAL_565;
  reg  _EVAL_566;
  wire  _EVAL_567;
  wire  _EVAL_568;
  wire  _EVAL_570;
  wire  _EVAL_572;
  wire  _EVAL_574;
  wire  _EVAL_575;
  wire  _EVAL_577;
  reg [7:0] _EVAL_578;
  wire  _EVAL_585;
  wire [63:0] _EVAL_586;
  wire  _EVAL_589;
  wire [1023:0] _EVAL_591;
  wire  _EVAL_592;
  wire  _EVAL_593;
  wire  _EVAL_595;
  wire  _EVAL_597;
  wire  _EVAL_600;
  wire  _EVAL_601;
  wire [20:0] _EVAL_603;
  wire [2:0] _EVAL_604;
  wire  _EVAL_605;
  reg [7:0] _EVAL_606;
  wire  _EVAL_607;
  wire [11:0] _EVAL_608;
  wire  _EVAL_609;
  wire  _EVAL_610;
  wire  _EVAL_611;
  wire  _EVAL_613;
  wire  _EVAL_614;
  wire  _EVAL_617;
  wire  _EVAL_618;
  wire [31:0] _EVAL_621;
  wire  _EVAL_623;
  reg [7:0] _EVAL_624;
  reg [2:0] _EVAL_625;
  wire  _EVAL_626;
  wire  _EVAL_628;
  wire  _EVAL_629;
  wire  _EVAL_631;
  wire  _EVAL_632;
  wire [7:0] _EVAL_634;
  wire  _EVAL_635;
  wire  _EVAL_636;
  wire  _EVAL_638;
  wire  _EVAL_639;
  wire [7:0] _EVAL_640;
  wire  _EVAL_641;
  wire  _EVAL_642;
  wire  _EVAL_643;
  reg  _EVAL_647;
  wire  _EVAL_648;
  wire  _EVAL_649;
  wire  _EVAL_650;
  wire [7:0] _EVAL_651;
  wire  _EVAL_653;
  wire  _EVAL_654;
  wire [15:0] _EVAL_655;
  wire  _EVAL_658;
  wire  _EVAL_660;
  wire  _EVAL_661;
  reg [7:0] _EVAL_664;
  wire  _EVAL_665;
  wire  _EVAL_666;
  wire  _EVAL_667;
  wire  _EVAL_668;
  wire  _EVAL_669;
  wire  _EVAL_670;
  wire  _EVAL_671;
  wire  _EVAL_673;
  wire  _EVAL_675;
  wire  _EVAL_676;
  wire [127:0] _EVAL_677;
  wire [3:0] _EVAL_678;
  wire  _EVAL_680;
  reg [7:0] _EVAL_684;
  wire  _EVAL_685;
  wire  _EVAL_686;
  wire  _EVAL_687;
  wire  _EVAL_688;
  wire  _EVAL_689;
  wire  _EVAL_690;
  wire  _EVAL_691;
  reg  _EVAL_692;
  wire  _EVAL_694;
  reg [7:0] _EVAL_696;
  wire  _EVAL_698;
  wire  _EVAL_699;
  wire [31:0] _EVAL_700;
  wire [7:0] _EVAL_701;
  wire  _EVAL_702;
  reg [7:0] _EVAL_704;
  wire  _EVAL_705;
  wire  _EVAL_707;
  wire  _EVAL_709;
  wire  _EVAL_710;
  wire  _EVAL_712;
  reg [7:0] _EVAL_713;
  wire  _EVAL_715;
  wire  _EVAL_716;
  wire  _EVAL_717;
  wire  _EVAL_718;
  wire [2:0] _EVAL_723;
  wire  _EVAL_724;
  wire  _EVAL_725;
  wire  _EVAL_726;
  wire  _EVAL_727;
  wire  _EVAL_729;
  wire  _EVAL_732;
  wire  _EVAL_733;
  reg [7:0] _EVAL_735;
  wire [7:0] _EVAL_736;
  wire [9:0] _EVAL_737;
  wire  _EVAL_739;
  wire  _EVAL_740;
  wire [31:0] _EVAL_741;
  wire  _EVAL_742;
  wire  _EVAL_743;
  reg [7:0] _EVAL_744;
  wire  _EVAL_747;
  wire  _EVAL_748;
  reg [7:0] _EVAL_749;
  wire  _EVAL_751;
  wire  _EVAL_753;
  reg [7:0] _EVAL_754;
  wire  _EVAL_755;
  wire [31:0] _EVAL_756;
  wire [31:0] _EVAL_757;
  wire  _EVAL_758;
  wire [31:0] _EVAL_761;
  wire  _EVAL_763;
  wire [7:0] _EVAL_765;
  wire  _EVAL_766;
  wire  _EVAL_767;
  wire  _EVAL_768;
  wire  _EVAL_769;
  wire  _EVAL_772;
  wire  _EVAL_773;
  wire [31:0] _EVAL_775;
  wire  _EVAL_776;
  reg [7:0] _EVAL_777;
  wire  _EVAL_778;
  wire  _EVAL_779;
  wire  _EVAL_781;
  wire [31:0] _EVAL_782;
  wire  _EVAL_783;
  wire  _EVAL_784;
  wire  _EVAL_785;
  wire  _EVAL_787;
  wire  _EVAL_788;
  wire  _EVAL_789;
  wire [31:0] _EVAL_791;
  wire [23:0] _EVAL_793;
  wire [31:0] _EVAL_794;
  wire  _EVAL_797;
  wire  _EVAL_801;
  wire  _EVAL_802;
  wire  _EVAL_803;
  wire  _EVAL_805;
  wire  _EVAL_811;
  wire  _EVAL_813;
  wire  _EVAL_814;
  wire [7:0] _EVAL_815;
  wire  _EVAL_817;
  wire  _EVAL_819;
  wire  _EVAL_821;
  reg [7:0] _EVAL_822;
  wire  _EVAL_823;
  wire  _EVAL_825;
  wire  _EVAL_827;
  wire [31:0] _EVAL_828;
  wire [28:0] _EVAL_830;
  wire  _EVAL_831;
  wire  _EVAL_832;
  wire [31:0] _EVAL_834;
  wire  _EVAL_836;
  wire  _EVAL_837;
  wire  _EVAL_838;
  wire  _EVAL_839;
  wire  _EVAL_841;
  wire  _EVAL_842;
  wire  _EVAL_844;
  wire  _EVAL_845;
  wire  _EVAL_846;
  wire  _EVAL_847;
  wire  _EVAL_848;
  wire  _EVAL_849;
  wire  _EVAL_850;
  wire  _EVAL_852;
  wire  _EVAL_854;
  reg [7:0] _EVAL_855;
  reg [7:0] _EVAL_856;
  wire  _EVAL_857;
  wire  _EVAL_858;
  wire  _EVAL_859;
  wire  _EVAL_861;
  wire [31:0] _EVAL_862;
  wire  _EVAL_863;
  wire  _EVAL_865;
  wire  _EVAL_866;
  wire  _EVAL_867;
  wire  _EVAL_868;
  wire  _EVAL_870;
  wire  _EVAL_871;
  wire  _EVAL_874;
  wire  _EVAL_875;
  wire  _EVAL_876;
  wire  _EVAL_880;
  wire  _EVAL_882;
  wire  _EVAL_883;
  wire  _EVAL_885;
  wire  _EVAL_886;
  wire  _EVAL_887;
  wire  _EVAL_888;
  wire  _EVAL_890;
  wire  _EVAL_891;
  wire  _EVAL_892;
  wire  _EVAL_894;
  wire  _EVAL_895;
  wire  _EVAL_896;
  wire  _EVAL_897;
  wire  _EVAL_898;
  wire  _EVAL_899;
  wire [31:0] _EVAL_901;
  reg [7:0] _EVAL_903;
  wire  _EVAL_904;
  wire [31:0] _EVAL_905;
  wire  _EVAL_906;
  wire  _EVAL_907;
  wire  _EVAL_908;
  wire  _EVAL_910;
  wire  _EVAL_911;
  wire  _EVAL_914;
  wire [31:0] _EVAL_915;
  wire  _EVAL_920;
  wire  _EVAL_921;
  reg [11:0] _EVAL_922;
  wire  _EVAL_923;
  wire  _EVAL_924;
  wire [31:0] _EVAL_925;
  wire [31:0] _EVAL_926;
  wire  _EVAL_927;
  wire  _EVAL_928;
  wire  _EVAL_929;
  wire  _EVAL_933;
  wire  _EVAL_934;
  wire  _EVAL_935;
  wire  _EVAL_936;
  wire [31:0] _EVAL_937;
  wire [9:0] _EVAL_939;
  wire [7:0] _EVAL_940;
  wire  _EVAL_942;
  wire  _EVAL_946;
  wire [7:0] _EVAL_949;
  wire  _EVAL_951;
  wire [31:0] _EVAL_954;
  wire  _EVAL_956;
  wire  _EVAL_957;
  wire  _EVAL_958;
  wire  _EVAL_959;
  wire  _EVAL_961;
  wire  _EVAL_963;
  wire  _EVAL_964;
  wire  _EVAL_966;
  wire [2:0] _EVAL_967;
  wire  _EVAL_968;
  wire [31:0] _EVAL_971;
  wire  _EVAL_972;
  wire  _EVAL_973;
  wire  _EVAL_974;
  wire  _EVAL_975;
  wire  _EVAL_976;
  wire  _EVAL_978;
  wire  _EVAL_979;
  reg [7:0] _EVAL_980;
  wire  _EVAL_981;
  wire  _EVAL_982;
  wire  _EVAL_984;
  wire  _EVAL_986;
  reg [7:0] _EVAL_988;
  wire  _EVAL_989;
  wire  _EVAL_991;
  wire [2:0] _EVAL_992;
  wire  _EVAL_994;
  wire  _EVAL_995;
  wire  _EVAL_996;
  wire  _EVAL_998;
  wire [31:0] _EVAL_999;
  wire [7:0] _EVAL_1000;
  wire  _EVAL_1001;
  wire  _EVAL_1002;
  wire  _EVAL_1007;
  reg [7:0] _EVAL_1008;
  reg [31:0] _EVAL_1009;
  wire  _EVAL_1010;
  reg [7:0] _EVAL_1011;
  wire  _EVAL_1012;
  wire  _EVAL_1013;
  wire  _EVAL_1014;
  wire  _EVAL_1015;
  wire  _EVAL_1016;
  wire  _EVAL_1019;
  wire  _EVAL_1020;
  wire  _EVAL_1022;
  wire  _EVAL_1023;
  wire  _EVAL_1024;
  wire  _EVAL_1025;
  wire  _EVAL_1026;
  wire  _EVAL_1028;
  wire  _EVAL_1030;
  wire  _EVAL_1032;
  wire  _EVAL_1033;
  wire  _EVAL_1035;
  wire  _EVAL_1036;
  wire  _EVAL_1038;
  wire [23:0] _EVAL_1040;
  wire  _EVAL_1042;
  wire  _EVAL_1043;
  wire  _EVAL_1044;
  wire  _EVAL_1045;
  wire  _EVAL_1046;
  wire  _EVAL_1047;
  reg [7:0] _EVAL_1048;
  wire  _EVAL_1050;
  reg [7:0] _EVAL_1051;
  wire  _EVAL_1052;
  wire  _EVAL_1053;
  wire  _EVAL_1054;
  wire  _EVAL_1055;
  wire  _EVAL_1056;
  wire  _EVAL_1057;
  wire  _EVAL_1058;
  wire  _EVAL_1059;
  wire  _EVAL_1061;
  wire  _EVAL_1062;
  reg [7:0] _EVAL_1063;
  wire  _EVAL_1068;
  wire  _EVAL_1070;
  wire  _EVAL_1071;
  wire  _EVAL_1072;
  wire  _EVAL_1073;
  wire  _EVAL_1074;
  wire  _EVAL_1075;
  wire  _EVAL_1077;
  wire  _EVAL_1078;
  wire  _EVAL_1079;
  wire  _EVAL_1080;
  wire  _EVAL_1081;
  wire  _EVAL_1083;
  wire  _EVAL_1084;
  wire [31:0] _EVAL_1085;
  wire  _EVAL_1086;
  wire  _EVAL_1087;
  wire  _EVAL_1088;
  wire  _EVAL_1089;
  wire  _EVAL_1090;
  wire  _EVAL_1091;
  wire  _EVAL_1092;
  wire  _EVAL_1094;
  reg [1:0] _EVAL_1096;
  wire  _EVAL_1099;
  wire  _EVAL_1102;
  wire  _EVAL_1104;
  wire  _EVAL_1105;
  wire [2:0] _EVAL_1107;
  wire  _EVAL_1108;
  wire  _EVAL_1109;
  wire  _EVAL_1111;
  wire  _EVAL_1112;
  wire  _EVAL_1113;
  wire  _EVAL_1116;
  reg [7:0] _EVAL_1118;
  wire  _EVAL_1123;
  wire [23:0] _EVAL_1124;
  wire  _EVAL_1125;
  wire  _EVAL_1126;
  wire  _EVAL_1127;
  wire [7:0] _EVAL_1128;
  wire  _EVAL_1129;
  wire  _EVAL_1130;
  wire  _EVAL_1131;
  wire  _EVAL_1132;
  wire [11:0] _EVAL_1133;
  wire [15:0] _EVAL_1136;
  wire  _EVAL_1138;
  wire  _EVAL_1139;
  wire  _EVAL_1140;
  wire  _EVAL_1141;
  wire  _EVAL_1142;
  wire [31:0] _EVAL_1144;
  wire  _EVAL_1146;
  wire [31:0] _EVAL_1147;
  wire  _EVAL_1148;
  wire  _EVAL_1149;
  reg [7:0] _EVAL_1151;
  wire  _EVAL_1153;
  wire  _EVAL_1154;
  wire  _EVAL_1155;
  wire [7:0] _EVAL_1156;
  wire  _EVAL_1158;
  wire  _EVAL_1159;
  wire  _EVAL_1160;
  wire  _EVAL_1162;
  reg [7:0] _EVAL_1163;
  wire  _EVAL_1164;
  wire  _EVAL_1166;
  wire  _EVAL_1168;
  reg [7:0] _EVAL_1169;
  wire  _EVAL_1173;
  wire  _EVAL_1176;
  wire [31:0] _EVAL_1177;
  wire  _EVAL_1178;
  wire [7:0] _EVAL_1180;
  wire  _EVAL_1181;
  wire  _EVAL_1183;
  wire  _EVAL_1184;
  wire  _EVAL_1185;
  wire  _EVAL_1187;
  wire [31:0] _EVAL_1188;
  wire  _EVAL_1189;
  reg [7:0] _EVAL_1192;
  wire  _EVAL_1196;
  wire [28:0] _EVAL_1200;
  wire  _EVAL_1201;
  wire  _EVAL_1202;
  wire  _EVAL_1203;
  wire  _EVAL_1204;
  wire  _EVAL_1207;
  wire [31:0] _EVAL_1208;
  wire [31:0] _EVAL_1209;
  wire  _EVAL_1210;
  reg [7:0] _EVAL_1211;
  wire  _EVAL_1213;
  wire  _EVAL_1215;
  wire  _EVAL_1219;
  wire  _EVAL_1220;
  wire [1:0] _EVAL_1222;
  wire [31:0] _EVAL_1223;
  wire  _EVAL_1224;
  reg [7:0] _EVAL_1226;
  wire  _EVAL_1227;
  wire  _EVAL_1229;
  reg [7:0] _EVAL_1230;
  wire  _EVAL_1232;
  wire  _EVAL_1233;
  wire  _EVAL_1236;
  wire  _EVAL_1238;
  wire  _EVAL_1239;
  wire  _EVAL_1240;
  wire  _EVAL_1241;
  wire [2:0] _EVAL_1242;
  wire [15:0] _EVAL_1244;
  wire  _EVAL_1245;
  wire  _EVAL_1247;
  wire  _EVAL_1249;
  wire [31:0] _EVAL_1251;
  wire  _EVAL_1253;
  wire  _EVAL_1254;
  wire  _EVAL_1255;
  wire  _EVAL_1256;
  wire  _EVAL_1257;
  wire  _EVAL_1260;
  wire [31:0] _EVAL_1261;
  wire  _EVAL_1262;
  wire  _EVAL_1263;
  wire  _EVAL_1264;
  wire  _EVAL_1267;
  wire [127:0] _EVAL_1268;
  wire [21:0] _EVAL_1269;
  wire  _EVAL_1271;
  wire  _EVAL_1272;
  reg [7:0] _EVAL_1273;
  reg [7:0] _EVAL_1274;
  wire  _EVAL_1275;
  wire [31:0] _EVAL_1276;
  wire  _EVAL_1278;
  wire  _EVAL_1280;
  wire [31:0] _EVAL_1281;
  wire  _EVAL_1282;
  wire  _EVAL_1283;
  wire [31:0] _EVAL_1284;
  reg [2:0] _EVAL_1285;
  wire  _EVAL_1286;
  wire  _EVAL_1288;
  wire  _EVAL_1289;
  wire  _EVAL_1290;
  wire  _EVAL_1295;
  wire  _EVAL_1296;
  wire  _EVAL_1297;
  wire  _EVAL_1298;
  wire  _EVAL_1300;
  wire  _EVAL_1301;
  wire  _EVAL_1302;
  reg  _EVAL_1304;
  reg  _EVAL_1305;
  wire  _EVAL_1307;
  wire  _EVAL_1311;
  reg [7:0] _EVAL_1312;
  wire  _EVAL_1313;
  wire  _EVAL_1314;
  wire  _EVAL_1315;
  wire  _EVAL_1316;
  wire  _EVAL_1317;
  reg [7:0] _EVAL_1318;
  wire  _EVAL_1321;
  wire  _EVAL_1322;
  wire  _EVAL_1325;
  wire  _EVAL_1326;
  wire  _EVAL_1327;
  wire [31:0] _EVAL_1329;
  wire  _EVAL_1331;
  wire [511:0] _EVAL_1333;
  wire  _EVAL_1334;
  wire  _EVAL_1335;
  wire  _EVAL_1336;
  wire  _EVAL_1337;
  wire  _EVAL_1338;
  wire [4:0] _EVAL_1339;
  wire  _EVAL_1342;
  wire  _EVAL_1343;
  wire  _EVAL_1345;
  wire  _EVAL_1346;
  reg  _EVAL_1347;
  wire  _EVAL_1348;
  wire  _EVAL_1349;
  wire  _EVAL_1350;
  wire  _EVAL_1352;
  wire  _EVAL_1353;
  wire  _EVAL_1355;
  wire  _EVAL_1356;
  wire [31:0] _EVAL_1358;
  wire  _EVAL_1359;
  wire [7:0] _EVAL_1361;
  wire  _EVAL_1363;
  wire  _EVAL_1364;
  wire  _EVAL_1365;
  wire  _EVAL_1367;
  wire  _EVAL_1368;
  wire [31:0] _EVAL_1369;
  wire  _EVAL_1370;
  wire  _EVAL_1371;
  wire  _EVAL_1372;
  wire  _EVAL_1373;
  reg  _EVAL_1374;
  wire  _EVAL_1375;
  wire  _EVAL_1376;
  wire [7:0] _EVAL_1378;
  wire  _EVAL_1379;
  wire  _EVAL_1380;
  wire  _EVAL_1381;
  reg [7:0] _EVAL_1384;
  wire  _EVAL_1386;
  wire  _EVAL_1388;
  wire  _EVAL_1389;
  wire  sb2tlOpt__EVAL;
  wire  sb2tlOpt__EVAL_0;
  wire  sb2tlOpt__EVAL_1;
  wire  sb2tlOpt__EVAL_2;
  wire [31:0] sb2tlOpt__EVAL_3;
  wire  sb2tlOpt__EVAL_4;
  wire  sb2tlOpt__EVAL_5;
  wire [7:0] sb2tlOpt__EVAL_6;
  wire  sb2tlOpt__EVAL_7;
  wire [7:0] sb2tlOpt__EVAL_8;
  wire  sb2tlOpt__EVAL_9;
  wire [3:0] sb2tlOpt__EVAL_10;
  wire  sb2tlOpt__EVAL_11;
  wire  sb2tlOpt__EVAL_12;
  wire  sb2tlOpt__EVAL_13;
  wire  sb2tlOpt__EVAL_14;
  wire [2:0] sb2tlOpt__EVAL_15;
  wire [2:0] sb2tlOpt__EVAL_16;
  wire [127:0] sb2tlOpt__EVAL_17;
  wire [2:0] sb2tlOpt__EVAL_18;
  wire  sb2tlOpt__EVAL_19;
  wire  sb2tlOpt__EVAL_20;
  wire  sb2tlOpt__EVAL_21;
  wire  sb2tlOpt__EVAL_22;
  wire  sb2tlOpt__EVAL_23;
  wire  sb2tlOpt__EVAL_24;
  wire [127:0] sb2tlOpt__EVAL_25;
  wire [7:0] sb2tlOpt__EVAL_26;
  wire  sb2tlOpt__EVAL_27;
  wire  _EVAL_1390;
  wire  _EVAL_1392;
  wire  _EVAL_1394;
  wire  _EVAL_1396;
  wire [31:0] _EVAL_1399;
  wire  _EVAL_1400;
  wire  _EVAL_1403;
  wire [31:0] _EVAL_1406;
  wire  _EVAL_1408;
  wire  _EVAL_1409;
  wire  _EVAL_1410;
  wire  _EVAL_1411;
  wire  _EVAL_1412;
  wire [31:0] _EVAL_1414;
  wire  _EVAL_1415;
  reg [15:0] _EVAL_1416;
  wire  _EVAL_1418;
  wire  _EVAL_1419;
  wire [7:0] _EVAL_1420;
  wire  _EVAL_1421;
  wire  _EVAL_1422;
  wire  _EVAL_1423;
  wire  _EVAL_1425;
  wire  _EVAL_1428;
  wire  _EVAL_1431;
  wire  _EVAL_1432;
  wire  _EVAL_1435;
  reg [7:0] _EVAL_1438;
  wire  _EVAL_1441;
  wire  _EVAL_1442;
  wire  _EVAL_1443;
  wire  _EVAL_1445;
  wire  _EVAL_1446;
  wire  _EVAL_1448;
  wire [2:0] _EVAL_1450;
  wire  _EVAL_1451;
  wire  _EVAL_1452;
  reg [7:0] _EVAL_1454;
  wire  _EVAL_1455;
  wire  _EVAL_1458;
  wire  _EVAL_1459;
  wire  _EVAL_1460;
  wire  _EVAL_1461;
  wire  _EVAL_1463;
  wire  _EVAL_1466;
  wire  _EVAL_1468;
  wire  _EVAL_1471;
  wire  _EVAL_1472;
  wire  _EVAL_1473;
  wire  _EVAL_1474;
  wire  _EVAL_1475;
  wire  _EVAL_1477;
  wire  _EVAL_1480;
  reg [7:0] _EVAL_1482;
  reg [7:0] _EVAL_1483;
  wire  _EVAL_1485;
  wire  _EVAL_1486;
  wire  _EVAL_1488;
  wire  _EVAL_1489;
  wire  _EVAL_1490;
  wire  _EVAL_1498;
  wire [31:0] _EVAL_1501;
  wire [31:0] _EVAL_1502;
  wire  _EVAL_1503;
  wire  _EVAL_1504;
  wire  _EVAL_1505;
  wire  _EVAL_1507;
  wire  _EVAL_1513;
  wire  _EVAL_1515;
  wire  _EVAL_1516;
  wire  _EVAL_1518;
  wire  _EVAL_1519;
  reg [7:0] _EVAL_1520;
  wire  _EVAL_1522;
  wire  _EVAL_1524;
  wire  _EVAL_1527;
  wire  _EVAL_1529;
  wire  _EVAL_1530;
  wire  _EVAL_1532;
  wire  _EVAL_1533;
  wire  _EVAL_1534;
  wire  _EVAL_1537;
  wire  _EVAL_1539;
  reg  _EVAL_1541;
  wire  _EVAL_1542;
  wire [1:0] _EVAL_1543;
  wire [31:0] _EVAL_1544;
  wire  _EVAL_1545;
  wire  _EVAL_1546;
  wire  _EVAL_1549;
  wire  _EVAL_1552;
  wire  _EVAL_1553;
  wire  _EVAL_1556;
  wire  _EVAL_1557;
  wire  _EVAL_1558;
  wire  _EVAL_1559;
  wire  _EVAL_1561;
  wire [1:0] _EVAL_1563;
  wire [6:0] _EVAL_1565;
  wire  _EVAL_1566;
  wire [22:0] _EVAL_1567;
  wire  _EVAL_1568;
  wire  _EVAL_1571;
  wire  _EVAL_1572;
  wire  _EVAL_1574;
  wire  _EVAL_1575;
  wire  _EVAL_1577;
  wire  _EVAL_1578;
  wire [31:0] _EVAL_1579;
  wire  _EVAL_1580;
  wire [3:0] _EVAL_1581;
  wire  _EVAL_1582;
  wire  _EVAL_1583;
  wire  _EVAL_1586;
  wire  _EVAL_1587;
  wire  _EVAL_1588;
  wire [2:0] _EVAL_1590;
  wire  _EVAL_1591;
  wire  _EVAL_1592;
  wire  _EVAL_1593;
  wire  _EVAL_1596;
  wire  _EVAL_1599;
  wire  _EVAL_1600;
  wire  _EVAL_1601;
  wire  _EVAL_1603;
  wire  _EVAL_1604;
  wire  _EVAL_1605;
  wire  _EVAL_1606;
  wire  _EVAL_1607;
  wire  _EVAL_1610;
  wire  _EVAL_1612;
  wire  _EVAL_1613;
  wire  _EVAL_1614;
  wire  _EVAL_1615;
  reg [7:0] _EVAL_1616;
  wire  _EVAL_1618;
  wire  _EVAL_1620;
  wire  _EVAL_1623;
  wire  _EVAL_1627;
  wire  _EVAL_1629;
  wire  _EVAL_1632;
  wire  _EVAL_1633;
  wire  _EVAL_1634;
  wire  _EVAL_1635;
  wire [7:0] _EVAL_1636;
  wire  _EVAL_1637;
  wire  _EVAL_1638;
  wire  _EVAL_1640;
  wire  _EVAL_1641;
  wire  _EVAL_1642;
  wire [31:0] _EVAL_1643;
  wire [31:0] _EVAL_1644;
  wire  _EVAL_1646;
  wire  _EVAL_1648;
  wire  _EVAL_1650;
  wire  _EVAL_1652;
  wire  _EVAL_1653;
  wire [31:0] _EVAL_1657;
  wire  _EVAL_1658;
  wire  _EVAL_1659;
  wire  _EVAL_1660;
  wire  _EVAL_1663;
  reg [7:0] _EVAL_1664;
  wire  _EVAL_1666;
  wire  _EVAL_1667;
  wire  _EVAL_1669;
  wire [7:0] _EVAL_1672;
  wire [31:0] _EVAL_1675;
  wire  _EVAL_1677;
  wire  _EVAL_1678;
  wire [31:0] _EVAL_1679;
  wire  _EVAL_1681;
  wire  _EVAL_1682;
  wire  _EVAL_1683;
  wire  _EVAL_1685;
  wire [31:0] _EVAL_1687;
  wire  _EVAL_1688;
  wire [31:0] _EVAL_1689;
  wire  _EVAL_1693;
  wire [31:0] _EVAL_1694;
  wire  _EVAL_1697;
  wire  _EVAL_1698;
  wire [128:0] _EVAL_1702;
  wire  _EVAL_1703;
  wire [2:0] _EVAL_1704;
  wire [31:0] _EVAL_1705;
  wire  _EVAL_1706;
  wire  _EVAL_1707;
  wire  _EVAL_1710;
  wire [31:0] _EVAL_1711;
  wire [15:0] _EVAL_1712;
  wire  _EVAL_1713;
  wire  _EVAL_1714;
  wire [7:0] _EVAL_1715;
  wire [7:0] _EVAL_1716;
  wire  _EVAL_1717;
  wire  _EVAL_1718;
  wire  _EVAL_1719;
  wire  _EVAL_1720;
  wire  _EVAL_1721;
  reg [7:0] _EVAL_1722;
  reg [7:0] _EVAL_1723;
  wire  _EVAL_1724;
  wire  _EVAL_1726;
  wire  _EVAL_1728;
  wire  _EVAL_1729;
  wire  _EVAL_1730;
  wire  _EVAL_1731;
  wire  _EVAL_1732;
  wire  _EVAL_1735;
  wire [1:0] _EVAL_1737;
  wire [31:0] _EVAL_1738;
  wire [31:0] _EVAL_1740;
  wire  _EVAL_1742;
  wire  _EVAL_1743;
  wire  _EVAL_1744;
  wire  _EVAL_1745;
  wire [31:0] _EVAL_1749;
  wire [16:0] _EVAL_1751;
  wire  _EVAL_1752;
  wire  _EVAL_1756;
  wire  _EVAL_1757;
  wire  _EVAL_1758;
  wire  _EVAL_1762;
  wire  _EVAL_1763;
  wire  _EVAL_1765;
  wire  _EVAL_1767;
  wire [31:0] _EVAL_1768;
  wire  _EVAL_1769;
  wire  _EVAL_1770;
  wire  _EVAL_1773;
  wire  _EVAL_1774;
  wire [15:0] _EVAL_1775;
  wire  _EVAL_1778;
  wire  _EVAL_1779;
  reg [7:0] _EVAL_1781;
  wire  _EVAL_1783;
  wire  _EVAL_1784;
  wire  _EVAL_1785;
  wire  _EVAL_1790;
  wire  _EVAL_1791;
  wire  _EVAL_1792;
  wire [1:0] _EVAL_1793;
  wire  _EVAL_1794;
  wire  _EVAL_1795;
  wire  _EVAL_1796;
  wire [31:0] _EVAL_1798;
  wire  _EVAL_1801;
  wire  _EVAL_1803;
  wire  _EVAL_1804;
  wire  _EVAL_1805;
  wire  _EVAL_1807;
  wire  _EVAL_1808;
  wire  _EVAL_1811;
  wire  _EVAL_1812;
  wire  _EVAL_1813;
  wire [31:0] _EVAL_1815;
  reg [7:0] _EVAL_1816;
  wire  _EVAL_1817;
  wire  _EVAL_1819;
  wire  _EVAL_1823;
  wire  _EVAL_1824;
  wire  _EVAL_1826;
  reg [7:0] _EVAL_1828;
  wire  _EVAL_1833;
  wire  _EVAL_1834;
  wire  _EVAL_1835;
  wire  _EVAL_1837;
  wire  _EVAL_1839;
  wire  _EVAL_1841;
  wire  _EVAL_1843;
  reg [7:0] _EVAL_1844;
  wire  _EVAL_1845;
  wire  _EVAL_1846;
  wire [31:0] _EVAL_1847;
  wire  _EVAL_1848;
  wire [31:0] _EVAL_1849;
  wire  _EVAL_1850;
  wire  _EVAL_1852;
  reg [7:0] _EVAL_1853;
  wire  _EVAL_1857;
  wire  _EVAL_1858;
  wire  _EVAL_1859;
  wire  _EVAL_1861;
  wire [31:0] _EVAL_1863;
  wire  _EVAL_1864;
  wire  _EVAL_1865;
  wire  _EVAL_1866;
  wire  _EVAL_1867;
  wire  _EVAL_1868;
  wire  _EVAL_1869;
  wire  _EVAL_1875;
  wire  _EVAL_1876;
  wire [7:0] _EVAL_1877;
  wire  _EVAL_1880;
  wire  _EVAL_1881;
  reg [7:0] _EVAL_1882;
  wire  _EVAL_1884;
  wire  _EVAL_1885;
  reg  _EVAL_1886;
  wire  _EVAL_1887;
  wire  _EVAL_1888;
  wire  _EVAL_1889;
  wire  _EVAL_1894;
  wire [31:0] _EVAL_1895;
  wire  _EVAL_1897;
  wire  _EVAL_1898;
  wire  _EVAL_1900;
  wire  _EVAL_1901;
  wire  _EVAL_1903;
  reg  _EVAL_1904;
  reg [7:0] _EVAL_1905;
  wire  _EVAL_1906;
  reg [7:0] _EVAL_1907;
  wire  _EVAL_1908;
  wire  _EVAL_1909;
  wire  _EVAL_1910;
  wire  _EVAL_1914;
  wire  _EVAL_1915;
  wire  _EVAL_1917;
  reg [7:0] _EVAL_1918;
  wire  _EVAL_1920;
  wire  _EVAL_1921;
  reg [7:0] _EVAL_1922;
  wire  _EVAL_1923;
  wire  _EVAL_1925;
  wire  _EVAL_1927;
  wire  _EVAL_1928;
  wire  _EVAL_1929;
  wire  _EVAL_1931;
  wire  _EVAL_1932;
  wire  _EVAL_1933;
  wire [31:0] _EVAL_1934;
  wire  _EVAL_1936;
  wire  _EVAL_1940;
  wire  _EVAL_1941;
  reg [31:0] _EVAL_1943;
  wire  _EVAL_1944;
  wire  _EVAL_1945;
  wire  _EVAL_1946;
  wire  _EVAL_1948;
  wire  _EVAL_1950;
  wire  _EVAL_1953;
  wire  _EVAL_1956;
  wire  _EVAL_1957;
  wire  _EVAL_1958;
  wire  _EVAL_1959;
  wire [31:0] _EVAL_1961;
  wire  _EVAL_1962;
  wire  _EVAL_1964;
  wire  _EVAL_1965;
  wire [31:0] _EVAL_1966;
  wire  _EVAL_1969;
  reg [7:0] _EVAL_1970;
  wire  _EVAL_1971;
  wire  _EVAL_1972;
  wire [31:0] _EVAL_1973;
  wire  _EVAL_1974;
  wire  _EVAL_1975;
  wire  _EVAL_1976;
  wire  _EVAL_1977;
  wire [5:0] _EVAL_1978;
  wire  _EVAL_1979;
  wire [7:0] _EVAL_1980;
  wire  _EVAL_1982;
  wire  _EVAL_1984;
  wire  _EVAL_1985;
  wire  _EVAL_1986;
  wire  _EVAL_1987;
  wire  _EVAL_1988;
  reg [23:0] _EVAL_1989;
  wire  _EVAL_1991;
  wire  _EVAL_1992;
  wire  _EVAL_1994;
  wire  _EVAL_1996;
  wire  _EVAL_1997;
  wire [31:0] _EVAL_1998;
  wire  _EVAL_2000;
  wire  _EVAL_2001;
  wire [31:0] _EVAL_2002;
  wire  _EVAL_2003;
  wire  _EVAL_2008;
  wire  _EVAL_2009;
  wire  _EVAL_2011;
  wire  _EVAL_2014;
  wire  _EVAL_2015;
  wire  _EVAL_2017;
  wire  _EVAL_2018;
  wire [31:0] _EVAL_2025;
  wire  _EVAL_2027;
  wire  _EVAL_2028;
  wire [7:0] _EVAL_2030;
  wire  _EVAL_2031;
  reg [7:0] _EVAL_2032;
  wire  _EVAL_2033;
  wire  _EVAL_2034;
  wire  _EVAL_2035;
  wire  _EVAL_2036;
  wire  _EVAL_2037;
  wire  _EVAL_2039;
  wire  _EVAL_2041;
  wire  _EVAL_2042;
  wire  _EVAL_2043;
  wire  _EVAL_2044;
  wire  _EVAL_2045;
  wire  _EVAL_2046;
  wire  _EVAL_2047;
  wire  _EVAL_2049;
  wire  _EVAL_2050;
  wire  _EVAL_2051;
  wire  _EVAL_2052;
  _EVAL_176 hartIsInResetSync_0_debug_hartReset_0 (
    ._EVAL(hartIsInResetSync_0_debug_hartReset_0__EVAL),
    ._EVAL_0(hartIsInResetSync_0_debug_hartReset_0__EVAL_0),
    ._EVAL_1(hartIsInResetSync_0_debug_hartReset_0__EVAL_1),
    ._EVAL_2(hartIsInResetSync_0_debug_hartReset_0__EVAL_2)
  );
  _EVAL_173 sb2tlOpt (
    ._EVAL(sb2tlOpt__EVAL),
    ._EVAL_0(sb2tlOpt__EVAL_0),
    ._EVAL_1(sb2tlOpt__EVAL_1),
    ._EVAL_2(sb2tlOpt__EVAL_2),
    ._EVAL_3(sb2tlOpt__EVAL_3),
    ._EVAL_4(sb2tlOpt__EVAL_4),
    ._EVAL_5(sb2tlOpt__EVAL_5),
    ._EVAL_6(sb2tlOpt__EVAL_6),
    ._EVAL_7(sb2tlOpt__EVAL_7),
    ._EVAL_8(sb2tlOpt__EVAL_8),
    ._EVAL_9(sb2tlOpt__EVAL_9),
    ._EVAL_10(sb2tlOpt__EVAL_10),
    ._EVAL_11(sb2tlOpt__EVAL_11),
    ._EVAL_12(sb2tlOpt__EVAL_12),
    ._EVAL_13(sb2tlOpt__EVAL_13),
    ._EVAL_14(sb2tlOpt__EVAL_14),
    ._EVAL_15(sb2tlOpt__EVAL_15),
    ._EVAL_16(sb2tlOpt__EVAL_16),
    ._EVAL_17(sb2tlOpt__EVAL_17),
    ._EVAL_18(sb2tlOpt__EVAL_18),
    ._EVAL_19(sb2tlOpt__EVAL_19),
    ._EVAL_20(sb2tlOpt__EVAL_20),
    ._EVAL_21(sb2tlOpt__EVAL_21),
    ._EVAL_22(sb2tlOpt__EVAL_22),
    ._EVAL_23(sb2tlOpt__EVAL_23),
    ._EVAL_24(sb2tlOpt__EVAL_24),
    ._EVAL_25(sb2tlOpt__EVAL_25),
    ._EVAL_26(sb2tlOpt__EVAL_26),
    ._EVAL_27(sb2tlOpt__EVAL_27)
  );
  assign _EVAL_561 = _EVAL_391 & _EVAL_116;
  assign _EVAL_1593 = _EVAL_204 ? _EVAL_959 : _EVAL_280;
  assign _EVAL_537 = _EVAL_883 | _EVAL_122;
  assign _EVAL_2014 = _EVAL_1730 & _EVAL_743;
  assign _EVAL_910 = _EVAL_427 & _EVAL_1603;
  assign _EVAL_259 = {{14'd0}, _EVAL_1563};
  assign _EVAL_548 = _EVAL_1140 & _EVAL_150;
  assign _EVAL_407 = _EVAL_311 & _EVAL_1522;
  assign _EVAL_666 = _EVAL_90 & _EVAL_1074;
  assign _EVAL_1908 = _EVAL_1841 & _EVAL_1024;
  assign _EVAL_144 = _EVAL_1719 | _EVAL_875;
  assign _EVAL_755 = _EVAL_1140 & _EVAL_923;
  assign _EVAL_668 = _EVAL_2000 & _EVAL_566;
  assign _EVAL_1991 = _EVAL_1342 | _EVAL_1898;
  assign _EVAL_1255 = _EVAL_626 & _EVAL_223;
  assign _EVAL_1682 = _EVAL_650 | _EVAL_942;
  assign sb2tlOpt__EVAL_15 = _EVAL_1285;
  assign _EVAL_1102 = 9'h108 == _EVAL_351;
  assign _EVAL_1572 = _EVAL_1176 & _EVAL_911;
  assign _EVAL_105 = _EVAL_589 | _EVAL_362;
  assign _EVAL_865 = ~_EVAL_385;
  assign _EVAL_640 = _EVAL_1177[7:0];
  assign _EVAL_604 = _EVAL_39[14:12];
  assign _EVAL_1166 = _EVAL_882 | _EVAL_83;
  assign _EVAL_650 = _EVAL_222 | _EVAL_513;
  assign _EVAL_310 = _EVAL_345 & _EVAL_177;
  assign _EVAL_354 = _EVAL_305 ? _EVAL_1086 : _EVAL_845;
  assign _EVAL_611 = _EVAL_348 | _EVAL_508;
  assign _EVAL_1773 = &_EVAL_554;
  assign _EVAL_1707 = _EVAL_276 & _EVAL_223;
  assign _EVAL_921 = _EVAL_1925 & _EVAL_1824;
  assign _EVAL_1164 = _EVAL_586[36];
  assign _EVAL_937 = _EVAL_555 ? _EVAL_347 : _EVAL_1643;
  assign _EVAL_1977 = _EVAL_670 & _EVAL_1001;
  assign _EVAL_297 = _EVAL_1635 | _EVAL_239;
  assign _EVAL_217 = _EVAL_1724 ? _EVAL_959 : _EVAL_148;
  assign _EVAL_1502 = {_EVAL_1128,_EVAL_1980,_EVAL_1378,_EVAL_1672};
  assign _EVAL_1028 = _EVAL_286 & _EVAL_223;
  assign _EVAL_613 = _EVAL_345 & _EVAL_1074;
  assign _EVAL_177 = &_EVAL_765;
  assign _EVAL_198 = _EVAL_707 | _EVAL_340;
  assign _EVAL_866 = _EVAL_287 & _EVAL_1928;
  assign _EVAL_131 = _EVAL_1607 | _EVAL_727;
  assign _EVAL_1104 = _EVAL_1333[64];
  assign _EVAL_883 = _EVAL_1372 & _EVAL_223;
  assign _EVAL_1688 = _EVAL_1737 != 2'h0;
  assign _EVAL_513 = _EVAL_1985 | _EVAL_216;
  assign _EVAL_844 = _EVAL_556 & _EVAL_1846;
  assign _EVAL_1477 = 9'h40 == _EVAL_351;
  assign _EVAL_1089 = _EVAL_1348 | _EVAL_109;
  assign _EVAL_928 = sb2tlOpt__EVAL_12 & _EVAL_1455;
  assign _EVAL_351 = {_EVAL_1591,_EVAL_1728,_EVAL_411,_EVAL_1969,_EVAL_574,_EVAL_162,_EVAL_671,_EVAL_776,_EVAL_857};
  assign _EVAL_1743 = _EVAL_568 & _EVAL_1007;
  assign _EVAL_1803 = 9'h113 == _EVAL_351;
  assign _EVAL_550 = _EVAL_680 & _EVAL_1796;
  assign _EVAL_685 = _EVAL_1062 & _EVAL_1001;
  assign _EVAL_905 = {17'h7000,_EVAL_1590,_EVAL_1339,7'h3};
  assign _EVAL_494 = |_EVAL_736;
  assign _EVAL_1296 = _EVAL_1166 | _EVAL_198;
  assign _EVAL_1650 = _EVAL_1386 | _EVAL_124;
  assign _EVAL_638 = _EVAL_724 & _EVAL_854;
  assign _EVAL_215 = _EVAL_1763 & _EVAL_1603;
  assign _EVAL_1843 = _EVAL_1403 & _EVAL_1086;
  assign _EVAL_361 = 6'h38 == _EVAL_1978;
  assign _EVAL_1140 = _EVAL_1183 & _EVAL_739;
  assign _EVAL_923 = _EVAL_586[37];
  assign hartIsInResetSync_0_debug_hartReset_0__EVAL_1 = _EVAL_30;
  assign _EVAL_1375 = _EVAL_1693 & _EVAL_1335;
  assign _EVAL_1724 = 9'hd6 == _EVAL_351;
  assign _EVAL_1185 = _EVAL_521 & _EVAL_1928;
  assign _EVAL_862 = {3'h1,_EVAL_1200};
  assign _EVAL_403 = {_EVAL_988,_EVAL_1169,_EVAL_1918,_EVAL_606};
  assign _EVAL_1149 = _EVAL_729 & _EVAL_2045;
  assign _EVAL_831 = _EVAL_767 & _EVAL_116;
  assign _EVAL_1720 = _EVAL_328 ? _EVAL_959 : _EVAL_1213;
  assign _EVAL_1055 = _EVAL_341 & _EVAL_393;
  assign _EVAL_586 = 64'h1 << _EVAL_1978;
  assign _EVAL_653 = 6'h2c == _EVAL_1978;
  assign _EVAL_761 = _EVAL_1334 ? 32'h30000067 : _EVAL_828;
  assign _EVAL_971 = _EVAL_936 ? _EVAL_121 : _EVAL_791;
  assign _EVAL_1612 = 9'hdf == _EVAL_351;
  assign _EVAL_1229 = _EVAL_228 & _EVAL_1824;
  assign _EVAL_219 = _EVAL_690 & _EVAL_854;
  assign _EVAL_438 = _EVAL_391 & _EVAL_1458;
  assign _EVAL_317 = _EVAL_1333[214];
  assign sb2tlOpt__EVAL_17 = sb2tlOpt__EVAL_27 ? _EVAL_242 : _EVAL_140;
  assign _EVAL_891 = _EVAL_1352 & _EVAL_1086;
  assign _EVAL_1567 = {1'h0,_EVAL_1269};
  assign _EVAL_1600 = _EVAL_1557 | _EVAL_1313;
  assign _EVAL_369 = _EVAL_1333[223];
  assign _EVAL_1244 = {{7'd0}, _EVAL_87};
  assign _EVAL_515 = _EVAL_1337 ? _EVAL_1086 : _EVAL_758;
  assign _EVAL_473 = _EVAL_225 | _EVAL_563;
  assign _EVAL_574 = _EVAL_939[4];
  assign _EVAL_776 = _EVAL_939[1];
  assign _EVAL_1183 = _EVAL_17 & _EVAL_36;
  assign _EVAL_718 = 6'h20 == _EVAL_1978;
  assign _EVAL_265 = {_EVAL_1416,_EVAL_259};
  assign _EVAL_180 = _EVAL_305 ? _EVAL_285 : _EVAL_281;
  assign _EVAL_886 = _EVAL_1338 & _EVAL_1603;
  assign _EVAL_817 = _EVAL_1565[4];
  assign _EVAL_1349 = 9'h104 == _EVAL_351;
  assign _EVAL_1672 = _EVAL_933 ? 8'hff : 8'h0;
  assign _EVAL_117 = ~_EVAL_1460;
  assign _EVAL_1897 = _EVAL_1561 | _EVAL_772;
  assign _EVAL_1223 = _EVAL_1146 ? _EVAL_476 : _EVAL_1687;
  assign _EVAL_430 = 8'h1 << _EVAL_1285;
  assign _EVAL_1313 = _EVAL_484 & _EVAL_1127;
  assign _EVAL_1557 = _EVAL_753 & _EVAL_675;
  assign _EVAL_1580 = _EVAL_827 | _EVAL_1123;
  assign _EVAL_976 = _EVAL_1843 & _EVAL_494;
  assign hartIsInResetSync_0_debug_hartReset_0__EVAL_0 = _EVAL_14;
  assign _EVAL_559 = _EVAL_1485 | _EVAL_577;
  assign _EVAL_1571 = _EVAL_1901 | _EVAL_74;
  assign _EVAL_474 = 9'h10c == _EVAL_351;
  assign _EVAL_1767 = _EVAL_1590 == 3'h3;
  assign _EVAL_1245 = _EVAL_712 & _EVAL_1522;
  assign _EVAL_115 = _EVAL_210 | _EVAL_1982;
  assign _EVAL_1002 = _EVAL_1502[20];
  assign _EVAL_1026 = _EVAL_276 & _EVAL_1971;
  assign _EVAL_906 = _EVAL_564 ? _EVAL_959 : _EVAL_258;
  assign _EVAL_1201 = _EVAL_28 & _EVAL_44;
  assign _EVAL_530 = _EVAL_84 & _EVAL_1603;
  assign _EVAL_1693 = _EVAL_1295 & _EVAL_1086;
  assign _EVAL_1159 = _EVAL_423 & _EVAL_494;
  assign _EVAL_1086 = _EVAL_200 == 7'h0;
  assign _EVAL_1373 = _EVAL_1263 ? _EVAL_959 : _EVAL_1720;
  assign _EVAL_1423 = _EVAL_1043 | _EVAL_227;
  assign _EVAL_676 = _EVAL_1979 | _EVAL_1784;
  assign _EVAL_373 = _EVAL_1848 ? 1'h0 : _EVAL_272;
  assign _EVAL_1941 = _EVAL_1757 & _EVAL_1603;
  assign _EVAL_1052 = 6'h28 == _EVAL_1978;
  assign _EVAL_237 = _EVAL_641 & _EVAL_959;
  assign _EVAL_631 = _EVAL_1565[1];
  assign _EVAL_1408 = _EVAL_842 & _EVAL_1603;
  assign _EVAL_811 = _EVAL_712 & _EVAL_1001;
  assign _EVAL_1934 = _EVAL_1953 ? 32'h0 : _EVAL_231;
  assign _EVAL_1280 = _EVAL_114 & _EVAL_494;
  assign _EVAL_1711 = _EVAL_417 ? _EVAL_1943 : _EVAL_954;
  assign _EVAL_1763 = _EVAL_1703 & _EVAL_116;
  assign _EVAL_867 = _EVAL_375 & _EVAL_959;
  assign _EVAL_1316 = _EVAL_1333[65];
  assign _EVAL_326 = _EVAL_1915 & _EVAL_2027;
  assign _EVAL_1083 = _EVAL_1062 & _EVAL_1522;
  assign _EVAL_1369 = _EVAL_718 ? _EVAL_999 : _EVAL_1085;
  assign _EVAL_1422 = _EVAL_1502[0];
  assign _EVAL_1184 = _EVAL_1471 & _EVAL_1472;
  assign _EVAL_228 = _EVAL_1132 & _EVAL_1012;
  assign _EVAL_651 = _EVAL_195 ? 8'hff : 8'h0;
  assign _EVAL_778 = _EVAL_586[23];
  assign _EVAL_1966 = _EVAL_1142 ? 32'h440006f : _EVAL_445;
  assign _EVAL_74 = _EVAL_1552 | _EVAL_1290;
  assign _EVAL_1527 = _EVAL_168 & _EVAL_1928;
  assign _EVAL_1389 = _EVAL_360 ? _EVAL_959 : _EVAL_733;
  assign _EVAL_1945 = _EVAL_1974 ? _EVAL_959 : _EVAL_1288;
  assign _EVAL_1667 = _EVAL_76 & _EVAL_1370;
  assign _EVAL_1714 = _EVAL_168 & _EVAL_177;
  assign _EVAL_1586 = _EVAL_1381 & _EVAL_1603;
  assign _EVAL_894 = 9'h105 == _EVAL_351;
  assign _EVAL_1365 = _EVAL_1785 | _EVAL_821;
  assign _EVAL_1903 = _EVAL_1486 & _EVAL_1078;
  assign _EVAL_290 = _EVAL_617 & _EVAL_1086;
  assign _EVAL_1153 = _EVAL_1325 & _EVAL_1045;
  assign _EVAL_1898 = _EVAL_1380 & _EVAL_1001;
  assign _EVAL_946 = _EVAL_126 | _EVAL_654;
  assign _EVAL_337 = _EVAL_972 & _EVAL_177;
  assign _EVAL_797 = _EVAL_1770 & _EVAL_959;
  assign _EVAL_429 = _EVAL_1416[6];
  assign _EVAL_383 = _EVAL_1177[31:24];
  assign _EVAL_1314 = 6'h17 == _EVAL_1978;
  assign _EVAL_1168 = 9'h10a == _EVAL_351;
  assign _EVAL_1971 = &_EVAL_68;
  assign _EVAL_1254 = _EVAL_84 | _EVAL_1958;
  assign _EVAL_455 = _EVAL_1549 | _EVAL_309;
  assign _EVAL_897 = _EVAL_400 & _EVAL_924;
  assign _EVAL_299 = _EVAL_632 ? _EVAL_121 : _EVAL_174;
  assign _EVAL_72 = _EVAL_709 & _EVAL_1773;
  assign _EVAL_996 = _EVAL_336 & _EVAL_1086;
  assign _EVAL_107 = _EVAL_182 & _EVAL_1928;
  assign _EVAL_782 = {{31'd0}, _EVAL_566};
  assign _EVAL_22 = sb2tlOpt__EVAL_22;
  assign _EVAL_291 = _EVAL_1013 | _EVAL_1229;
  assign _EVAL_821 = _EVAL_1451 & _EVAL_1012;
  assign _EVAL_390 = _EVAL_1168 ? 32'h147413 : _EVAL_441;
  assign _EVAL_1090 = _EVAL_526 | _EVAL_1300;
  assign _EVAL_1213 = _EVAL_1953 ? _EVAL_959 : _EVAL_1945;
  assign _EVAL_1073 = _EVAL_1416[7];
  assign _EVAL_57 = sb2tlOpt__EVAL_27 & _EVAL_1839;
  assign _EVAL_1486 = _EVAL_831 | _EVAL_607;
  assign _EVAL_1380 = _EVAL_453 & _EVAL_1086;
  assign _EVAL_467 = _EVAL_1127 ? 1'h0 : _EVAL_332;
  assign _EVAL_104 = _EVAL_400 & _EVAL_1316;
  assign _EVAL_1030 = _EVAL_1610 | _EVAL_660;
  assign _EVAL_97 = _EVAL_1176 | _EVAL_108;
  assign _EVAL_1480 = _EVAL_1669 | _EVAL_1904;
  assign _EVAL_1623 = _EVAL_1346 & _EVAL_1353;
  assign _EVAL_1652 = _EVAL_1416[1];
  assign _EVAL_975 = _EVAL_1428 | _EVAL_447;
  assign _EVAL_366 = _EVAL_1285 == 3'h2;
  assign _EVAL_1635 = _EVAL_291 | _EVAL_1461;
  assign _EVAL_623 = _EVAL_920 & _EVAL_177;
  assign _EVAL_1932 = _EVAL_1342 & _EVAL_1603;
  assign _EVAL_1658 = _EVAL_867 & _EVAL_177;
  assign _EVAL_658 = _EVAL_586[56];
  assign _EVAL_933 = _EVAL_43[0];
  assign _EVAL_1794 = _EVAL_413 & _EVAL_1928;
  assign _EVAL_1793 = _EVAL_332 ? 2'h0 : 2'h2;
  assign _EVAL_2003 = _EVAL_450 & _EVAL_223;
  assign _EVAL_466 = 6'h25 == _EVAL_1978;
  assign _EVAL_1563 = {1'h0,_EVAL_1253};
  assign _EVAL_1317 = _EVAL_891 & _EVAL_1971;
  assign _EVAL_1666 = &_EVAL_737;
  assign _EVAL_322 = _EVAL_438 & _EVAL_1603;
  assign _EVAL_1138 = _EVAL_1333[215];
  assign _EVAL_1504 = 9'h10f == _EVAL_351;
  assign sb2tlOpt__EVAL_14 = _EVAL_4;
  assign _EVAL_272 = _EVAL_1355 | _EVAL_647;
  assign _EVAL_2043 = _EVAL_1515 & _EVAL_177;
  assign _EVAL_307 = _EVAL_678[2:0];
  assign _EVAL_1566 = _EVAL_888 & _EVAL_1603;
  assign _EVAL_736 = _EVAL_1502[7:0];
  assign _EVAL_1132 = _EVAL_665 & _EVAL_1086;
  assign _EVAL_654 = _EVAL_888 | _EVAL_1744;
  assign _EVAL_727 = _EVAL_510 & _EVAL_958;
  assign _EVAL_688 = _EVAL_689 ? _EVAL_2018 : _EVAL_515;
  assign _EVAL_1415 = _EVAL_273 & _EVAL_1086;
  assign _EVAL_982 = _EVAL_1653 ? _EVAL_1086 : _EVAL_1894;
  assign _EVAL_973 = _EVAL_1380 & _EVAL_1522;
  assign _EVAL_1173 = _EVAL_1853 == 8'h0;
  assign _EVAL_723 = _EVAL_1502[10:8];
  assign _EVAL_1534 = _EVAL_767 & _EVAL_223;
  assign _EVAL_1141 = 9'hd8 == _EVAL_351;
  assign _EVAL_1321 = _EVAL_1333[218];
  assign _EVAL_2011 = _EVAL_2003 & _EVAL_1603;
  assign _EVAL_400 = _EVAL_904 & _EVAL_1518;
  assign _EVAL_1678 = _EVAL_1765 | _EVAL_1903;
  assign _EVAL_1592 = |_EVAL_782;
  assign _EVAL_1394 = _EVAL_586[42];
  assign _EVAL_437 = _EVAL_1046 | _EVAL_563;
  assign _EVAL_182 = _EVAL_1301 & _EVAL_959;
  assign _EVAL_2000 = _EVAL_1541 | _EVAL_870;
  assign _EVAL_1247 = _EVAL_797 & _EVAL_1773;
  assign _EVAL_1973 = _EVAL_1337 ? _EVAL_1740 : _EVAL_1849;
  assign _EVAL_1411 = _EVAL_920 & _EVAL_1074;
  assign _EVAL_133 = _EVAL_766 & _EVAL_1603;
  assign _EVAL_1704 = _EVAL_1502[14:12];
  assign _EVAL_1774 = _EVAL_1726 | _EVAL_1909;
  assign _EVAL_557 = _EVAL_1325 & _EVAL_1936;
  assign _EVAL_37 = _EVAL_36;
  assign _EVAL_1703 = _EVAL_636 & _EVAL_1086;
  assign _EVAL_763 = _EVAL_1717 & _EVAL_223;
  assign _EVAL_1410 = _EVAL_315 == 10'h100;
  assign _EVAL_1443 = _EVAL_1141 ? _EVAL_959 : _EVAL_1202;
  assign _EVAL_1515 = _EVAL_1130 & _EVAL_959;
  assign _EVAL_783 = _EVAL_1448 | _EVAL_963;
  assign _EVAL_1868 = _EVAL_1757 | _EVAL_219;
  assign _EVAL_227 = _EVAL_423 & _EVAL_854;
  assign _EVAL_925 = {_EVAL_749,_EVAL_1063,_EVAL_545,_EVAL_664};
  assign _EVAL_898 = _EVAL_1016 & _EVAL_116;
  assign _EVAL_1689 = _EVAL_1139 ? _EVAL_2002 : _EVAL_1406;
  assign _EVAL_116 = &_EVAL_736;
  assign _EVAL_204 = 9'hd0 == _EVAL_351;
  assign _EVAL_605 = 6'h27 == _EVAL_1978;
  assign _EVAL_1959 = _EVAL_1327 & _EVAL_1127;
  assign _EVAL_998 = _EVAL_400 & _EVAL_1575;
  assign _EVAL_1367 = _EVAL_521 & _EVAL_1773;
  assign _EVAL_707 = _EVAL_1641 & _EVAL_1458;
  assign _EVAL_1128 = _EVAL_1577 ? 8'hff : 8'h0;
  assign _EVAL_1679 = _EVAL_876 ? _EVAL_1863 : _EVAL_139;
  assign _EVAL_1124 = {{10'd0}, _EVAL_188};
  assign _EVAL_1738 = _EVAL_282 ? _EVAL_1740 : _EVAL_700;
  assign _EVAL_1282 = ~_EVAL_1904;
  assign _EVAL_1740 = {_EVAL_980,_EVAL_713,_EVAL_1828,_EVAL_1011};
  assign _EVAL_1940 = &_EVAL_1704;
  assign _EVAL_2047 = _EVAL_797 & _EVAL_177;
  assign _EVAL_1532 = _EVAL_996 & _EVAL_1971;
  assign _EVAL_1286 = _EVAL_1581 != 4'h0;
  assign _EVAL_572 = _EVAL_229 & _EVAL_1522;
  assign _EVAL_339 = _EVAL_635 | _EVAL_685;
  assign _EVAL_2045 = _EVAL_343 == 10'h0;
  assign _EVAL_1805 = _EVAL_311 & _EVAL_1001;
  assign _EVAL_2041 = _EVAL_413 & _EVAL_177;
  assign _EVAL_1577 = _EVAL_43[3];
  assign _EVAL_1062 = _EVAL_1887 & _EVAL_1086;
  assign _EVAL_1729 = _EVAL_484 & _EVAL_1173;
  assign _EVAL_834 = _EVAL_1102 ? 32'h347413 : _EVAL_501;
  assign _EVAL_1591 = _EVAL_939[9];
  assign _EVAL_1455 = ~sb2tlOpt__EVAL;
  assign _EVAL_1798 = _EVAL_474 ? 32'h7b202473 : _EVAL_1579;
  assign _EVAL_1061 = _EVAL_1717 & _EVAL_1458;
  assign _EVAL_1770 = _EVAL_400 & _EVAL_1239;
  assign _EVAL_1751 = {_EVAL_1732,1'h0,1'h0,1'h0,1'h0,_EVAL_1007,_EVAL_1007,_EVAL_566,_EVAL_566,8'ha2};
  assign _EVAL_1307 = _EVAL_691 & _EVAL_1603;
  assign _EVAL_787 = _EVAL_876 ? _EVAL_959 : _EVAL_1389;
  assign _EVAL_162 = _EVAL_939[3];
  assign _EVAL_567 = _EVAL_1016 & _EVAL_1458;
  assign _EVAL_1343 = _EVAL_1888 & _EVAL_177;
  assign _EVAL_1240 = _EVAL_1923 & _EVAL_959;
  assign _EVAL_1915 = _EVAL_1131 & _EVAL_1094;
  assign _EVAL_2037 = _EVAL_1884 & _EVAL_1074;
  assign _EVAL_1289 = _EVAL_114 & _EVAL_1001;
  assign _EVAL_479 = _EVAL_1256 & _EVAL_494;
  assign _EVAL_1236 = _EVAL_290 & _EVAL_494;
  assign _EVAL_305 = 6'h26 == _EVAL_1978;
  assign _EVAL_935 = _EVAL_859 & _EVAL_1603;
  assign _EVAL_511 = _EVAL_1515 & _EVAL_1773;
  assign _EVAL_1975 = _EVAL_1111 | _EVAL_1058;
  assign _EVAL_428 = _EVAL_748 ? 32'h10802423 : _EVAL_203;
  assign _EVAL_1575 = _EVAL_1333[212];
  assign _EVAL_1817 = _EVAL_1376 ? _EVAL_1086 : _EVAL_1808;
  assign _EVAL_2008 = _EVAL_852 ? _EVAL_959 : _EVAL_374;
  assign _EVAL_870 = _EVAL_1109 ? 1'h0 : _EVAL_1623;
  assign _EVAL_1578 = _EVAL_1327 ? 1'h0 : _EVAL_570;
  assign _EVAL_1614 = _EVAL_1232 ? _EVAL_1086 : 1'h1;
  assign _EVAL_1475 = _EVAL_168 & _EVAL_1074;
  assign _EVAL_450 = _EVAL_1113 & _EVAL_1086;
  assign _EVAL_1498 = _EVAL_586[57];
  assign _EVAL_1040 = _EVAL_756[23:0];
  assign _EVAL_1249 = _EVAL_1087 & _EVAL_481;
  assign _EVAL_186 = _EVAL_1477 ? 32'h0 : _EVAL_173;
  assign _EVAL_904 = _EVAL_51 & _EVAL_19;
  assign _EVAL_1835 = _EVAL_498 & _EVAL_1305;
  assign _EVAL_0 = {{2'd0}, _EVAL_1876};
  assign _EVAL_1863 = {_EVAL_1922,_EVAL_1882,_EVAL_1723,_EVAL_1722};
  assign _EVAL_1400 = _EVAL_1140 & _EVAL_137;
  assign _EVAL_1885 = _EVAL_14;
  assign _EVAL_103 = _EVAL_1052 ? _EVAL_1705 : _EVAL_79;
  assign _EVAL_830 = {5'h10,_EVAL_1124};
  assign _EVAL_836 = _EVAL_1416[4];
  assign _EVAL_1441 = _EVAL_1565[2];
  assign _EVAL_1956 = _EVAL_1201 & _EVAL_45;
  assign _EVAL_422 = _EVAL_1325 & _EVAL_923;
  assign _EVAL_1409 = _EVAL_237 & _EVAL_1074;
  assign _EVAL_1607 = _EVAL_1054 | _EVAL_71;
  assign _EVAL_1925 = _EVAL_585 & _EVAL_1762;
  assign _EVAL_1582 = _EVAL_586[47];
  assign _EVAL_1130 = _EVAL_400 & _EVAL_1138;
  assign _EVAL_1537 = _EVAL_1380 & _EVAL_494;
  assign _EVAL_699 = _EVAL_1683 | _EVAL_784;
  assign _EVAL_1275 = _EVAL_1108 ? _EVAL_959 : _EVAL_1412;
  assign _EVAL_1474 = _EVAL_1565[3];
  assign _EVAL_1845 = _EVAL_1730 & _EVAL_274;
  assign _EVAL_1376 = 6'h22 == _EVAL_1978;
  assign _EVAL_331 = _EVAL_568 ? 1'h0 : 1'h1;
  assign _EVAL_1406 = _EVAL_564 ? _EVAL_925 : _EVAL_1657;
  assign _EVAL_1071 = _EVAL_1140 & _EVAL_187;
  assign _EVAL_1297 = 6'h16 == _EVAL_1978;
  assign _EVAL_280 = _EVAL_1139 ? _EVAL_959 : _EVAL_906;
  assign _EVAL_974 = _EVAL_991 | _EVAL_302;
  assign _EVAL_154 = _EVAL_544 & _EVAL_494;
  assign _EVAL_1839 = ~sb2tlOpt__EVAL_19;
  assign _EVAL_1333 = 512'h1 << _EVAL_351;
  assign _EVAL_192 = _EVAL_1325 & _EVAL_137;
  assign _EVAL_726 = _EVAL_724 & _EVAL_1522;
  assign sb2tlOpt__EVAL_9 = _EVAL_38;
  assign _EVAL_789 = _EVAL_676 | _EVAL_814;
  assign _EVAL_393 = ~_EVAL_1823;
  assign _EVAL_689 = 6'h0 == _EVAL_1978;
  assign _EVAL_1784 = _EVAL_763 | _EVAL_63;
  assign _EVAL_1300 = _EVAL_2033 | _EVAL_1977;
  assign _EVAL_475 = _EVAL_1502[19:17];
  assign _EVAL_1078 = _EVAL_1416[9];
  assign _EVAL_304 = _EVAL_1552 & _EVAL_1603;
  assign _EVAL_441 = _EVAL_1108 ? 32'h40863 : _EVAL_1798;
  assign _EVAL_443 = _EVAL_690 & _EVAL_494;
  assign _EVAL_1765 = _EVAL_432 | _EVAL_1667;
  assign _EVAL_1775 = _EVAL_1502[31:16];
  assign _EVAL_992 = _EVAL_1745 ? 3'h4 : _EVAL_463;
  assign _EVAL_691 = _EVAL_425 & _EVAL_223;
  assign _EVAL_742 = _EVAL_141 | _EVAL_1423;
  assign _EVAL_66 = _EVAL_1196 & _EVAL_1224;
  assign _EVAL_190 = _EVAL_104 & _EVAL_959;
  assign _EVAL_1657 = _EVAL_1660 ? _EVAL_1188 : _EVAL_1261;
  assign _EVAL_359 = _EVAL_418 & _EVAL_1086;
  assign _EVAL_229 = _EVAL_1533 & _EVAL_1086;
  assign _EVAL_249 = _EVAL_466 ? _EVAL_1086 : _EVAL_354;
  assign _EVAL_1762 = &_EVAL_723;
  assign _EVAL_41 = _EVAL_33;
  assign _EVAL_1088 = _EVAL_1158 & _EVAL_393;
  assign _EVAL_737 = _EVAL_1815[9:0];
  assign _EVAL_462 = _EVAL_311 & _EVAL_494;
  assign _EVAL_1281 = _EVAL_1297 ? {{3'd0}, _EVAL_830} : _EVAL_621;
  assign _EVAL_593 = _EVAL_1028 & _EVAL_1603;
  assign _EVAL_597 = _EVAL_247 & _EVAL_494;
  assign _EVAL_1473 = 9'hdb == _EVAL_351;
  assign _EVAL_148 = _EVAL_536 ? _EVAL_959 : _EVAL_1443;
  assign _EVAL_1147 = _EVAL_1220 ? _EVAL_1188 : _EVAL_926;
  assign _EVAL_262 = _EVAL_566 | _EVAL_446;
  assign _EVAL_264 = _EVAL_586[33];
  assign _EVAL_413 = _EVAL_956 & _EVAL_959;
  assign _EVAL_839 = _EVAL_115 | _EVAL_344;
  assign _EVAL_1539 = _EVAL_521 & _EVAL_177;
  assign _EVAL_741 = _EVAL_1473 ? _EVAL_347 : _EVAL_1679;
  assign _EVAL_1519 = _EVAL_1448 & _EVAL_1603;
  assign _EVAL_876 = 9'hdc == _EVAL_351;
  assign _EVAL_1272 = _EVAL_1388 ? _EVAL_959 : _EVAL_1336;
  assign _EVAL_1643 = _EVAL_653 ? _EVAL_1863 : _EVAL_540;
  assign _EVAL_1435 = _EVAL_400 & _EVAL_895;
  assign _EVAL_875 = _EVAL_505 | _EVAL_1289;
  assign _EVAL_1142 = 9'h102 == _EVAL_351;
  assign _EVAL_1446 = _EVAL_643 | _EVAL_1350;
  assign _EVAL_753 = _EVAL_228 & _EVAL_1603;
  assign _EVAL_1961 = {_EVAL_684,_EVAL_397,_EVAL_855,_EVAL_1048};
  assign _EVAL_959 = _EVAL_315 == 10'h0;
  assign _EVAL_482 = _EVAL_1473 ? _EVAL_959 : _EVAL_787;
  assign _EVAL_562 = _EVAL_984 | _EVAL_1559;
  assign _EVAL_1227 = _EVAL_2001 & _EVAL_116;
  assign _EVAL_2035 = _EVAL_247 & _EVAL_854;
  assign _EVAL_794 = _EVAL_328 ? 32'h0 : _EVAL_1934;
  assign sb2tlOpt__EVAL_26 = _EVAL_8;
  assign _EVAL_1826 = 6'h21 == _EVAL_1978;
  assign _EVAL_191 = _EVAL_400 & _EVAL_1807;
  assign _EVAL_1546 = _EVAL_1271 | _EVAL_1875;
  assign _EVAL_1979 = _EVAL_1126 | _EVAL_892;
  assign _EVAL_1485 = _EVAL_1703 & _EVAL_223;
  assign _EVAL_1490 = _EVAL_1421 ? _EVAL_959 : _EVAL_500;
  assign _EVAL_84 = _EVAL_1703 & _EVAL_1971;
  assign _EVAL_516 = _EVAL_144 | _EVAL_1262;
  assign _EVAL_195 = _EVAL_32[3];
  assign _EVAL_639 = _EVAL_1285 == 3'h3;
  assign _EVAL_1895 = _EVAL_127 ? 32'h100073 : 32'h0;
  assign _EVAL_934 = _EVAL_1325 & _EVAL_150;
  assign _EVAL_669 = _EVAL_1534 & _EVAL_1603;
  assign _EVAL_555 = 6'h2b == _EVAL_1978;
  assign _EVAL_635 = _EVAL_626 & _EVAL_1458;
  assign _EVAL_2018 = _EVAL_200 == 7'h40;
  assign _EVAL_243 = _EVAL_1653 ? _EVAL_1749 : _EVAL_1281;
  assign _EVAL_231 = _EVAL_1974 ? 32'h380006f : _EVAL_1711;
  assign _EVAL_1627 = _EVAL_555 ? _EVAL_1086 : _EVAL_868;
  assign _EVAL_485 = _EVAL_1376 ? _EVAL_925 : _EVAL_1147;
  assign _EVAL_1298 = _EVAL_263 | _EVAL_1486;
  assign _EVAL_1982 = _EVAL_523 | _EVAL_407;
  assign _EVAL_837 = _EVAL_450 & _EVAL_1971;
  assign _EVAL_1331 = _EVAL_972 & _EVAL_1928;
  assign _EVAL_621 = _EVAL_1314 ? _EVAL_2025 : _EVAL_1768;
  assign _EVAL_1288 = _EVAL_417 ? _EVAL_959 : _EVAL_1238;
  assign _EVAL_134 = {{120'd0}, _EVAL_430};
  assign _EVAL_1471 = _EVAL_898 | _EVAL_462;
  assign _EVAL_939 = _EVAL_54[11:2];
  assign _EVAL_705 = _EVAL_1062 & _EVAL_494;
  assign _EVAL_618 = _EVAL_1375 & _EVAL_1603;
  assign _EVAL_1016 = _EVAL_1400 & _EVAL_1086;
  assign _EVAL_1505 = _EVAL_996 & _EVAL_116;
  assign _EVAL_1687 = _EVAL_1724 ? _EVAL_285 : _EVAL_1644;
  assign _EVAL_1368 = _EVAL_1502[16];
  assign _EVAL_1461 = _EVAL_516 & _EVAL_1824;
  assign _EVAL_823 = _EVAL_345 & _EVAL_1773;
  assign _EVAL_436 = _EVAL_1079 ? _EVAL_1329 : _EVAL_1399;
  assign _EVAL_660 = _EVAL_2031 | _EVAL_801;
  assign _EVAL_426 = _EVAL_1641 & _EVAL_116;
  assign _EVAL_127 = 9'h114 == _EVAL_351;
  assign _EVAL_98 = _EVAL_670 & _EVAL_1522;
  assign _EVAL_245 = _EVAL_135 & _EVAL_1603;
  assign _EVAL_1202 = _EVAL_1079 ? _EVAL_959 : _EVAL_241;
  assign _EVAL_1859 = _EVAL_287 & _EVAL_177;
  assign _EVAL_347 = {_EVAL_856,_EVAL_1664,_EVAL_1192,_EVAL_1211};
  assign _EVAL_1804 = _EVAL_883 & _EVAL_1603;
  assign _EVAL_585 = _EVAL_1706 & _EVAL_1086;
  assign _EVAL_1276 = _EVAL_528 ? 32'h10802023 : _EVAL_73;
  assign _EVAL_1045 = _EVAL_586[45];
  assign _EVAL_1154 = &_EVAL_1368;
  assign _EVAL_1596 = _EVAL_544 & _EVAL_854;
  assign _EVAL_288 = _EVAL_821 | _EVAL_1881;
  assign _EVAL_1632 = _EVAL_1327 & _EVAL_841;
  assign _EVAL_1345 = _EVAL_1355 | _EVAL_692;
  assign _EVAL_984 = _EVAL_1641 & _EVAL_1971;
  assign _EVAL_1336 = _EVAL_1349 ? _EVAL_959 : _EVAL_751;
  assign _EVAL_1256 = _EVAL_1153 & _EVAL_1086;
  assign _EVAL_496 = _EVAL_1612 ? _EVAL_959 : _EVAL_2042;
  assign _EVAL_1965 = _EVAL_400 & _EVAL_356;
  assign _EVAL_1984 = _EVAL_1848 ? 1'h0 : _EVAL_1489;
  assign _EVAL_1399 = _EVAL_1929 ? _EVAL_1998 : _EVAL_741;
  assign _EVAL_907 = _EVAL_1333[209];
  assign _EVAL_825 = _EVAL_767 & _EVAL_1971;
  assign _EVAL_1337 = 6'h4 == _EVAL_1978;
  assign _EVAL_914 = _EVAL_586[22];
  assign _EVAL_345 = _EVAL_1965 & _EVAL_959;
  assign _EVAL_498 = sb2tlOpt__EVAL_11 | sb2tlOpt__EVAL_1;
  assign _EVAL_29 = _EVAL_688 ? _EVAL_775 : 32'h0;
  assign _EVAL_717 = _EVAL_1906 & _EVAL_1603;
  assign _EVAL_491 = _EVAL_1888 & _EVAL_1928;
  assign _EVAL_1808 = _EVAL_1220 ? _EVAL_1086 : _EVAL_896;
  assign _EVAL_534 = _EVAL_1392 & _EVAL_1282;
  assign _EVAL_871 = _EVAL_1219 & _EVAL_1773;
  assign _EVAL_1877 = _EVAL_40[31:24];
  assign _EVAL_412 = &_EVAL_1987;
  assign _EVAL_1615 = _EVAL_544 & _EVAL_1001;
  assign _EVAL_1036 = _EVAL_725 | _EVAL_1159;
  assign _EVAL_1824 = ~_EVAL_1603;
  assign _EVAL_1978 = {_EVAL_1642,_EVAL_817,_EVAL_1474,_EVAL_1441,_EVAL_631,_EVAL_964};
  assign _EVAL_1718 = _EVAL_648 | _EVAL_169;
  assign _EVAL_665 = _EVAL_1140 & _EVAL_778;
  assign _EVAL_1986 = _EVAL_1325 & _EVAL_89;
  assign _EVAL_677 = _EVAL_1702[127:0];
  assign _EVAL_1848 = _EVAL_288 & _EVAL_1823;
  assign _EVAL_1074 = &_EVAL_949;
  assign _EVAL_1880 = _EVAL_972 & _EVAL_1773;
  assign _EVAL_1823 = _EVAL_1663 | _EVAL_1162;
  assign _EVAL_2042 = _EVAL_282 ? _EVAL_959 : _EVAL_1068;
  assign _EVAL_1013 = _EVAL_1769 | _EVAL_464;
  assign _EVAL_1900 = _EVAL_2025[17];
  assign _EVAL_2025 = {_EVAL_1853,_EVAL_1989};
  assign _EVAL_1948 = _EVAL_556 & _EVAL_1599;
  assign _EVAL_1207 = _EVAL_709 & _EVAL_1074;
  assign _EVAL_281 = _EVAL_605 ? _EVAL_1358 : _EVAL_103;
  assign _EVAL_1796 = _EVAL_1416[10];
  assign _EVAL_756 = _EVAL_228 ? _EVAL_39 : 32'h0;
  assign _EVAL_690 = _EVAL_422 & _EVAL_1086;
  assign _EVAL_1177 = _EVAL_821 ? _EVAL_39 : 32'h0;
  assign _EVAL_2052 = _EVAL_114 & _EVAL_854;
  assign _EVAL_880 = _EVAL_858 & _EVAL_1286;
  assign _EVAL_642 = _EVAL_1077 ? _EVAL_1410 : _EVAL_1419;
  assign _EVAL_203 = _EVAL_852 ? 32'h7b202473 : _EVAL_1209;
  assign _EVAL_112 = _EVAL_1028 | _EVAL_961;
  assign _EVAL_671 = _EVAL_939[2];
  assign _EVAL_1488 = _EVAL_1348 & _EVAL_1603;
  assign _EVAL_1015 = _EVAL_1648 & _EVAL_1603;
  assign _EVAL_1224 = _EVAL_625 == 3'h0;
  assign _EVAL_525 = _EVAL_1532 | _EVAL_1992;
  assign _EVAL_1985 = _EVAL_271 & _EVAL_223;
  assign _EVAL_374 = _EVAL_846 ? _EVAL_959 : _EVAL_565;
  assign _EVAL_1325 = _EVAL_1183 & _EVAL_1452;
  assign _EVAL_1371 = _EVAL_837 | _EVAL_439;
  assign _EVAL_1732 = _EVAL_1346 ? _EVAL_1249 : _EVAL_1087;
  assign _EVAL_716 = _EVAL_766 | _EVAL_1537;
  assign _EVAL_546 = _EVAL_1349 ? 32'h7b241073 : _EVAL_1847;
  assign _EVAL_1378 = _EVAL_503 ? 8'hff : 8'h0;
  assign _EVAL_1350 = _EVAL_247 & _EVAL_1001;
  assign _EVAL_1640 = _EVAL_1888 & _EVAL_1074;
  assign _EVAL_848 = _EVAL_1693 & _EVAL_363;
  assign _EVAL_1044 = _EVAL_1485 & _EVAL_1603;
  assign _EVAL_1561 = _EVAL_1682 | _EVAL_319;
  assign _EVAL_1084 = _EVAL_2033 & _EVAL_1603;
  assign _EVAL_791 = _EVAL_382 ? _EVAL_1961 : _EVAL_1251;
  assign _EVAL_846 = 9'h112 == _EVAL_351;
  assign _EVAL_1239 = _EVAL_1333[222];
  assign _EVAL_954 = _EVAL_358 ? _EVAL_199 : _EVAL_517;
  assign _EVAL_484 = _EVAL_353 | _EVAL_131;
  assign _EVAL_2002 = {_EVAL_1384,_EVAL_754,_EVAL_372,_EVAL_578};
  assign _EVAL_532 = _EVAL_611 | _EVAL_1254;
  assign _EVAL_67 = _EVAL_400 & _EVAL_369;
  assign _EVAL_978 = ~_EVAL_1900;
  assign _EVAL_1059 = _EVAL_1219 & _EVAL_1928;
  assign _EVAL_247 = _EVAL_146 & _EVAL_1086;
  assign _EVAL_1466 = _EVAL_563 | _EVAL_575;
  assign _EVAL_434 = _EVAL_1325 & _EVAL_2009;
  assign _EVAL_140 = {64'h0,32'h0,_EVAL_448,_EVAL_1520,_EVAL_1273,_EVAL_1230};
  assign _EVAL_187 = _EVAL_586[60];
  assign _EVAL_94 = _EVAL_248 & _EVAL_1603;
  assign _EVAL_1653 = 6'h13 == _EVAL_1978;
  assign _EVAL_521 = _EVAL_1944 & _EVAL_959;
  assign _EVAL_1352 = _EVAL_1140 & _EVAL_538;
  assign _EVAL_287 = _EVAL_1756 & _EVAL_959;
  assign _EVAL_1032 = _EVAL_1038 | _EVAL_1583;
  assign _EVAL_156 = _EVAL_543 & _EVAL_1073;
  assign _EVAL_1012 = &_EVAL_1502;
  assign _EVAL_568 = _EVAL_978 | _EVAL_326;
  assign _EVAL_564 = 9'hd2 == _EVAL_351;
  assign _EVAL_1204 = _EVAL_1504 ? _EVAL_959 : _EVAL_230;
  assign _EVAL_470 = _EVAL_392 | _EVAL_779;
  assign _EVAL_1109 = ~_EVAL_20;
  assign _EVAL_261 = _EVAL_797 & _EVAL_1928;
  assign _EVAL_1681 = 6'h29 == _EVAL_1978;
  assign _EVAL_464 = _EVAL_848 & _EVAL_1824;
  assign _EVAL_410 = _EVAL_789 | _EVAL_1868;
  assign _EVAL_213 = _EVAL_1468 ? _EVAL_1086 : _EVAL_342;
  assign _EVAL_1887 = _EVAL_1325 & _EVAL_264;
  assign _EVAL_901 = _EVAL_1730 ? _EVAL_1144 : _EVAL_1009;
  assign _EVAL_1326 = _EVAL_182 & _EVAL_1773;
  assign _EVAL_244 = _EVAL_1985 & _EVAL_1603;
  assign _EVAL_76 = _EVAL_1022 | _EVAL_2039;
  assign _EVAL_1953 = 9'h43 == _EVAL_351;
  assign _EVAL_418 = _EVAL_1140 & _EVAL_1498;
  assign _EVAL_628 = _EVAL_1314 ? _EVAL_1086 : _EVAL_1758;
  assign _EVAL_523 = _EVAL_1016 & _EVAL_223;
  assign _EVAL_649 = _EVAL_39[15];
  assign _EVAL_389 = _EVAL_271 & _EVAL_1458;
  assign _EVAL_258 = _EVAL_1660 ? _EVAL_959 : _EVAL_1812;
  assign _EVAL_1964 = _EVAL_586[46];
  assign _EVAL_1133 = _EVAL_608 & 12'h1;
  assign _EVAL_174 = _EVAL_1612 ? _EVAL_1961 : _EVAL_1738;
  assign _EVAL_283 = _EVAL_1168 ? _EVAL_959 : _EVAL_1275;
  assign _EVAL_1420 = _EVAL_40[7:0];
  assign _EVAL_1189 = _EVAL_974 | _EVAL_296;
  assign _EVAL_343 = _EVAL_40[9:0];
  assign _EVAL_284 = _EVAL_1416[13];
  assign _EVAL_1849 = _EVAL_301 ? {{9'd0}, _EVAL_1567} : _EVAL_243;
  assign _EVAL_447 = _EVAL_1379 | _EVAL_973;
  assign _EVAL_1418 = _EVAL_848 & _EVAL_1603;
  assign _EVAL_986 = _EVAL_532 | _EVAL_76;
  assign _EVAL_242 = {64'h0,32'h0,_EVAL_1177};
  assign _EVAL_271 = _EVAL_661 & _EVAL_1086;
  assign _EVAL_712 = _EVAL_234 & _EVAL_1086;
  assign _EVAL_1790 = _EVAL_1333[66];
  assign _EVAL_356 = _EVAL_1333[221];
  assign _EVAL_1111 = _EVAL_1813 | _EVAL_1446;
  assign _EVAL_743 = _EVAL_307 == 3'h0;
  assign _EVAL_850 = _EVAL_1026 & _EVAL_1603;
  assign _EVAL_1712 = _EVAL_2025[15:0];
  assign _EVAL_1713 = _EVAL_400 & _EVAL_449;
  assign _EVAL_1200 = {{5'd0}, _EVAL_793};
  assign _EVAL_1181 = _EVAL_1416[2];
  assign _EVAL_432 = _EVAL_1014 | _EVAL_156;
  assign _EVAL_1364 = _EVAL_920 & _EVAL_1928;
  assign _EVAL_1962 = _EVAL_586[32];
  assign _EVAL_352 = _EVAL_426 | _EVAL_1396;
  assign _EVAL_1372 = _EVAL_1033 & _EVAL_1086;
  assign _EVAL_1301 = _EVAL_400 & _EVAL_1795;
  assign _EVAL_908 = _EVAL_686 | _EVAL_673;
  assign _EVAL_632 = 9'hde == _EVAL_351;
  assign _EVAL_956 = _EVAL_400 & _EVAL_552;
  assign _EVAL_1719 = _EVAL_1025 | _EVAL_537;
  assign _EVAL_595 = _EVAL_159 | _EVAL_507;
  assign _EVAL_1819 = _EVAL_300 ? 1'h0 : _EVAL_1600;
  assign _EVAL_360 = 9'hdd == _EVAL_351;
  assign _EVAL_1545 = _EVAL_237 & _EVAL_1928;
  assign _EVAL_686 = _EVAL_1507 | _EVAL_456;
  assign _EVAL_285 = {_EVAL_506,_EVAL_2032,_EVAL_1483,_EVAL_333};
  assign _EVAL_263 = _EVAL_1090 | _EVAL_1371;
  assign _EVAL_1283 = _EVAL_1036 & _EVAL_429;
  assign _EVAL_1522 = |_EVAL_1361;
  assign _EVAL_1683 = _EVAL_286 & _EVAL_1458;
  assign _EVAL_1053 = _EVAL_803 ? _EVAL_959 : _EVAL_283;
  assign _EVAL_1099 = _EVAL_1219 & _EVAL_177;
  assign _EVAL_1641 = _EVAL_1677 & _EVAL_1086;
  assign _EVAL_887 = _EVAL_825 & _EVAL_1603;
  assign _EVAL_2027 = _EVAL_1606 | _EVAL_1767;
  assign _EVAL_1503 = _EVAL_1416[5];
  assign _EVAL_1094 = _EVAL_1712 <= 16'h101f;
  assign _EVAL_1269 = {{1'd0}, _EVAL_603};
  assign _EVAL_420 = _EVAL_635 & _EVAL_1603;
  assign _EVAL_813 = _EVAL_1502[22];
  assign _EVAL_129 = _EVAL_39[19:17];
  assign _EVAL_949 = _EVAL_1815[23:16];
  assign _EVAL_1715 = _EVAL_39[7:0];
  assign _EVAL_1944 = _EVAL_400 & _EVAL_907;
  assign _EVAL_1702 = _EVAL_295 + _EVAL_134;
  assign _EVAL_592 = _EVAL_1605 & _EVAL_1154;
  assign _EVAL_2015 = _EVAL_1603 ? 1'h0 : _EVAL_1632;
  assign _EVAL_966 = _EVAL_32[0];
  assign _EVAL_502 = _EVAL_1678 | _EVAL_550;
  assign _EVAL_892 = _EVAL_1264 | _EVAL_443;
  assign _EVAL_1717 = _EVAL_755 & _EVAL_1086;
  assign _EVAL_64 = _EVAL_1931 ? _EVAL_1086 : _EVAL_1627;
  assign _EVAL_60 = _EVAL_1416[3];
  assign _EVAL_1791 = _EVAL_972 & _EVAL_1074;
  assign _EVAL_888 = _EVAL_996 & _EVAL_1458;
  assign _EVAL_453 = _EVAL_1325 & _EVAL_538;
  assign _EVAL_1648 = _EVAL_240 & _EVAL_223;
  assign _EVAL_1390 = _EVAL_400 & _EVAL_1790;
  assign _EVAL_793 = {1'h0,_EVAL_1904,_EVAL_768,_EVAL_274,_EVAL_1285,_EVAL_1305,_EVAL_1304,_EVAL_307,12'h407};
  assign _EVAL_118 = _EVAL_1996 | _EVAL_1596;
  assign _EVAL_1783 = _EVAL_648 & _EVAL_1603;
  assign _EVAL_202 = _EVAL_1375 & _EVAL_1824;
  assign _EVAL_1136 = _EVAL_39[31:16];
  assign _EVAL_1458 = &_EVAL_1180;
  assign _EVAL_1459 = _EVAL_1146 ? _EVAL_959 : _EVAL_217;
  assign _EVAL_868 = _EVAL_653 ? _EVAL_1086 : _EVAL_213;
  assign _EVAL_1046 = _EVAL_196[0];
  assign _EVAL_1917 = &_EVAL_813;
  assign _EVAL_1866 = _EVAL_1374 & _EVAL_1466;
  assign _EVAL_1425 = ~_EVAL_437;
  assign _EVAL_1370 = _EVAL_1416[8];
  assign _EVAL_895 = _EVAL_1333[213];
  assign _EVAL_12 = {{2'd0}, _EVAL_1452};
  assign _EVAL_1876 = _EVAL_9 == 3'h4;
  assign _EVAL_364 = &_EVAL_475;
  assign _EVAL_1431 = _EVAL_1605 & _EVAL_364;
  assign _EVAL_421 = _EVAL_2014 & _EVAL_865;
  assign _EVAL_1929 = 9'hda == _EVAL_351;
  assign _EVAL_1927 = _EVAL_1325 & _EVAL_444;
  assign _EVAL_222 = _EVAL_979 | _EVAL_278;
  assign _EVAL_1996 = _EVAL_2001 & _EVAL_1971;
  assign _EVAL_1187 = _EVAL_225 & _EVAL_481;
  assign _EVAL_1579 = _EVAL_1811 ? 32'h10002223 : _EVAL_761;
  assign _EVAL_2033 = _EVAL_450 & _EVAL_1458;
  assign _EVAL_1846 = _EVAL_604[1];
  assign _EVAL_510 = _EVAL_1957 | _EVAL_1236;
  assign _EVAL_926 = _EVAL_1920 ? _EVAL_1694 : _EVAL_1675;
  assign _EVAL_698 = _EVAL_1142 ? _EVAL_959 : _EVAL_1272;
  assign _EVAL_1208 = _EVAL_1232 ? _EVAL_1414 : 32'h0;
  assign _EVAL_1209 = _EVAL_846 ? 32'h7b200073 : _EVAL_56;
  assign _EVAL_306 = _EVAL_1650 | _EVAL_339;
  assign _EVAL_920 = _EVAL_998 & _EVAL_959;
  assign _EVAL_336 = _EVAL_1140 & _EVAL_1045;
  assign _EVAL_1988 = _EVAL_1515 & _EVAL_1074;
  assign _EVAL_276 = _EVAL_298 & _EVAL_1086;
  assign _EVAL_911 = _EVAL_1416[0];
  assign _EVAL_963 = _EVAL_229 & _EVAL_1001;
  assign _EVAL_591 = 1024'h1 << _EVAL_343;
  assign _EVAL_301 = 6'h11 == _EVAL_1978;
  assign _EVAL_626 = _EVAL_1779 & _EVAL_1086;
  assign _EVAL_1588 = _EVAL_1227 & _EVAL_1603;
  assign _EVAL_1807 = _EVAL_1333[67];
  assign _EVAL_1019 = _EVAL_1629 | _EVAL_373;
  assign _EVAL_617 = _EVAL_1325 & _EVAL_1582;
  assign _EVAL_929 = _EVAL_1884 & _EVAL_177;
  assign sb2tlOpt__EVAL_25 = _EVAL_1730 ? _EVAL_1268 : _EVAL_295;
  assign _EVAL_1889 = 9'h101 == _EVAL_351;
  assign _EVAL_958 = _EVAL_1416[15];
  assign _EVAL_841 = _EVAL_1127 ? 1'h0 : _EVAL_1553;
  assign _EVAL_1238 = _EVAL_358 ? _EVAL_959 : _EVAL_1593;
  assign _EVAL_501 = _EVAL_803 ? 32'hfe0408e3 : _EVAL_390;
  assign _EVAL_1263 = 9'h41 == _EVAL_351;
  assign _EVAL_211 = _EVAL_271 & _EVAL_1971;
  assign _EVAL_1023 = _EVAL_413 & _EVAL_1074;
  assign _EVAL_603 = {1'h0,_EVAL_225,_EVAL_225,_EVAL_1732,_EVAL_1751};
  assign _EVAL_1533 = _EVAL_1325 & _EVAL_1964;
  assign _EVAL_311 = _EVAL_192 & _EVAL_1086;
  assign _EVAL_805 = _EVAL_1603 ? 1'h0 : _EVAL_1578;
  assign _EVAL_358 = 9'hcf == _EVAL_351;
  assign _EVAL_858 = _EVAL_1285 == 3'h4;
  assign _EVAL_1768 = _EVAL_740 ? _EVAL_265 : _EVAL_1369;
  assign _EVAL_915 = _EVAL_1931 ? _EVAL_1998 : _EVAL_937;
  assign _EVAL_216 = _EVAL_1035 & _EVAL_1522;
  assign _EVAL_670 = _EVAL_1986 & _EVAL_1086;
  assign _EVAL_1342 = _EVAL_891 & _EVAL_1458;
  assign _EVAL_802 = _EVAL_1925 & _EVAL_1603;
  assign _EVAL_972 = _EVAL_702 & _EVAL_959;
  assign _EVAL_832 = _EVAL_278 & _EVAL_1634;
  assign _EVAL_1038 = _EVAL_1016 & _EVAL_1971;
  assign _EVAL_538 = _EVAL_586[34];
  assign _EVAL_252 = _EVAL_2036 ? _EVAL_1009 : _EVAL_1208;
  assign _EVAL_1697 = _EVAL_39[22];
  assign _EVAL_1583 = _EVAL_311 & _EVAL_854;
  assign _EVAL_694 = _EVAL_290 & _EVAL_1522;
  assign _EVAL_1210 = _EVAL_366 & _EVAL_1688;
  assign _EVAL_395 = _EVAL_120 & _EVAL_1666;
  assign _EVAL_1587 = _EVAL_262 & _EVAL_1425;
  assign _EVAL_1513 = ~_EVAL_388;
  assign _EVAL_1468 = 6'h2d == _EVAL_1978;
  assign _EVAL_1812 = _EVAL_1042 ? _EVAL_959 : _EVAL_1459;
  assign _EVAL_1921 = _EVAL_1187 | _EVAL_563;
  assign _EVAL_544 = _EVAL_899 & _EVAL_1086;
  assign _EVAL_2 = _EVAL;
  assign _EVAL_2009 = _EVAL_586[44];
  assign _EVAL_419 = _EVAL_1884 & _EVAL_1773;
  assign _EVAL_1852 = _EVAL_797 & _EVAL_1074;
  assign _EVAL_380 = _EVAL_400 & _EVAL_890;
  assign _EVAL_549 = _EVAL_287 & _EVAL_1074;
  assign _EVAL_536 = 9'hd7 == _EVAL_351;
  assign _EVAL_427 = _EVAL_1703 & _EVAL_1458;
  assign _EVAL_141 = _EVAL_610 | _EVAL_699;
  assign _EVAL_1112 = _EVAL_1096 == 2'h2;
  assign _EVAL_1160 = _EVAL_229 & _EVAL_494;
  assign _EVAL_135 = _EVAL_1372 & _EVAL_116;
  assign _EVAL_2017 = _EVAL_1219 & _EVAL_1074;
  assign _EVAL_73 = _EVAL_1421 ? 32'h40044403 : _EVAL_834;
  assign _EVAL_340 = _EVAL_1091 & _EVAL_1001;
  assign _EVAL_417 = 9'hce == _EVAL_351;
  assign _EVAL_1861 = _EVAL_2015 | _EVAL_2051;
  assign _EVAL_2046 = _EVAL_32[2];
  assign _EVAL_1795 = _EVAL_1333[211];
  assign _EVAL_842 = _EVAL_1372 & _EVAL_1971;
  assign _EVAL_169 = _EVAL_1062 & _EVAL_854;
  assign _EVAL_1196 = _EVAL_753 & _EVAL_1659;
  assign _EVAL_863 = _EVAL_1148 & _EVAL_1603;
  assign _EVAL_2039 = _EVAL_670 & _EVAL_494;
  assign _EVAL_1946 = _EVAL_1240 & _EVAL_1666;
  assign _EVAL_1155 = _EVAL_127 ? _EVAL_959 : 1'h1;
  assign _EVAL_951 = _EVAL_1333[220];
  assign sb2tlOpt__EVAL_12 = _EVAL_1088 & _EVAL_117;
  assign _EVAL_1392 = _EVAL_821 & _EVAL_865;
  assign _EVAL_773 = _EVAL_1296 | _EVAL_562;
  assign _EVAL_885 = _EVAL_1189 | _EVAL_680;
  assign _EVAL_1629 = _EVAL_288 & _EVAL_1460;
  assign _EVAL_541 = _EVAL_946 | _EVAL_525;
  assign _EVAL_25 = _EVAL_6;
  assign _EVAL_497 = _EVAL_182 & _EVAL_177;
  assign _EVAL_575 = _EVAL_1886 & _EVAL_1007;
  assign _EVAL_1516 = _EVAL_767 & _EVAL_1458;
  assign _EVAL_927 = _EVAL_742 | _EVAL_543;
  assign _EVAL_1460 = _EVAL_105 | _EVAL_880;
  assign _EVAL_375 = _EVAL_400 & _EVAL_1321;
  assign _EVAL_1257 = _EVAL_1603 ? _EVAL_1819 : _EVAL_1959;
  assign _EVAL_1603 = _EVAL_1096 == 2'h0;
  assign _EVAL_184 = _EVAL_643 & _EVAL_1603;
  assign _EVAL_1553 = _EVAL_332 ? 1'h0 : 1'h1;
  assign _EVAL_1811 = 9'h10d == _EVAL_351;
  assign _EVAL_715 = _EVAL_1264 & _EVAL_1603;
  assign _EVAL_1726 = _EVAL_276 & _EVAL_1458;
  assign _EVAL_1544 = _EVAL_1077 ? {{16'd0}, _EVAL_1244} : _EVAL_186;
  assign _EVAL_1105 = _EVAL_1884 & _EVAL_1928;
  assign _EVAL_309 = _EVAL_1707 | _EVAL_694;
  assign _EVAL_300 = _EVAL_66 | _EVAL_334;
  assign _EVAL_781 = _EVAL_2036 ? _EVAL_1086 : _EVAL_1614;
  assign _EVAL_1264 = _EVAL_1717 & _EVAL_116;
  assign _EVAL_80 = _EVAL_438 | _EVAL_811;
  assign _EVAL_125 = _EVAL_724 & _EVAL_1001;
  assign _EVAL_1452 = _EVAL_3 == 3'h4;
  assign _EVAL_1638 = _EVAL_1648 | _EVAL_454;
  assign _EVAL_1241 = _EVAL_984 & _EVAL_1603;
  assign _EVAL_2028 = _EVAL_690 & _EVAL_1001;
  assign _EVAL_775 = _EVAL_689 ? _EVAL_782 : _EVAL_1973;
  assign _EVAL_1448 = _EVAL_425 & _EVAL_1458;
  assign _EVAL_1123 = _EVAL_1026 | _EVAL_1834;
  assign _EVAL_1847 = _EVAL_894 ? 32'hf1402473 : _EVAL_1276;
  assign _EVAL_1000 = _EVAL_1177[15:8];
  assign _EVAL_1057 = _EVAL_1785 & _EVAL_1304;
  assign _EVAL_767 = _EVAL_548 & _EVAL_1086;
  assign _EVAL_52 = _EVAL_19;
  assign _EVAL_803 = 9'h109 == _EVAL_351;
  assign _EVAL_1262 = _EVAL_842 | _EVAL_2052;
  assign _EVAL_1220 = 6'h23 == _EVAL_1978;
  assign _EVAL_1188 = {_EVAL_379,_EVAL_308,_EVAL_1781,_EVAL_822};
  assign _EVAL_733 = _EVAL_632 ? _EVAL_959 : _EVAL_496;
  assign _EVAL_270 = _EVAL_709 & _EVAL_1928;
  assign _EVAL_981 = _EVAL_32[1];
  assign _EVAL_1348 = _EVAL_391 & _EVAL_1971;
  assign _EVAL_874 = _EVAL_1811 ? _EVAL_959 : _EVAL_732;
  assign _EVAL_610 = _EVAL_1857 | _EVAL_112;
  assign _EVAL_1322 = _EVAL_1865 | _EVAL_832;
  assign _EVAL_278 = _EVAL_1148 | _EVAL_1646;
  assign _EVAL_519 = _EVAL_235 & _EVAL_1666;
  assign _EVAL_1278 = _EVAL_1035 & _EVAL_1001;
  assign _EVAL_1158 = _EVAL_667 & _EVAL_743;
  assign _EVAL_240 = _EVAL_1864 & _EVAL_1086;
  assign _EVAL_1338 = _EVAL_240 & _EVAL_116;
  assign _EVAL_1875 = _EVAL_1256 & _EVAL_1522;
  assign _EVAL_282 = 9'he0 == _EVAL_351;
  assign _EVAL_554 = _EVAL_1815[7:0];
  assign _EVAL_751 = _EVAL_894 ? _EVAL_959 : _EVAL_1081;
  assign _EVAL_859 = _EVAL_2001 & _EVAL_1458;
  assign _EVAL_709 = _EVAL_67 & _EVAL_959;
  assign _EVAL_556 = _EVAL_1605 & _EVAL_1940;
  assign _EVAL_1976 = _EVAL_541 | _EVAL_1125;
  assign _EVAL_1108 = 9'h10b == _EVAL_351;
  assign _EVAL_86 = _EVAL_831 & _EVAL_1603;
  assign sb2tlOpt__EVAL_24 = _EVAL_50;
  assign _EVAL_1472 = _EVAL_1416[11];
  assign _EVAL_178 = _EVAL_39[31:24];
  assign _EVAL_1047 = _EVAL_1091 & _EVAL_1522;
  assign _EVAL_643 = _EVAL_240 & _EVAL_1458;
  assign _EVAL_814 = _EVAL_1061 | _EVAL_2028;
  assign _EVAL_109 = _EVAL_712 & _EVAL_854;
  assign _EVAL_1077 = 9'h0 == _EVAL_351;
  assign _EVAL_1745 = _EVAL_1603 ? 1'h0 : _EVAL_1010;
  assign _EVAL_1901 = _EVAL_773 | _EVAL_710;
  assign _EVAL_989 = _EVAL_861 & _EVAL_1603;
  assign _EVAL_316 = _EVAL_1255 & _EVAL_1603;
  assign _EVAL_1778 = _EVAL_1271 & _EVAL_1603;
  assign _EVAL_362 = _EVAL_639 & _EVAL_2050;
  assign _EVAL_854 = |_EVAL_68;
  assign _EVAL_16 = _EVAL_17;
  assign _EVAL_847 = _EVAL_892 & _EVAL_1503;
  assign _EVAL_1033 = _EVAL_1140 & _EVAL_1936;
  assign _EVAL_1605 = _EVAL_957 & _EVAL_1086;
  assign _EVAL_367 = |_EVAL_1502;
  assign _EVAL_1888 = _EVAL_1713 & _EVAL_959;
  assign _EVAL_1785 = _EVAL_1415 & _EVAL_367;
  assign _EVAL_188 = {1'h0,_EVAL_1432,1'h0,_EVAL_625,8'h1};
  assign _EVAL_1412 = _EVAL_474 ? _EVAL_959 : _EVAL_874;
  assign _EVAL_298 = _EVAL_1140 & _EVAL_1582;
  assign _EVAL_732 = _EVAL_1334 ? _EVAL_959 : _EVAL_1204;
  assign _EVAL_1974 = 9'hc0 == _EVAL_351;
  assign _EVAL_328 = 9'h42 == _EVAL_351;
  assign _EVAL_210 = _EVAL_1975 | _EVAL_1471;
  assign _EVAL_382 = 6'h2f == _EVAL_1978;
  assign _EVAL_535 = _EVAL_561 & _EVAL_1603;
  assign _EVAL_1998 = {_EVAL_1163,_EVAL_1816,_EVAL_777,_EVAL_553};
  assign _EVAL_739 = ~_EVAL_1452;
  assign _EVAL_1909 = _EVAL_290 & _EVAL_1001;
  assign _EVAL_1749 = {{31'd0}, _EVAL_1592};
  assign _EVAL_230 = _EVAL_748 ? _EVAL_959 : _EVAL_2008;
  assign _EVAL_766 = _EVAL_891 & _EVAL_116;
  assign _EVAL_2001 = _EVAL_1633 & _EVAL_1086;
  assign _EVAL_1085 = _EVAL_1826 ? _EVAL_2002 : _EVAL_485;
  assign _EVAL_608 = {{11'd0}, _EVAL_995};
  assign _EVAL_120 = _EVAL_1390 & _EVAL_959;
  assign _EVAL_1419 = _EVAL_1477 ? _EVAL_959 : _EVAL_1373;
  assign _EVAL_673 = _EVAL_352 & _EVAL_60;
  assign _EVAL_563 = hartIsInResetSync_0_debug_hartReset_0__EVAL;
  assign _EVAL_463 = _EVAL_802 ? _EVAL_1242 : _EVAL_625;
  assign _EVAL_1706 = _EVAL_1140 & _EVAL_914;
  assign _EVAL_504 = _EVAL_710 & _EVAL_836;
  assign _EVAL_1075 = _EVAL_1837 & _EVAL_1603;
  assign _EVAL_196 = _EVAL_395 ? _EVAL_591 : 1024'h0;
  assign _EVAL_1705 = {_EVAL_1118,_EVAL_1616,_EVAL_624,_EVAL_1051};
  assign _EVAL_1268 = {96'h0,_EVAL_1144};
  assign _EVAL_335 = _EVAL_1726 & _EVAL_1603;
  assign _EVAL_629 = _EVAL_920 & _EVAL_1773;
  assign _EVAL_423 = _EVAL_1933 & _EVAL_1086;
  assign _EVAL_1559 = _EVAL_1091 & _EVAL_854;
  assign _EVAL_968 = _EVAL_361 ? _EVAL_1086 : _EVAL_781;
  assign _EVAL_1050 = _EVAL_1826 ? _EVAL_1086 : _EVAL_1817;
  assign _EVAL_1558 = _EVAL_1889 ? _EVAL_959 : _EVAL_698;
  assign _EVAL_827 = _EVAL_455 | _EVAL_1774;
  assign _EVAL_600 = _EVAL_1463 & _EVAL_1697;
  assign _EVAL_327 = _EVAL_39[20];
  assign _EVAL_896 = _EVAL_1920 ? _EVAL_1086 : _EVAL_249;
  assign _EVAL_1997 = _EVAL_1052 ? _EVAL_1086 : _EVAL_1260;
  assign _EVAL_1379 = _EVAL_891 & _EVAL_223;
  assign _EVAL_1928 = &_EVAL_1716;
  assign _EVAL_964 = _EVAL_1565[0];
  assign _EVAL_319 = _EVAL_211 | _EVAL_1267;
  assign _EVAL_146 = _EVAL_1325 & _EVAL_1394;
  assign _EVAL_565 = _EVAL_1803 ? _EVAL_959 : _EVAL_1155;
  assign _EVAL_724 = _EVAL_934 & _EVAL_1086;
  assign _EVAL_1518 = ~_EVAL_1876;
  assign _EVAL_1957 = _EVAL_276 & _EVAL_116;
  assign _EVAL_1675 = _EVAL_466 ? _EVAL_476 : _EVAL_180;
  assign _EVAL_1233 = _EVAL_1848 | _EVAL_1345;
  assign _EVAL_1042 = 9'hd4 == _EVAL_351;
  assign sb2tlOpt__EVAL_27 = _EVAL_1055 & _EVAL_117;
  assign _EVAL_315 = _EVAL_939 & 10'h100;
  assign _EVAL_1599 = _EVAL_604[0];
  assign sb2tlOpt__EVAL_20 = _EVAL_18;
  assign _EVAL_124 = _EVAL_1255 | _EVAL_1083;
  assign _EVAL_1081 = _EVAL_528 ? _EVAL_959 : _EVAL_1490;
  assign _EVAL_1068 = _EVAL_785 ? _EVAL_959 : _EVAL_1558;
  assign _EVAL_1581 = _EVAL_901[3:0];
  assign _EVAL_505 = _EVAL_1372 & _EVAL_1458;
  assign _EVAL_1920 = 6'h24 == _EVAL_1978;
  assign _EVAL_425 = _EVAL_1618 & _EVAL_1086;
  assign _EVAL_1450 = _EVAL_901[2:0];
  assign _EVAL_28 = 1'h1;
  assign _EVAL_296 = _EVAL_825 | _EVAL_638;
  assign _EVAL_678 = {1'h0,_EVAL_692,_EVAL_1347,_EVAL_647};
  assign _EVAL_995 = _EVAL_39[0];
  assign _EVAL_439 = _EVAL_670 & _EVAL_854;
  assign _EVAL_648 = _EVAL_626 & _EVAL_1971;
  assign _EVAL_1131 = _EVAL_1712 >= 16'h1000;
  assign _EVAL_1295 = _EVAL_1140 & _EVAL_416;
  assign _EVAL_1290 = _EVAL_544 & _EVAL_1522;
  assign _EVAL_1730 = _EVAL_359 & _EVAL_1012;
  assign _EVAL_757 = _EVAL_677[31:0];
  assign _EVAL_1660 = 9'hd3 == _EVAL_351;
  assign _EVAL_132 = _EVAL_1317 & _EVAL_1603;
  assign _EVAL_170 = _EVAL_97 | _EVAL_80;
  assign _EVAL_1931 = 6'h2a == _EVAL_1978;
  assign _EVAL_1864 = _EVAL_1140 & _EVAL_1394;
  assign _EVAL_1568 = _EVAL_1333[224];
  assign _EVAL_991 = _EVAL_1298 | _EVAL_1072;
  assign _EVAL_1139 = 9'hd1 == _EVAL_351;
  assign _EVAL_2049 = _EVAL_43[2];
  assign sb2tlOpt__EVAL_5 = _EVAL_34;
  assign _EVAL_223 = &_EVAL_1361;
  assign _EVAL_758 = _EVAL_301 ? _EVAL_1086 : _EVAL_982;
  assign _EVAL_979 = _EVAL_839 | _EVAL_1032;
  assign _EVAL_472 = _EVAL_867 & _EVAL_1074;
  assign _EVAL_289 = _EVAL_1043 & _EVAL_1603;
  assign _EVAL_845 = _EVAL_605 ? _EVAL_1086 : _EVAL_1997;
  assign _EVAL_342 = _EVAL_936 ? _EVAL_1086 : _EVAL_1972;
  assign _EVAL_1035 = _EVAL_434 & _EVAL_1086;
  assign _EVAL_601 = _EVAL_1516 & _EVAL_1603;
  assign _EVAL_1327 = _EVAL_1096 == 2'h1;
  assign _EVAL_1113 = _EVAL_1140 & _EVAL_89;
  assign _EVAL_1742 = _EVAL_306 | _EVAL_1718;
  assign _EVAL_92 = _EVAL_712 & _EVAL_494;
  assign _EVAL_1549 = _EVAL_1030 | _EVAL_510;
  assign _EVAL_607 = _EVAL_724 & _EVAL_494;
  assign _EVAL_1020 = _EVAL_586[38];
  assign _EVAL_1950 = _EVAL_211 & _EVAL_1603;
  assign _EVAL_961 = _EVAL_423 & _EVAL_1522;
  assign _EVAL_1906 = _EVAL_391 & _EVAL_223;
  assign _EVAL_1869 = _EVAL_1605 & _EVAL_486;
  assign _EVAL_1054 = _EVAL_1322 | _EVAL_1710;
  assign _EVAL_801 = _EVAL_229 & _EVAL_854;
  assign _EVAL_344 = _EVAL_567 | _EVAL_1805;
  assign _EVAL_155 = _EVAL_1946 ? _EVAL_591 : 1024'h0;
  assign _EVAL_1127 = _EVAL_1173 ? _EVAL_331 : 1'h1;
  assign _EVAL_1837 = _EVAL_425 & _EVAL_116;
  assign _EVAL_1850 = _EVAL_1380 & _EVAL_854;
  assign _EVAL_1253 = _EVAL_922[0];
  assign _EVAL_79 = _EVAL_1681 ? _EVAL_1329 : _EVAL_915;
  assign _EVAL_1302 = _EVAL_898 & _EVAL_1603;
  assign _EVAL_161 = _EVAL_505 & _EVAL_1603;
  assign _EVAL_890 = _EVAL_1333[208];
  assign _EVAL_940 = _EVAL_2046 ? 8'hff : 8'h0;
  assign _EVAL_507 = _EVAL_1629 | _EVAL_1984;
  assign _EVAL_1721 = _EVAL_1505 & _EVAL_1603;
  assign _EVAL_1107 = ~_EVAL_967;
  assign _EVAL_1463 = _EVAL_1605 & _EVAL_1917;
  assign _EVAL_1043 = _EVAL_286 & _EVAL_1971;
  assign _EVAL_363 = &_EVAL_1775;
  assign _EVAL_936 = 6'h2e == _EVAL_1978;
  assign _EVAL_334 = _EVAL_1729 & _EVAL_1224;
  assign _EVAL_675 = ~_EVAL_1659;
  assign _EVAL_2034 = _EVAL_1532 & _EVAL_1603;
  assign _EVAL_1178 = _EVAL_426 & _EVAL_1603;
  assign _EVAL_1403 = _EVAL_1325 & _EVAL_1529;
  assign _EVAL_1865 = _EVAL_502 | _EVAL_1184;
  assign _EVAL_449 = _EVAL_1333[210];
  assign _EVAL_1346 = _EVAL_1201 & _EVAL_48;
  assign _EVAL_1358 = {_EVAL_1226,_EVAL_1905,_EVAL_1970,_EVAL_451};
  assign _EVAL_1260 = _EVAL_1681 ? _EVAL_1086 : _EVAL_64;
  assign _EVAL_1080 = _EVAL_763 & _EVAL_1603;
  assign _EVAL_150 = _EVAL_586[41];
  assign _EVAL_1359 = _EVAL_867 & _EVAL_1773;
  assign _EVAL_2031 = _EVAL_425 & _EVAL_1971;
  assign _EVAL_1744 = _EVAL_1256 & _EVAL_1001;
  assign _EVAL_2044 = _EVAL_725 & _EVAL_1603;
  assign _EVAL_1601 = _EVAL_718 ? _EVAL_1086 : _EVAL_1050;
  assign _EVAL_47 = sb2tlOpt__EVAL_16;
  assign _EVAL_1007 = ~_EVAL_566;
  assign _EVAL_1334 = 9'h10e == _EVAL_351;
  assign _EVAL_248 = _EVAL_1641 & _EVAL_223;
  assign _EVAL_286 = _EVAL_1530 & _EVAL_1086;
  assign _EVAL_1329 = {_EVAL_1274,_EVAL_1482,_EVAL_1312,_EVAL_744};
  assign _EVAL_1634 = _EVAL_1416[12];
  assign _EVAL_1125 = _EVAL_1837 | _EVAL_1160;
  assign _EVAL_253 = _EVAL_981 ? 8'hff : 8'h0;
  assign _EVAL_114 = _EVAL_557 & _EVAL_1086;
  assign _EVAL_772 = _EVAL_1505 | _EVAL_479;
  assign _EVAL_522 = _EVAL_237 & _EVAL_177;
  assign _EVAL_445 = _EVAL_1388 ? 32'hff0000f : _EVAL_546;
  assign _EVAL_1779 = _EVAL_1140 & _EVAL_264;
  assign _EVAL_46 = _EVAL_1886;
  assign _EVAL_1881 = _EVAL_1845 | _EVAL_1057;
  assign _EVAL_1442 = _EVAL_1022 & _EVAL_1603;
  assign _EVAL_1677 = _EVAL_1140 & _EVAL_444;
  assign _EVAL_1489 = _EVAL_1355 | _EVAL_1347;
  assign _EVAL_1024 = _EVAL_901[0];
  assign _EVAL_1070 = _EVAL_90 & _EVAL_1773;
  assign _EVAL_87 = {1'h0,6'h0,_EVAL_1541,_EVAL_388};
  assign _EVAL_667 = _EVAL_1801 & _EVAL_1282;
  assign _EVAL_96 = _EVAL_190 & _EVAL_1666;
  assign _EVAL_24 = _EVAL_51;
  assign _EVAL_1923 = _EVAL_400 & _EVAL_1104;
  assign _EVAL_1242 = _EVAL_625 & _EVAL_1107;
  assign _EVAL_1126 = _EVAL_819 | _EVAL_118;
  assign _EVAL_386 = _EVAL_287 & _EVAL_1773;
  assign _EVAL_1014 = _EVAL_408 | _EVAL_1283;
  assign _EVAL_701 = _EVAL_1177[23:16];
  assign _EVAL_21 = _EVAL_49;
  assign _EVAL_765 = _EVAL_1815[31:24];
  assign _EVAL_1339 = _EVAL_655[4:0];
  assign _EVAL_235 = _EVAL_191 & _EVAL_959;
  assign _EVAL_481 = ~_EVAL_1353;
  assign _EVAL_1261 = _EVAL_1042 ? _EVAL_1694 : _EVAL_1223;
  assign _EVAL_1414 = {_EVAL_448,_EVAL_1520,_EVAL_1273,_EVAL_1230};
  assign _EVAL_1079 = 9'hd9 == _EVAL_351;
  assign _EVAL_1698 = _EVAL_908 | _EVAL_504;
  assign _EVAL_1833 = _EVAL_556 & _EVAL_128;
  assign _EVAL_1933 = _EVAL_1325 & _EVAL_1020;
  assign _EVAL_321 = _EVAL_1957 & _EVAL_1603;
  assign _EVAL_63 = _EVAL_690 & _EVAL_1522;
  assign _EVAL_725 = _EVAL_286 & _EVAL_116;
  assign _EVAL_1284 = _EVAL_1141 ? _EVAL_1705 : _EVAL_436;
  assign _EVAL_702 = _EVAL_400 & _EVAL_788;
  assign _EVAL_1659 = _EVAL_1156 == 8'h0;
  assign _EVAL_7 = sb2tlOpt__EVAL_3;
  assign _EVAL_1315 = _EVAL_691 | _EVAL_572;
  assign _EVAL_560 = _EVAL_39[15:8];
  assign _EVAL_302 = _EVAL_1516 | _EVAL_125;
  assign _EVAL_589 = _EVAL_1908 | _EVAL_1210;
  assign _EVAL_486 = &_EVAL_1002;
  assign _EVAL_1058 = _EVAL_861 | _EVAL_2035;
  assign _EVAL_108 = _EVAL_1906 | _EVAL_1245;
  assign _EVAL_1421 = 9'h107 == _EVAL_351;
  assign _EVAL_444 = _EVAL_586[35];
  assign _EVAL_1203 = _EVAL_413 & _EVAL_1773;
  assign _EVAL_1087 = ~_EVAL_1541;
  assign _EVAL_200 = _EVAL_1565 & 7'h40;
  assign _EVAL_852 = 9'h111 == _EVAL_351;
  assign _EVAL_1813 = _EVAL_885 | _EVAL_1638;
  assign _EVAL_785 = 9'h100 == _EVAL_351;
  assign _EVAL_416 = _EVAL_586[24];
  assign _EVAL_1710 = _EVAL_772 & _EVAL_284;
  assign _EVAL_173 = _EVAL_1263 ? 32'h0 : _EVAL_794;
  assign _EVAL_1156 = _EVAL_756[31:24];
  assign _EVAL_636 = _EVAL_1140 & _EVAL_1529;
  assign _EVAL_710 = _EVAL_1227 | _EVAL_154;
  assign _EVAL_1756 = _EVAL_400 & _EVAL_317;
  assign _EVAL_526 = _EVAL_986 | _EVAL_1914;
  assign _EVAL_241 = _EVAL_1929 ? _EVAL_959 : _EVAL_482;
  assign _EVAL_1633 = _EVAL_1140 & _EVAL_1164;
  assign _EVAL_408 = _EVAL_1698 | _EVAL_847;
  assign _EVAL_1857 = _EVAL_410 | _EVAL_1036;
  assign _EVAL_5 = sb2tlOpt__EVAL_10;
  assign _EVAL_999 = {_EVAL_1008,_EVAL_529,_EVAL_903,_EVAL_696};
  assign _EVAL_128 = _EVAL_604[2];
  assign _EVAL_1355 = _EVAL_498 & sb2tlOpt__EVAL_0;
  assign _EVAL_769 = _EVAL_837 & _EVAL_1603;
  assign _EVAL_942 = _EVAL_389 | _EVAL_1278;
  assign _EVAL_71 = _EVAL_1125 & _EVAL_1735;
  assign _EVAL_471 = _EVAL_1996 & _EVAL_1603;
  assign _EVAL_1180 = _EVAL_1502[23:16];
  assign _EVAL_415 = _EVAL_1889 ? 32'h380006f : _EVAL_1966;
  assign _EVAL_139 = _EVAL_360 ? _EVAL_403 : _EVAL_299;
  assign _EVAL_634 = _EVAL_39[23:16];
  assign _EVAL_570 = _EVAL_1112 & _EVAL_519;
  assign _EVAL_1758 = _EVAL_740 ? _EVAL_1086 : _EVAL_1601;
  assign _EVAL_1987 = _EVAL_1502[15];
  assign _EVAL_1072 = _EVAL_1534 | _EVAL_726;
  assign _EVAL_1565 = _EVAL_42[8:2];
  assign _EVAL_1022 = _EVAL_450 & _EVAL_116;
  assign _EVAL_503 = _EVAL_43[1];
  assign _EVAL_1146 = 9'hd5 == _EVAL_351;
  assign _EVAL_56 = _EVAL_1803 ? 32'h10002623 : _EVAL_1895;
  assign _EVAL_1025 = _EVAL_135 | _EVAL_1280;
  assign _EVAL_1841 = _EVAL_1285 == 3'h1;
  assign _EVAL_1311 = _EVAL_345 & _EVAL_1928;
  assign _EVAL_239 = _EVAL_1580 & _EVAL_1824;
  assign _EVAL_1335 = &_EVAL_1422;
  assign _EVAL_1644 = _EVAL_536 ? _EVAL_1358 : _EVAL_1284;
  assign _EVAL_748 = 9'h110 == _EVAL_351;
  assign _EVAL_1091 = _EVAL_1927 & _EVAL_1086;
  assign _EVAL_13 = _EVAL_642 ? _EVAL_1544 : 32'h0;
  assign _EVAL_517 = _EVAL_204 ? _EVAL_999 : _EVAL_1689;
  assign _EVAL_1694 = {_EVAL_325,_EVAL_158,_EVAL_520,_EVAL_1318};
  assign _EVAL_1267 = _EVAL_1035 & _EVAL_854;
  assign _EVAL_1972 = _EVAL_382 ? _EVAL_1086 : _EVAL_968;
  assign _EVAL_1271 = _EVAL_996 & _EVAL_223;
  assign _EVAL_1834 = _EVAL_290 & _EVAL_854;
  assign _EVAL_2050 = _EVAL_1450 != 3'h0;
  assign _EVAL_1543 = _EVAL_1149 ? 2'h0 : _EVAL_1096;
  assign hartIsInResetSync_0_debug_hartReset_0__EVAL_2 = _EVAL_35;
  assign _EVAL_1606 = _EVAL_1590 == 3'h2;
  assign _EVAL_543 = _EVAL_1763 | _EVAL_976;
  assign _EVAL_137 = _EVAL_586[43];
  assign _EVAL_500 = _EVAL_1102 ? _EVAL_959 : _EVAL_1053;
  assign _EVAL_1507 = _EVAL_1572 | _EVAL_1910;
  assign _EVAL_460 = _EVAL_709 & _EVAL_177;
  assign _EVAL_121 = {_EVAL_1454,_EVAL_1438,_EVAL_1907,_EVAL_704};
  assign _EVAL_1574 = _EVAL_859 | _EVAL_1615;
  assign _EVAL_661 = _EVAL_1140 & _EVAL_2009;
  assign _EVAL_1388 = 9'h103 == _EVAL_351;
  assign _EVAL_819 = _EVAL_1571 | _EVAL_1574;
  assign _EVAL_1529 = _EVAL_586[39];
  assign _EVAL_1222 = _EVAL_519 ? 2'h0 : _EVAL_1543;
  assign _EVAL_899 = _EVAL_1325 & _EVAL_1164;
  assign _EVAL_1556 = _EVAL_2025[18];
  assign _EVAL_1992 = _EVAL_1256 & _EVAL_854;
  assign _EVAL_680 = _EVAL_1338 | _EVAL_597;
  assign _EVAL_838 = _EVAL_1381 | _EVAL_705;
  assign _EVAL_68 = _EVAL_1502[31:24];
  assign _EVAL_89 = _EVAL_586[40];
  assign _EVAL_1530 = _EVAL_1140 & _EVAL_1020;
  assign _EVAL_508 = _EVAL_427 | _EVAL_1613;
  assign _EVAL_446 = _EVAL_155[0];
  assign _EVAL_957 = _EVAL_1140 & _EVAL_658;
  assign _EVAL_552 = _EVAL_1333[219];
  assign _EVAL_528 = 9'h106 == _EVAL_351;
  assign _EVAL_1386 = _EVAL_1994 | _EVAL_838;
  assign _EVAL_168 = _EVAL_380 & _EVAL_959;
  assign _EVAL_348 = _EVAL_927 | _EVAL_559;
  assign _EVAL_1361 = _EVAL_1502[15:8];
  assign _EVAL_1646 = _EVAL_1035 & _EVAL_494;
  assign _EVAL_1669 = _EVAL_1365 & _EVAL_768;
  assign _EVAL_1618 = _EVAL_1140 & _EVAL_1964;
  assign _EVAL_83 = _EVAL_248 | _EVAL_1047;
  assign _EVAL_779 = _EVAL_1317 | _EVAL_1850;
  assign _EVAL_1428 = _EVAL_1742 | _EVAL_716;
  assign _EVAL_1056 = _EVAL_523 & _EVAL_1603;
  assign _EVAL_1501 = {7'h1c,_EVAL_1339,5'h0,_EVAL_1590,5'h0,7'h23};
  assign _EVAL_90 = _EVAL_897 & _EVAL_959;
  assign _EVAL_341 = _EVAL_534 & _EVAL_743;
  assign _EVAL_1969 = _EVAL_939[5];
  assign _EVAL_740 = 6'h18 == _EVAL_1978;
  assign _EVAL_456 = _EVAL_716 & _EVAL_1181;
  assign _EVAL_1757 = _EVAL_1717 & _EVAL_1971;
  assign _EVAL_994 = _EVAL_567 & _EVAL_1603;
  assign _EVAL_411 = _EVAL_939[6];
  assign _EVAL_788 = _EVAL_1333[217];
  assign _EVAL_1613 = _EVAL_1843 & _EVAL_1001;
  assign _EVAL_267 = _EVAL_389 & _EVAL_1603;
  assign _EVAL_577 = _EVAL_1843 & _EVAL_1522;
  assign _EVAL_1792 = _EVAL_1515 & _EVAL_1928;
  assign _EVAL_273 = _EVAL_1325 & _EVAL_187;
  assign _EVAL_1381 = _EVAL_626 & _EVAL_116;
  assign _EVAL_1637 = _EVAL_39[16];
  assign _EVAL_747 = _EVAL_1605 & _EVAL_412;
  assign _EVAL_2030 = _EVAL_966 ? 8'hff : 8'h0;
  assign _EVAL_1219 = _EVAL_1435 & _EVAL_959;
  assign _EVAL_1731 = _EVAL_1888 & _EVAL_1773;
  assign _EVAL_476 = {_EVAL_458,_EVAL_1844,_EVAL_735,_EVAL_1151};
  assign _EVAL_1910 = _EVAL_838 & _EVAL_1652;
  assign _EVAL_967 = _EVAL_39[10:8];
  assign _EVAL_882 = _EVAL_470 | _EVAL_352;
  assign _EVAL_1451 = _EVAL_1071 & _EVAL_1086;
  assign _EVAL_353 = _EVAL_1025 & _EVAL_1253;
  assign sb2tlOpt__EVAL_2 = _EVAL_15;
  assign _EVAL_1769 = _EVAL_921 | _EVAL_202;
  assign _EVAL_1642 = _EVAL_1565[5];
  assign _EVAL_1129 = _EVAL_90 & _EVAL_1928;
  assign _EVAL_266 = _EVAL_2025[16];
  assign _EVAL_609 = _EVAL_421 & _EVAL_1282;
  assign _EVAL_641 = _EVAL_400 & _EVAL_1568;
  assign _EVAL_159 = _EVAL_57 | _EVAL_928;
  assign _EVAL_1590 = _EVAL_2025[22:20];
  assign _EVAL_768 = sb2tlOpt__EVAL_18 != 3'h0;
  assign _EVAL_655 = _EVAL_1712 & 16'h1f;
  assign _EVAL_1980 = _EVAL_2049 ? 8'hff : 8'h0;
  assign _EVAL_924 = _EVAL_1333[216];
  assign _EVAL_1801 = _EVAL_1881 & _EVAL_865;
  assign _EVAL_1728 = _EVAL_939[7];
  assign _EVAL_1363 = _EVAL_1683 & _EVAL_1603;
  assign _EVAL_1604 = _EVAL_2031 & _EVAL_1603;
  assign _EVAL_126 = _EVAL_1897 | _EVAL_1546;
  assign _EVAL_391 = _EVAL_1092 & _EVAL_1086;
  assign _EVAL_346 = _EVAL_90 & _EVAL_177;
  assign _EVAL_122 = _EVAL_114 & _EVAL_1522;
  assign _EVAL_1716 = _EVAL_1815[15:8];
  assign _EVAL_10 = sb2tlOpt__EVAL_7;
  assign _EVAL_687 = _EVAL_867 & _EVAL_1928;
  assign _EVAL_1144 = _EVAL_1730 ? _EVAL_39 : 32'h0;
  assign _EVAL_1936 = _EVAL_586[4];
  assign _EVAL_295 = {64'h0,32'h0,_EVAL_1009};
  assign _EVAL_815 = _EVAL_40[15:8];
  assign _EVAL_1894 = _EVAL_1297 ? _EVAL_1086 : _EVAL_628;
  assign _EVAL_729 = _EVAL_1513 & _EVAL_1946;
  assign _EVAL_2051 = _EVAL_96 ? 1'h0 : _EVAL_388;
  assign _EVAL_1685 = _EVAL_1976 | _EVAL_1315;
  assign _EVAL_1552 = _EVAL_2001 & _EVAL_223;
  assign _EVAL_1176 = _EVAL_561 | _EVAL_92;
  assign _EVAL_1445 = _EVAL_521 & _EVAL_1074;
  assign _EVAL_849 = _EVAL_182 & _EVAL_1074;
  assign _EVAL_1815 = {_EVAL_651,_EVAL_940,_EVAL_253,_EVAL_2030};
  assign _EVAL_1636 = _EVAL_40[23:16];
  assign _EVAL_1735 = _EVAL_1416[14];
  assign _EVAL_1162 = _EVAL_1285 > 3'h4;
  assign _EVAL_392 = _EVAL_975 | _EVAL_1991;
  assign _EVAL_332 = _EVAL_1173 & _EVAL_1743;
  assign _EVAL_1001 = |_EVAL_1180;
  assign _EVAL_1432 = _EVAL_1096 != 2'h0;
  assign _EVAL_1867 = _EVAL_1379 & _EVAL_1603;
  assign _EVAL_1663 = _EVAL_639 | _EVAL_858;
  assign _EVAL_1092 = _EVAL_1140 & _EVAL_1962;
  assign _EVAL_828 = _EVAL_1504 ? 32'hf1402473 : _EVAL_428;
  assign _EVAL_1994 = _EVAL_170 | _EVAL_1089;
  assign _EVAL_1524 = _EVAL_1542 | _EVAL_1480;
  assign _EVAL_700 = _EVAL_785 ? 32'hc0006f : _EVAL_415;
  assign _EVAL_614 = _EVAL_168 & _EVAL_1773;
  assign _EVAL_857 = _EVAL_939[0];
  assign _EVAL_1396 = _EVAL_1091 & _EVAL_494;
  assign _EVAL_1353 = _EVAL_11 == 10'h0;
  assign _EVAL_454 = _EVAL_247 & _EVAL_1522;
  assign _EVAL_861 = _EVAL_240 & _EVAL_1971;
  assign _EVAL_1914 = _EVAL_2003 | _EVAL_98;
  assign _EVAL_1148 = _EVAL_271 & _EVAL_116;
  assign _EVAL_1232 = 6'h3c == _EVAL_1978;
  assign _EVAL_1215 = _EVAL_1061 & _EVAL_1603;
  assign _EVAL_234 = _EVAL_1325 & _EVAL_1962;
  assign _EVAL_540 = _EVAL_1468 ? _EVAL_403 : _EVAL_971;
  assign _EVAL_2036 = 6'h39 == _EVAL_1978;
  assign _EVAL_1542 = _EVAL_1730 & _EVAL_768;
  assign _EVAL_1610 = _EVAL_1685 | _EVAL_783;
  assign _EVAL_1752 = _EVAL_400 & _EVAL_951;
  assign _EVAL_23 = sb2tlOpt__EVAL_6;
  assign _EVAL_1116 = _EVAL_707 & _EVAL_1603;
  assign _EVAL_1251 = _EVAL_361 ? _EVAL_862 : _EVAL_252;
  assign _EVAL_1858 = _EVAL_237 & _EVAL_1773;
  assign _EVAL_1620 = _EVAL_1038 & _EVAL_1603;
  assign _EVAL_1010 = _EVAL_1327 & _EVAL_467;
  assign _EVAL_784 = _EVAL_423 & _EVAL_1001;
  assign _EVAL_1884 = _EVAL_1752 & _EVAL_959;
  assign _EVAL_1958 = _EVAL_1843 & _EVAL_854;
  assign _EVAL_1737 = _EVAL_901[1:0];
  assign _EVAL_1356 = _EVAL_1707 & _EVAL_1603;
  always @(posedge _EVAL_30) begin
    if (_EVAL_1109) begin
      _EVAL_158 <= 8'h0;
    end else if (_EVAL_1411) begin
      _EVAL_158 <= _EVAL_1636;
    end else if (_EVAL_935) begin
      if (_EVAL_859) begin
        _EVAL_158 <= _EVAL_634;
      end
    end
    if (_EVAL_2015) begin
      if (_EVAL_1556) begin
        _EVAL_199 <= 32'h13;
      end else begin
        _EVAL_199 <= 32'h100073;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_225 <= 1'h0;
    end else if (_EVAL_1956) begin
      _EVAL_225 <= _EVAL_1921;
    end else begin
      _EVAL_225 <= _EVAL_473;
    end
    if (_EVAL_1109) begin
      _EVAL_274 <= 1'h0;
    end else if (_EVAL_1869) begin
      _EVAL_274 <= _EVAL_327;
    end
    if (_EVAL_1109) begin
      _EVAL_308 <= 8'h0;
    end else if (_EVAL_849) begin
      _EVAL_308 <= _EVAL_1636;
    end else if (_EVAL_1116) begin
      if (_EVAL_707) begin
        _EVAL_308 <= _EVAL_634;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_325 <= 8'h0;
    end else if (_EVAL_623) begin
      _EVAL_325 <= _EVAL_1877;
    end else if (_EVAL_471) begin
      if (_EVAL_1996) begin
        _EVAL_325 <= _EVAL_178;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_333 <= 8'h0;
    end else if (_EVAL_386) begin
      _EVAL_333 <= _EVAL_1420;
    end else if (_EVAL_2044) begin
      if (_EVAL_725) begin
        _EVAL_333 <= _EVAL_1715;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_372 <= 8'h0;
    end else if (_EVAL_1185) begin
      _EVAL_372 <= _EVAL_815;
    end else if (_EVAL_316) begin
      if (_EVAL_1255) begin
        _EVAL_372 <= _EVAL_560;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_379 <= 8'h0;
    end else if (_EVAL_497) begin
      _EVAL_379 <= _EVAL_1877;
    end else if (_EVAL_1241) begin
      if (_EVAL_984) begin
        _EVAL_379 <= _EVAL_178;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_385 <= _EVAL_768;
    end
    if (_EVAL_1109) begin
      _EVAL_388 <= 1'h0;
    end else begin
      _EVAL_388 <= _EVAL_1861;
    end
    if (_EVAL_1109) begin
      _EVAL_397 <= 8'h0;
    end else if (_EVAL_1207) begin
      _EVAL_397 <= _EVAL_1636;
    end else if (_EVAL_335) begin
      if (_EVAL_1726) begin
        _EVAL_397 <= _EVAL_634;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_448 <= 8'h0;
    end else if (_EVAL_341) begin
      _EVAL_448 <= _EVAL_383;
    end else if (sb2tlOpt__EVAL_21) begin
      _EVAL_448 <= sb2tlOpt__EVAL_8;
    end
    if (_EVAL_1109) begin
      _EVAL_451 <= 8'h0;
    end else if (_EVAL_511) begin
      _EVAL_451 <= _EVAL_1420;
    end else if (_EVAL_215) begin
      if (_EVAL_1763) begin
        _EVAL_451 <= _EVAL_1715;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_458 <= 8'h0;
    end else if (_EVAL_1099) begin
      _EVAL_458 <= _EVAL_1877;
    end else if (_EVAL_1941) begin
      if (_EVAL_1757) begin
        _EVAL_458 <= _EVAL_178;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_506 <= 8'h0;
    end else if (_EVAL_1859) begin
      _EVAL_506 <= _EVAL_1877;
    end else if (_EVAL_289) begin
      if (_EVAL_1043) begin
        _EVAL_506 <= _EVAL_178;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_520 <= 8'h0;
    end else if (_EVAL_1364) begin
      _EVAL_520 <= _EVAL_815;
    end else if (_EVAL_304) begin
      if (_EVAL_1552) begin
        _EVAL_520 <= _EVAL_560;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_529 <= 8'h0;
    end else if (_EVAL_1475) begin
      _EVAL_529 <= _EVAL_1636;
    end else if (_EVAL_322) begin
      if (_EVAL_438) begin
        _EVAL_529 <= _EVAL_634;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_545 <= 8'h0;
    end else if (_EVAL_491) begin
      _EVAL_545 <= _EVAL_815;
    end else if (_EVAL_1867) begin
      if (_EVAL_1379) begin
        _EVAL_545 <= _EVAL_560;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_553 <= 8'h0;
    end else if (_EVAL_1359) begin
      _EVAL_553 <= _EVAL_1420;
    end else if (_EVAL_886) begin
      if (_EVAL_1338) begin
        _EVAL_553 <= _EVAL_1715;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_566 <= 1'h0;
    end else begin
      _EVAL_566 <= _EVAL_1587;
    end
    if (_EVAL_1109) begin
      _EVAL_578 <= 8'h0;
    end else if (_EVAL_1367) begin
      _EVAL_578 <= _EVAL_1420;
    end else if (_EVAL_1586) begin
      if (_EVAL_1381) begin
        _EVAL_578 <= _EVAL_1715;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_606 <= 8'h0;
    end else if (_EVAL_823) begin
      _EVAL_606 <= _EVAL_1420;
    end else if (_EVAL_1721) begin
      if (_EVAL_1505) begin
        _EVAL_606 <= _EVAL_1715;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_624 <= 8'h0;
    end else if (_EVAL_1129) begin
      _EVAL_624 <= _EVAL_815;
    end else if (_EVAL_2011) begin
      if (_EVAL_2003) begin
        _EVAL_624 <= _EVAL_560;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_625 <= 3'h0;
    end else if (_EVAL_297) begin
      _EVAL_625 <= 3'h1;
    end else if (_EVAL_805) begin
      _EVAL_625 <= 3'h3;
    end else if (_EVAL_1257) begin
      _EVAL_625 <= 3'h2;
    end else begin
      _EVAL_625 <= _EVAL_992;
    end
    if (_EVAL_1109) begin
      _EVAL_647 <= 1'h0;
    end else if (_EVAL_1948) begin
      _EVAL_647 <= 1'h0;
    end else if (_EVAL_159) begin
      _EVAL_647 <= 1'h0;
    end else begin
      _EVAL_647 <= _EVAL_1019;
    end
    if (_EVAL_1109) begin
      _EVAL_664 <= 8'h0;
    end else if (_EVAL_1731) begin
      _EVAL_664 <= _EVAL_1420;
    end else if (_EVAL_133) begin
      if (_EVAL_766) begin
        _EVAL_664 <= _EVAL_1715;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_684 <= 8'h0;
    end else if (_EVAL_460) begin
      _EVAL_684 <= _EVAL_1877;
    end else if (_EVAL_850) begin
      if (_EVAL_1026) begin
        _EVAL_684 <= _EVAL_178;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_692 <= 1'h0;
    end else if (_EVAL_1833) begin
      _EVAL_692 <= 1'h0;
    end else if (_EVAL_159) begin
      _EVAL_692 <= 1'h0;
    end else if (_EVAL_1629) begin
      _EVAL_692 <= 1'h0;
    end else begin
      _EVAL_692 <= _EVAL_1233;
    end
    if (_EVAL_1109) begin
      _EVAL_696 <= 8'h0;
    end else if (_EVAL_614) begin
      _EVAL_696 <= _EVAL_1420;
    end else if (_EVAL_535) begin
      if (_EVAL_561) begin
        _EVAL_696 <= _EVAL_1715;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_704 <= 8'h0;
    end else if (_EVAL_1247) begin
      _EVAL_704 <= _EVAL_1420;
    end else if (_EVAL_1075) begin
      if (_EVAL_1837) begin
        _EVAL_704 <= _EVAL_1715;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_713 <= 8'h0;
    end else if (_EVAL_1409) begin
      _EVAL_713 <= _EVAL_1636;
    end else if (_EVAL_161) begin
      if (_EVAL_505) begin
        _EVAL_713 <= _EVAL_634;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_735 <= 8'h0;
    end else if (_EVAL_1059) begin
      _EVAL_735 <= _EVAL_815;
    end else if (_EVAL_1080) begin
      if (_EVAL_763) begin
        _EVAL_735 <= _EVAL_560;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_744 <= 8'h0;
    end else if (_EVAL_1880) begin
      _EVAL_744 <= _EVAL_1420;
    end else if (_EVAL_86) begin
      if (_EVAL_831) begin
        _EVAL_744 <= _EVAL_1715;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_749 <= 8'h0;
    end else if (_EVAL_1343) begin
      _EVAL_749 <= _EVAL_1877;
    end else if (_EVAL_132) begin
      if (_EVAL_1317) begin
        _EVAL_749 <= _EVAL_178;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_754 <= 8'h0;
    end else if (_EVAL_1445) begin
      _EVAL_754 <= _EVAL_1636;
    end else if (_EVAL_420) begin
      if (_EVAL_635) begin
        _EVAL_754 <= _EVAL_634;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_777 <= 8'h0;
    end else if (_EVAL_687) begin
      _EVAL_777 <= _EVAL_815;
    end else if (_EVAL_1015) begin
      if (_EVAL_1648) begin
        _EVAL_777 <= _EVAL_560;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_822 <= 8'h0;
    end else if (_EVAL_1326) begin
      _EVAL_822 <= _EVAL_1420;
    end else if (_EVAL_1178) begin
      if (_EVAL_426) begin
        _EVAL_822 <= _EVAL_1715;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_855 <= 8'h0;
    end else if (_EVAL_270) begin
      _EVAL_855 <= _EVAL_815;
    end else if (_EVAL_1356) begin
      if (_EVAL_1707) begin
        _EVAL_855 <= _EVAL_560;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_856 <= 8'h0;
    end else if (_EVAL_2041) begin
      _EVAL_856 <= _EVAL_1877;
    end else if (_EVAL_1620) begin
      if (_EVAL_1038) begin
        _EVAL_856 <= _EVAL_178;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_903 <= 8'h0;
    end else if (_EVAL_1527) begin
      _EVAL_903 <= _EVAL_815;
    end else if (_EVAL_717) begin
      if (_EVAL_1906) begin
        _EVAL_903 <= _EVAL_560;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_922 <= 12'h0;
    end else if (_EVAL_618) begin
      _EVAL_922 <= _EVAL_1133;
    end
    if (_EVAL_1109) begin
      _EVAL_980 <= 8'h0;
    end else if (_EVAL_522) begin
      _EVAL_980 <= _EVAL_1877;
    end else if (_EVAL_1408) begin
      if (_EVAL_842) begin
        _EVAL_980 <= _EVAL_178;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_988 <= 8'h0;
    end else if (_EVAL_310) begin
      _EVAL_988 <= _EVAL_1877;
    end else if (_EVAL_2034) begin
      if (_EVAL_1532) begin
        _EVAL_988 <= _EVAL_178;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1008 <= 8'h0;
    end else if (_EVAL_1714) begin
      _EVAL_1008 <= _EVAL_1877;
    end else if (_EVAL_1488) begin
      if (_EVAL_1348) begin
        _EVAL_1008 <= _EVAL_178;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1009 <= 32'h0;
    end else if (_EVAL_609) begin
      if (_EVAL_1730) begin
        _EVAL_1009 <= _EVAL_39;
      end else begin
        _EVAL_1009 <= 32'h0;
      end
    end else if (_EVAL_1835) begin
      _EVAL_1009 <= _EVAL_757;
    end
    if (_EVAL_1109) begin
      _EVAL_1011 <= 8'h0;
    end else if (_EVAL_1858) begin
      _EVAL_1011 <= _EVAL_1420;
    end else if (_EVAL_245) begin
      if (_EVAL_135) begin
        _EVAL_1011 <= _EVAL_1715;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1048 <= 8'h0;
    end else if (_EVAL_72) begin
      _EVAL_1048 <= _EVAL_1420;
    end else if (_EVAL_321) begin
      if (_EVAL_1957) begin
        _EVAL_1048 <= _EVAL_1715;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1051 <= 8'h0;
    end else if (_EVAL_1070) begin
      _EVAL_1051 <= _EVAL_1420;
    end else if (_EVAL_1442) begin
      if (_EVAL_1022) begin
        _EVAL_1051 <= _EVAL_1715;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1063 <= 8'h0;
    end else if (_EVAL_1640) begin
      _EVAL_1063 <= _EVAL_1636;
    end else if (_EVAL_1932) begin
      if (_EVAL_1342) begin
        _EVAL_1063 <= _EVAL_634;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1096 <= 2'h0;
    end else if (_EVAL_1603) begin
      if (_EVAL_300) begin
        _EVAL_1096 <= 2'h1;
      end
    end else if (_EVAL_1327) begin
      if (_EVAL_1127) begin
        _EVAL_1096 <= 2'h0;
      end else begin
        _EVAL_1096 <= _EVAL_1793;
      end
    end else if (_EVAL_1112) begin
      _EVAL_1096 <= _EVAL_1222;
    end
    if (_EVAL_1109) begin
      _EVAL_1118 <= 8'h0;
    end else if (_EVAL_346) begin
      _EVAL_1118 <= _EVAL_1877;
    end else if (_EVAL_769) begin
      if (_EVAL_837) begin
        _EVAL_1118 <= _EVAL_178;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1151 <= 8'h0;
    end else if (_EVAL_871) begin
      _EVAL_1151 <= _EVAL_1420;
    end else if (_EVAL_715) begin
      if (_EVAL_1264) begin
        _EVAL_1151 <= _EVAL_1715;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1163 <= 8'h0;
    end else if (_EVAL_1658) begin
      _EVAL_1163 <= _EVAL_1877;
    end else if (_EVAL_989) begin
      if (_EVAL_861) begin
        _EVAL_1163 <= _EVAL_178;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1169 <= 8'h0;
    end else if (_EVAL_613) begin
      _EVAL_1169 <= _EVAL_1636;
    end else if (_EVAL_1566) begin
      if (_EVAL_888) begin
        _EVAL_1169 <= _EVAL_634;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1192 <= 8'h0;
    end else if (_EVAL_1794) begin
      _EVAL_1192 <= _EVAL_815;
    end else if (_EVAL_1056) begin
      if (_EVAL_523) begin
        _EVAL_1192 <= _EVAL_560;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1211 <= 8'h0;
    end else if (_EVAL_1203) begin
      _EVAL_1211 <= _EVAL_1420;
    end else if (_EVAL_1302) begin
      if (_EVAL_898) begin
        _EVAL_1211 <= _EVAL_1715;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1226 <= 8'h0;
    end else if (_EVAL_2043) begin
      _EVAL_1226 <= _EVAL_1877;
    end else if (_EVAL_530) begin
      if (_EVAL_84) begin
        _EVAL_1226 <= _EVAL_178;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1230 <= 8'h0;
    end else if (_EVAL_341) begin
      _EVAL_1230 <= _EVAL_640;
    end else if (sb2tlOpt__EVAL_4) begin
      _EVAL_1230 <= sb2tlOpt__EVAL_8;
    end
    if (_EVAL_1109) begin
      _EVAL_1273 <= 8'h0;
    end else if (_EVAL_341) begin
      _EVAL_1273 <= _EVAL_1000;
    end else if (sb2tlOpt__EVAL_23) begin
      _EVAL_1273 <= sb2tlOpt__EVAL_8;
    end
    if (_EVAL_1109) begin
      _EVAL_1274 <= 8'h0;
    end else if (_EVAL_337) begin
      _EVAL_1274 <= _EVAL_1877;
    end else if (_EVAL_887) begin
      if (_EVAL_825) begin
        _EVAL_1274 <= _EVAL_178;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1285 <= 3'h2;
    end else if (_EVAL_1431) begin
      _EVAL_1285 <= _EVAL_129;
    end
    if (_EVAL_1109) begin
      _EVAL_1304 <= 1'h0;
    end else if (_EVAL_747) begin
      _EVAL_1304 <= _EVAL_649;
    end
    if (_EVAL_1109) begin
      _EVAL_1305 <= 1'h0;
    end else if (_EVAL_592) begin
      _EVAL_1305 <= _EVAL_1637;
    end
    if (_EVAL_1109) begin
      _EVAL_1312 <= 8'h0;
    end else if (_EVAL_1331) begin
      _EVAL_1312 <= _EVAL_815;
    end else if (_EVAL_669) begin
      if (_EVAL_1534) begin
        _EVAL_1312 <= _EVAL_560;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1318 <= 8'h0;
    end else if (_EVAL_629) begin
      _EVAL_1318 <= _EVAL_1420;
    end else if (_EVAL_1588) begin
      if (_EVAL_1227) begin
        _EVAL_1318 <= _EVAL_1715;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1347 <= 1'h0;
    end else if (_EVAL_844) begin
      _EVAL_1347 <= 1'h0;
    end else begin
      _EVAL_1347 <= _EVAL_595;
    end
    if (_EVAL_14) begin
      _EVAL_1374 <= 1'h0;
    end else if (_EVAL_1109) begin
      _EVAL_1374 <= 1'h0;
    end else if (_EVAL_1201) begin
      _EVAL_1374 <= _EVAL_53;
    end
    if (_EVAL_1109) begin
      _EVAL_1384 <= 8'h0;
    end else if (_EVAL_1539) begin
      _EVAL_1384 <= _EVAL_1877;
    end else if (_EVAL_1783) begin
      if (_EVAL_648) begin
        _EVAL_1384 <= _EVAL_178;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1416 <= 16'h0;
    end else if (_EVAL_1418) begin
      _EVAL_1416 <= _EVAL_1136;
    end
    if (_EVAL_1109) begin
      _EVAL_1438 <= 8'h0;
    end else if (_EVAL_1852) begin
      _EVAL_1438 <= _EVAL_1636;
    end else if (_EVAL_1519) begin
      if (_EVAL_1448) begin
        _EVAL_1438 <= _EVAL_634;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1454 <= 8'h0;
    end else if (_EVAL_2047) begin
      _EVAL_1454 <= _EVAL_1877;
    end else if (_EVAL_1604) begin
      if (_EVAL_2031) begin
        _EVAL_1454 <= _EVAL_178;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1482 <= 8'h0;
    end else if (_EVAL_1791) begin
      _EVAL_1482 <= _EVAL_1636;
    end else if (_EVAL_601) begin
      if (_EVAL_1516) begin
        _EVAL_1482 <= _EVAL_634;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1483 <= 8'h0;
    end else if (_EVAL_866) begin
      _EVAL_1483 <= _EVAL_815;
    end else if (_EVAL_593) begin
      if (_EVAL_1028) begin
        _EVAL_1483 <= _EVAL_560;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1520 <= 8'h0;
    end else if (_EVAL_341) begin
      _EVAL_1520 <= _EVAL_701;
    end else if (sb2tlOpt__EVAL_13) begin
      _EVAL_1520 <= sb2tlOpt__EVAL_8;
    end
    if (_EVAL_1109) begin
      _EVAL_1541 <= 1'h0;
    end else begin
      _EVAL_1541 <= _EVAL_668;
    end
    if (_EVAL_1109) begin
      _EVAL_1616 <= 8'h0;
    end else if (_EVAL_666) begin
      _EVAL_1616 <= _EVAL_1636;
    end else if (_EVAL_1084) begin
      if (_EVAL_2033) begin
        _EVAL_1616 <= _EVAL_634;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1664 <= 8'h0;
    end else if (_EVAL_1023) begin
      _EVAL_1664 <= _EVAL_1636;
    end else if (_EVAL_994) begin
      if (_EVAL_567) begin
        _EVAL_1664 <= _EVAL_634;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1722 <= 8'h0;
    end else if (_EVAL_419) begin
      _EVAL_1722 <= _EVAL_1420;
    end else if (_EVAL_863) begin
      if (_EVAL_1148) begin
        _EVAL_1722 <= _EVAL_1715;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1723 <= 8'h0;
    end else if (_EVAL_1105) begin
      _EVAL_1723 <= _EVAL_815;
    end else if (_EVAL_244) begin
      if (_EVAL_1985) begin
        _EVAL_1723 <= _EVAL_560;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1781 <= 8'h0;
    end else if (_EVAL_107) begin
      _EVAL_1781 <= _EVAL_815;
    end else if (_EVAL_94) begin
      if (_EVAL_248) begin
        _EVAL_1781 <= _EVAL_560;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1816 <= 8'h0;
    end else if (_EVAL_472) begin
      _EVAL_1816 <= _EVAL_1636;
    end else if (_EVAL_184) begin
      if (_EVAL_643) begin
        _EVAL_1816 <= _EVAL_634;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1828 <= 8'h0;
    end else if (_EVAL_1545) begin
      _EVAL_1828 <= _EVAL_815;
    end else if (_EVAL_1804) begin
      if (_EVAL_883) begin
        _EVAL_1828 <= _EVAL_560;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1844 <= 8'h0;
    end else if (_EVAL_2017) begin
      _EVAL_1844 <= _EVAL_1636;
    end else if (_EVAL_1215) begin
      if (_EVAL_1061) begin
        _EVAL_1844 <= _EVAL_634;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1853 <= 8'h0;
    end else if (_EVAL_753) begin
      _EVAL_1853 <= _EVAL_1156;
    end
    if (_EVAL_1109) begin
      _EVAL_1882 <= 8'h0;
    end else if (_EVAL_2037) begin
      _EVAL_1882 <= _EVAL_1636;
    end else if (_EVAL_267) begin
      if (_EVAL_389) begin
        _EVAL_1882 <= _EVAL_634;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1904 <= 1'h0;
    end else if (_EVAL_600) begin
      _EVAL_1904 <= 1'h0;
    end else begin
      _EVAL_1904 <= _EVAL_1524;
    end
    if (_EVAL_1109) begin
      _EVAL_1905 <= 8'h0;
    end else if (_EVAL_1988) begin
      _EVAL_1905 <= _EVAL_1636;
    end else if (_EVAL_910) begin
      if (_EVAL_427) begin
        _EVAL_1905 <= _EVAL_634;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1907 <= 8'h0;
    end else if (_EVAL_261) begin
      _EVAL_1907 <= _EVAL_815;
    end else if (_EVAL_1307) begin
      if (_EVAL_691) begin
        _EVAL_1907 <= _EVAL_560;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1918 <= 8'h0;
    end else if (_EVAL_1311) begin
      _EVAL_1918 <= _EVAL_815;
    end else if (_EVAL_1778) begin
      if (_EVAL_1271) begin
        _EVAL_1918 <= _EVAL_560;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1922 <= 8'h0;
    end else if (_EVAL_929) begin
      _EVAL_1922 <= _EVAL_1877;
    end else if (_EVAL_1950) begin
      if (_EVAL_211) begin
        _EVAL_1922 <= _EVAL_178;
      end
    end
    if (_EVAL_2015) begin
      if (_EVAL_1900) begin
        if (_EVAL_266) begin
          _EVAL_1943 <= _EVAL_905;
        end else begin
          _EVAL_1943 <= _EVAL_1501;
        end
      end else begin
        _EVAL_1943 <= 32'h13;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1970 <= 8'h0;
    end else if (_EVAL_1792) begin
      _EVAL_1970 <= _EVAL_815;
    end else if (_EVAL_1044) begin
      if (_EVAL_1485) begin
        _EVAL_1970 <= _EVAL_560;
      end
    end
    if (_EVAL_1109) begin
      _EVAL_1989 <= 24'h0;
    end else if (_EVAL_753) begin
      _EVAL_1989 <= _EVAL_1040;
    end
    if (_EVAL_1109) begin
      _EVAL_2032 <= 8'h0;
    end else if (_EVAL_549) begin
      _EVAL_2032 <= _EVAL_1636;
    end else if (_EVAL_1363) begin
      if (_EVAL_1683) begin
        _EVAL_2032 <= _EVAL_634;
      end
    end
  end
  always @(posedge _EVAL_30 or posedge _EVAL_1885) begin
    if (_EVAL_1885) begin
      _EVAL_1886 <= 1'h0;
    end else if (_EVAL_1109) begin
      _EVAL_1886 <= 1'h0;
    end else begin
      _EVAL_1886 <= _EVAL_1866;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_158 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_199 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_225 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_274 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_308 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_325 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_333 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_372 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_379 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_385 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_388 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_397 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_448 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_451 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_458 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_506 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_520 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  _EVAL_529 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  _EVAL_545 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  _EVAL_553 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  _EVAL_566 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _EVAL_578 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  _EVAL_606 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  _EVAL_624 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  _EVAL_625 = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  _EVAL_647 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  _EVAL_664 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  _EVAL_684 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  _EVAL_692 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  _EVAL_696 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  _EVAL_704 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  _EVAL_713 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  _EVAL_735 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  _EVAL_744 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  _EVAL_749 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  _EVAL_754 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  _EVAL_777 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  _EVAL_822 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  _EVAL_855 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  _EVAL_856 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  _EVAL_903 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  _EVAL_922 = _RAND_41[11:0];
  _RAND_42 = {1{`RANDOM}};
  _EVAL_980 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  _EVAL_988 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  _EVAL_1008 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  _EVAL_1009 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  _EVAL_1011 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  _EVAL_1048 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  _EVAL_1051 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  _EVAL_1063 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  _EVAL_1096 = _RAND_50[1:0];
  _RAND_51 = {1{`RANDOM}};
  _EVAL_1118 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  _EVAL_1151 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  _EVAL_1163 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  _EVAL_1169 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  _EVAL_1192 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  _EVAL_1211 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  _EVAL_1226 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  _EVAL_1230 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  _EVAL_1273 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  _EVAL_1274 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  _EVAL_1285 = _RAND_61[2:0];
  _RAND_62 = {1{`RANDOM}};
  _EVAL_1304 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  _EVAL_1305 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  _EVAL_1312 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  _EVAL_1318 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  _EVAL_1347 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  _EVAL_1374 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  _EVAL_1384 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  _EVAL_1416 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  _EVAL_1438 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  _EVAL_1454 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  _EVAL_1482 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  _EVAL_1483 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  _EVAL_1520 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  _EVAL_1541 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  _EVAL_1616 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  _EVAL_1664 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  _EVAL_1722 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  _EVAL_1723 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  _EVAL_1781 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  _EVAL_1816 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  _EVAL_1828 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  _EVAL_1844 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  _EVAL_1853 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  _EVAL_1882 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  _EVAL_1886 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  _EVAL_1904 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  _EVAL_1905 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  _EVAL_1907 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  _EVAL_1918 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  _EVAL_1922 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  _EVAL_1943 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  _EVAL_1970 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  _EVAL_1989 = _RAND_94[23:0];
  _RAND_95 = {1{`RANDOM}};
  _EVAL_2032 = _RAND_95[7:0];
`endif // RANDOMIZE_REG_INIT
  if (_EVAL_1885) begin
    _EVAL_1886 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
