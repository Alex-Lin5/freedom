//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_163_assert(
  input        _EVAL,
  input        _EVAL_0,
  input  [1:0] _EVAL_1,
  input        _EVAL_2,
  input  [2:0] _EVAL_3,
  input        _EVAL_4,
  input  [2:0] _EVAL_5,
  input        _EVAL_6,
  input        _EVAL_7,
  input  [8:0] _EVAL_8,
  input        _EVAL_9,
  input        _EVAL_10,
  input        _EVAL_11,
  input        _EVAL_12,
  input  [1:0] _EVAL_13
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_14;
  wire  _EVAL_15;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire [8:0] _EVAL_31;
  wire  _EVAL_32;
  wire [9:0] _EVAL_33;
  wire  _EVAL_34;
  wire [1:0] _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire [9:0] _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire [9:0] _EVAL_52;
  wire  _EVAL_53;
  reg  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire [9:0] _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire [9:0] _EVAL_62;
  wire  _EVAL_63;
  wire [8:0] _EVAL_64;
  wire [9:0] _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire [8:0] _EVAL_76;
  wire  _EVAL_77;
  wire [1:0] _EVAL_78;
  wire  _EVAL_79;
  wire [9:0] _EVAL_80;
  reg [1:0] _EVAL_81;
  wire  _EVAL_83;
  wire [9:0] _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire [8:0] _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire [9:0] _EVAL_90;
  wire [9:0] _EVAL_91;
  reg  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire [31:0] _EVAL_95;
  wire  _EVAL_96;
  wire [1:0] _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire [1:0] _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  reg [2:0] _EVAL_106;
  wire  _EVAL_107;
  reg  _EVAL_108;
  wire  _EVAL_109;
  wire [9:0] _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_120;
  wire [9:0] _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  reg [8:0] _EVAL_125;
  wire  _EVAL_126;
  wire [9:0] _EVAL_127;
  wire [1:0] _EVAL_128;
  wire  _EVAL_129;
  reg  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  reg  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire [8:0] _EVAL_142;
  wire  _EVAL_143;
  reg  _EVAL_144;
  wire  _EVAL_145;
  wire [32:0] _EVAL_146;
  wire  _EVAL_147;
  wire [9:0] _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire [9:0] _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  reg [31:0] _EVAL_155;
  wire  _EVAL_156;
  wire [9:0] _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire [9:0] _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire [8:0] _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  reg  _EVAL_177;
  wire  _EVAL_178;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_182;
  reg  _EVAL_183;
  wire [1:0] _EVAL_184;
  wire  _EVAL_185;
  wire [1:0] _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  reg [1:0] _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  reg [2:0] _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire [9:0] _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_93 = ~_EVAL_129;
  assign _EVAL_169 = ~_EVAL_57;
  assign _EVAL_112 = _EVAL_0 & _EVAL_56;
  assign _EVAL_195 = _EVAL_155 < plusarg_reader_out;
  assign _EVAL_114 = ~_EVAL_150;
  assign _EVAL_149 = _EVAL_4 == _EVAL_138;
  assign _EVAL_190 = _EVAL_58 | _EVAL_143;
  assign _EVAL_18 = _EVAL_186[0];
  assign _EVAL_131 = ~_EVAL_12;
  assign _EVAL_61 = _EVAL_35[0];
  assign _EVAL_107 = _EVAL_3 == 3'h2;
  assign _EVAL_147 = _EVAL_9 & _EVAL_73;
  assign _EVAL_14 = _EVAL_5 == 3'h4;
  assign _EVAL_36 = ~_EVAL_158;
  assign _EVAL_26 = _EVAL_11 & _EVAL_9;
  assign _EVAL_59 = _EVAL_45;
  assign _EVAL_19 = _EVAL_145 | _EVAL_143;
  assign _EVAL_87 = _EVAL_8 ^ 9'h80;
  assign _EVAL_72 = plusarg_reader_out == 32'h0;
  assign _EVAL_71 = _EVAL_3 == 3'h1;
  assign _EVAL_161 = ~_EVAL_4;
  assign _EVAL_166 = _EVAL_78[0];
  assign _EVAL_48 = _EVAL_9 & _EVAL_126;
  assign _EVAL_126 = _EVAL_5 == 3'h2;
  assign _EVAL_40 = ~_EVAL_43;
  assign _EVAL_113 = _EVAL_13 == _EVAL_191;
  assign _EVAL_33 = _EVAL_121;
  assign _EVAL_85 = _EVAL_154 | _EVAL_143;
  assign _EVAL_150 = _EVAL_161 | _EVAL_143;
  assign _EVAL_179 = ~_EVAL_86;
  assign _EVAL_105 = _EVAL_60 | _EVAL_72;
  assign _EVAL_90 = {1'b0,$signed(_EVAL_76)};
  assign _EVAL_170 = _EVAL_8 ^ 9'h100;
  assign _EVAL_176 = _EVAL_118 | _EVAL_134;
  assign _EVAL_76 = _EVAL_8 ^ 9'h58;
  assign _EVAL_203 = _EVAL_184[0];
  assign _EVAL_146 = _EVAL_155 + 32'h1;
  assign _EVAL_172 = _EVAL_103[0];
  assign _EVAL_63 = _EVAL_0 & _EVAL_196;
  assign _EVAL_189 = ~_EVAL_164;
  assign _EVAL_182 = _EVAL_39 | _EVAL_132;
  assign _EVAL_184 = _EVAL_92 - 1'h1;
  assign _EVAL_21 = _EVAL_8 == _EVAL_125;
  assign _EVAL_151 = |_EVAL_183;
  assign _EVAL_157 = $signed(_EVAL_52) & -10'sh20;
  assign _EVAL_175 = ~_EVAL_183;
  assign _EVAL_160 = ~_EVAL_83;
  assign _EVAL_28 = _EVAL_17 >> _EVAL_12;
  assign _EVAL_64 = _EVAL_8 & 9'h3;
  assign _EVAL_50 = ~_EVAL_51;
  assign _EVAL_163 = _EVAL_1 == _EVAL_81;
  assign _EVAL_204 = _EVAL_24 | _EVAL_143;
  assign _EVAL_178 = ~_EVAL_190;
  assign _EVAL_62 = _EVAL_157;
  assign _EVAL_35 = _EVAL_116 ? _EVAL_128 : 2'h0;
  assign _EVAL_100 = ~_EVAL_171;
  assign _EVAL_127 = _EVAL_66;
  assign _EVAL_16 = _EVAL_123 | _EVAL_143;
  assign _EVAL_94 = _EVAL & _EVAL_0;
  assign _EVAL_115 = _EVAL_172 != _EVAL_61;
  assign _EVAL_49 = _EVAL_94 & _EVAL_79;
  assign _EVAL_84 = $signed(_EVAL_90) & -10'sh8;
  assign _EVAL_188 = _EVAL_5 == 3'h1;
  assign _EVAL_141 = _EVAL_137 | _EVAL_143;
  assign _EVAL_135 = ~_EVAL_42;
  assign _EVAL_122 = ~_EVAL_47;
  assign _EVAL_153 = ~_EVAL_19;
  assign _EVAL_45 = $signed(_EVAL_91) & -10'sh100;
  assign _EVAL_103 = _EVAL_173 ? 2'h1 : 2'h0;
  assign _EVAL_51 = _EVAL_175 | _EVAL_143;
  assign _EVAL_83 = _EVAL_3 == 3'h6;
  assign _EVAL_34 = _EVAL_149 | _EVAL_143;
  assign _EVAL_197 = ~_EVAL_85;
  assign _EVAL_38 = _EVAL_21 | _EVAL_143;
  assign _EVAL_55 = ~_EVAL_136;
  assign _EVAL_133 = ~_EVAL_168;
  assign _EVAL_198 = ~_EVAL_104;
  assign _EVAL_24 = _EVAL_88 | _EVAL_206;
  assign _EVAL_174 = _EVAL_13 >= 2'h2;
  assign _EVAL_75 = _EVAL_0 & _EVAL_107;
  assign _EVAL_164 = _EVAL_163 | _EVAL_143;
  assign _EVAL_15 = ~_EVAL_68;
  assign _EVAL_39 = $signed(_EVAL_33) == 10'sh0;
  assign _EVAL_154 = _EVAL_1 != 2'h2;
  assign _EVAL_102 = ~_EVAL_54;
  assign _EVAL_43 = _EVAL_53 | _EVAL_143;
  assign _EVAL_202 = ~_EVAL_143;
  assign _EVAL_77 = _EVAL_94 & _EVAL_136;
  assign _EVAL_22 = _EVAL_161 | _EVAL_2;
  assign _EVAL_41 = ~_EVAL_16;
  assign _EVAL_162 = _EVAL_152;
  assign _EVAL_56 = _EVAL_3 == 3'h0;
  assign _EVAL_27 = ~_EVAL_141;
  assign _EVAL_96 = $signed(_EVAL_110) == 10'sh0;
  assign _EVAL_31 = _EVAL_8 ^ 9'h60;
  assign _EVAL_99 = _EVAL_5 == 3'h3;
  assign _EVAL_29 = _EVAL_0 & _EVAL_55;
  assign _EVAL_199 = ~_EVAL_38;
  assign _EVAL_148 = {1'b0,$signed(_EVAL_142)};
  assign _EVAL_200 = {1'b0,$signed(_EVAL_8)};
  assign _EVAL_88 = _EVAL_176 | _EVAL_187;
  assign _EVAL_17 = _EVAL_172 | _EVAL_183;
  assign _EVAL_57 = _EVAL_174 | _EVAL_143;
  assign _EVAL_167 = _EVAL_12 == _EVAL_108;
  assign _EVAL_110 = _EVAL_84;
  assign _EVAL_30 = _EVAL_9 & _EVAL_15;
  assign _EVAL_23 = ~_EVAL_61;
  assign _EVAL_207 = _EVAL_183 | _EVAL_172;
  assign _EVAL_101 = ~_EVAL_98;
  assign _EVAL_205 = ~_EVAL_204;
  assign _EVAL_196 = _EVAL_3 == 3'h5;
  assign _EVAL_186 = _EVAL_54 - 1'h1;
  assign _EVAL_104 = _EVAL_131 | _EVAL_143;
  assign _EVAL_201 = _EVAL_3 == _EVAL_106;
  assign _EVAL_97 = _EVAL_177 - 1'h1;
  assign _EVAL_128 = 2'h1 << _EVAL_12;
  assign _EVAL_140 = _EVAL_64 == 9'h0;
  assign _EVAL_89 = _EVAL_0 & _EVAL_180;
  assign _EVAL_47 = _EVAL_22 | _EVAL_143;
  assign _EVAL_165 = _EVAL_97[0];
  assign _EVAL_44 = _EVAL_113 | _EVAL_143;
  assign _EVAL_42 = _EVAL_201 | _EVAL_143;
  assign _EVAL_67 = _EVAL_26 & _EVAL_68;
  assign _EVAL_37 = _EVAL_9 & _EVAL_20;
  assign _EVAL_60 = ~_EVAL_151;
  assign _EVAL_120 = _EVAL_6 == _EVAL_130;
  assign _EVAL_124 = _EVAL_0 & _EVAL_71;
  assign _EVAL_173 = _EVAL_26 & _EVAL_102;
  assign _EVAL_159 = _EVAL_9 & _EVAL_99;
  assign _EVAL_180 = _EVAL_3 == 3'h4;
  assign _EVAL_145 = _EVAL_1 == 2'h0;
  assign _EVAL_129 = _EVAL_185 | _EVAL_143;
  assign _EVAL_80 = {1'b0,$signed(_EVAL_87)};
  assign _EVAL_109 = _EVAL_9 & _EVAL_139;
  assign _EVAL_152 = $signed(_EVAL_148) & -10'shc;
  assign _EVAL_69 = _EVAL_0 & _EVAL_83;
  assign _EVAL_137 = _EVAL_3 <= 3'h6;
  assign _EVAL_142 = _EVAL_8 ^ 9'h44;
  assign _EVAL_66 = $signed(_EVAL_80) & -10'sh80;
  assign _EVAL_168 = _EVAL_120 | _EVAL_143;
  assign _EVAL_117 = _EVAL_5 == 3'h6;
  assign _EVAL_206 = $signed(_EVAL_59) == 10'sh0;
  assign _EVAL_68 = ~_EVAL_92;
  assign _EVAL_118 = _EVAL_182 | _EVAL_96;
  assign _EVAL_78 = _EVAL_144 - 1'h1;
  assign _EVAL_116 = _EVAL_49 & _EVAL_160;
  assign _EVAL_192 = _EVAL_9 & _EVAL_188;
  assign _EVAL_46 = _EVAL_26 | _EVAL_94;
  assign _EVAL_70 = ~_EVAL_44;
  assign _EVAL_91 = {1'b0,$signed(_EVAL_170)};
  assign _EVAL_95 = _EVAL_146[31:0];
  assign _EVAL_98 = _EVAL_167 | _EVAL_143;
  assign _EVAL_53 = _EVAL_5 == _EVAL_194;
  assign _EVAL_134 = $signed(_EVAL_62) == 10'sh0;
  assign _EVAL_74 = _EVAL_9 & _EVAL_14;
  assign _EVAL_58 = _EVAL_105 | _EVAL_195;
  assign _EVAL_111 = _EVAL_9 & _EVAL_117;
  assign _EVAL_32 = _EVAL_193 | _EVAL_143;
  assign _EVAL_139 = _EVAL_5 == 3'h5;
  assign _EVAL_79 = ~_EVAL_144;
  assign _EVAL_136 = ~_EVAL_177;
  assign _EVAL_121 = $signed(_EVAL_200) & -10'sh40;
  assign _EVAL_20 = _EVAL_5 == 3'h0;
  assign _EVAL_132 = $signed(_EVAL_162) == 10'sh0;
  assign _EVAL_52 = {1'b0,$signed(_EVAL_31)};
  assign _EVAL_25 = ~_EVAL_32;
  assign _EVAL_193 = _EVAL_115 | _EVAL_179;
  assign _EVAL_185 = ~_EVAL_2;
  assign _EVAL_143 = _EVAL_10;
  assign _EVAL_123 = _EVAL_1 <= 2'h2;
  assign _EVAL_86 = |_EVAL_172;
  assign _EVAL_171 = _EVAL_140 | _EVAL_143;
  assign _EVAL_73 = _EVAL_5 == 3'h7;
  assign _EVAL_158 = _EVAL_28 | _EVAL_143;
  assign _EVAL_156 = ~_EVAL_34;
  assign _EVAL_187 = $signed(_EVAL_127) == 10'sh0;
  always @(posedge _EVAL_7) begin
    if (_EVAL_77) begin
      _EVAL_81 <= _EVAL_1;
    end
    if (_EVAL_77) begin
      _EVAL_106 <= _EVAL_3;
    end
    if (_EVAL_77) begin
      _EVAL_108 <= _EVAL_12;
    end
    if (_EVAL_67) begin
      _EVAL_125 <= _EVAL_8;
    end
    if (_EVAL_77) begin
      _EVAL_130 <= _EVAL_6;
    end
    if (_EVAL_77) begin
      _EVAL_138 <= _EVAL_4;
    end
    if (_EVAL_77) begin
      _EVAL_191 <= _EVAL_13;
    end
    if (_EVAL_67) begin
      _EVAL_194 <= _EVAL_5;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c38865e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9570cb7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7ef7d83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a53c826d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa1e1a6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(559c67b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0cdc3bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9375ba8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88836edf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(773989ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87ce0fe4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e975dd5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1edd5314)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb1b2d60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(531e2c18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd066a2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d8f66a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9bdc898)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b00579c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eef5a83d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9647312e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4f4fec4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ffc180e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a2aef9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd1fe1df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c077e061)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0cdc3bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bead8409)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2494d575)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69863c14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(570b388b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9cdd086)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9adcb2b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be977c17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f78ea4aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13da3376)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(171184d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0b5465d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5674b2ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14dac17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e4447dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf8c94fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(715abdbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24804db2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f7890d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36adcb92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8057fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(450e5e9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d438878)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6d24c5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd1b7b4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6384e5c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be0abb80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3fe17d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_199) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(811cd5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e7dbe60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30 & _EVAL_199) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd5b00c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f7b2cc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(718fa646)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf237ef8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(912b307c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_202) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_202) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9c9022d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c86515bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8d9d3a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f0f9f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge _EVAL_7 or posedge _EVAL_10) begin
    if (_EVAL_10) begin
      _EVAL_54 <= 1'h0;
    end else if (_EVAL_26) begin
      if (_EVAL_102) begin
        _EVAL_54 <= 1'h0;
      end else begin
        _EVAL_54 <= _EVAL_18;
      end
    end
  end
  always @(posedge _EVAL_7 or posedge _EVAL_10) begin
    if (_EVAL_10) begin
      _EVAL_92 <= 1'h0;
    end else if (_EVAL_26) begin
      if (_EVAL_68) begin
        _EVAL_92 <= 1'h0;
      end else begin
        _EVAL_92 <= _EVAL_203;
      end
    end
  end
  always @(posedge _EVAL_7 or posedge _EVAL_10) begin
    if (_EVAL_10) begin
      _EVAL_144 <= 1'h0;
    end else if (_EVAL_94) begin
      if (_EVAL_79) begin
        _EVAL_144 <= 1'h0;
      end else begin
        _EVAL_144 <= _EVAL_166;
      end
    end
  end
  always @(posedge _EVAL_7 or posedge _EVAL_10) begin
    if (_EVAL_10) begin
      _EVAL_155 <= 32'h0;
    end else if (_EVAL_46) begin
      _EVAL_155 <= 32'h0;
    end else begin
      _EVAL_155 <= _EVAL_95;
    end
  end
  always @(posedge _EVAL_7 or posedge _EVAL_10) begin
    if (_EVAL_10) begin
      _EVAL_177 <= 1'h0;
    end else if (_EVAL_94) begin
      if (_EVAL_136) begin
        _EVAL_177 <= 1'h0;
      end else begin
        _EVAL_177 <= _EVAL_165;
      end
    end
  end
  always @(posedge _EVAL_7 or posedge _EVAL_10) begin
    if (_EVAL_10) begin
      _EVAL_183 <= 1'h0;
    end else begin
      _EVAL_183 <= _EVAL_207 & _EVAL_23;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_54 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_81 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_92 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_106 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_108 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_125 = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_130 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_138 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_144 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_155 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_177 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_183 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_191 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_194 = _RAND_13[2:0];
`endif // RANDOMIZE_REG_INIT
  if (_EVAL_10) begin
    _EVAL_54 = 1'h0;
  end
  if (_EVAL_10) begin
    _EVAL_92 = 1'h0;
  end
  if (_EVAL_10) begin
    _EVAL_144 = 1'h0;
  end
  if (_EVAL_10) begin
    _EVAL_155 = 32'h0;
  end
  if (_EVAL_10) begin
    _EVAL_177 = 1'h0;
  end
  if (_EVAL_10) begin
    _EVAL_183 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
