//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_3_assert(
  input         _EVAL,
  input  [3:0]  _EVAL_5,
  input  [3:0]  _EVAL_6,
  input  [2:0]  _EVAL_9,
  input         _EVAL_10,
  input  [2:0]  _EVAL_11,
  input  [31:0] _EVAL_16,
  input  [31:0] _EVAL_18,
  input  [3:0]  _EVAL_29,
  input         _EVAL_30,
  input         _EVAL_39,
  input  [2:0]  _EVAL_54,
  input  [2:0]  _EVAL_58,
  input         _EVAL_61,
  input         _EVAL_64,
  input  [3:0]  _EVAL_70,
  input         _EVAL_74,
  input         _EVAL_75,
  input         _EVAL_89,
  input  [3:0]  _EVAL_91,
  input         _EVAL_114,
  input         _EVAL_122,
  input         _EVAL_123,
  input  [1:0]  _EVAL_135,
  input  [2:0]  _EVAL_142,
  input         _EVAL_153,
  input         _EVAL_157,
  input         _EVAL_177,
  input         _EVAL_178,
  input         _EVAL_197,
  input         _EVAL_206,
  input         _EVAL_212,
  input         _EVAL_220,
  input  [3:0]  _EVAL_224,
  input         _EVAL_232,
  input         _EVAL_258,
  input         _EVAL_264,
  input  [2:0]  _EVAL_265,
  input         _EVAL_268,
  input  [1:0]  _EVAL_282,
  input         _EVAL_284,
  input         _EVAL_290,
  input  [3:0]  _EVAL_296,
  input         _EVAL_297,
  input         _EVAL_301,
  input         _EVAL_307,
  input  [2:0]  _EVAL_308,
  input  [4:0]  _EVAL_315,
  input  [3:0]  _EVAL_316,
  input  [4:0]  _EVAL_326,
  input         _EVAL_330,
  input         _EVAL_332,
  input         _EVAL_366,
  input         _EVAL_368,
  input  [1:0]  _EVAL_374,
  input         _EVAL_380,
  input         _EVAL_382,
  input         _EVAL_384,
  input         _EVAL_392,
  input         _EVAL_424,
  input         _EVAL_429,
  input  [3:0]  _EVAL_488,
  input         _EVAL_492,
  input  [2:0]  _EVAL_493,
  input  [1:0]  _EVAL_498,
  input         _EVAL_506
);
  wire  _EVAL_98;
  wire  _EVAL_101;
  wire  _EVAL_104;
  wire  _EVAL_108;
  wire  monitor__EVAL;
  wire  monitor__EVAL_0;
  wire [1:0] monitor__EVAL_1;
  wire [2:0] monitor__EVAL_2;
  wire  monitor__EVAL_3;
  wire  monitor__EVAL_4;
  wire [3:0] monitor__EVAL_5;
  wire [31:0] monitor__EVAL_6;
  wire [2:0] monitor__EVAL_7;
  wire  monitor__EVAL_8;
  wire  monitor__EVAL_9;
  wire [3:0] monitor__EVAL_10;
  wire  monitor__EVAL_11;
  wire [2:0] monitor__EVAL_12;
  wire  monitor__EVAL_13;
  wire  monitor__EVAL_14;
  wire  monitor__EVAL_15;
  wire  monitor__EVAL_16;
  wire [3:0] monitor__EVAL_17;
  wire  monitor__EVAL_18;
  wire  _EVAL_125;
  wire  _EVAL_129;
  wire  _EVAL_134;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_182;
  wire  _EVAL_204;
  wire  _EVAL_207;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_226;
  wire  _EVAL_228;
  wire  _EVAL_235;
  wire  _EVAL_253;
  wire  _EVAL_257;
  wire  _EVAL_261;
  wire  _EVAL_274;
  wire  _EVAL_278;
  wire  _EVAL_280;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_289;
  wire  _EVAL_293;
  wire  _EVAL_295;
  wire  _EVAL_302;
  wire  _EVAL_327;
  wire  _EVAL_328;
  wire  _EVAL_344;
  wire  _EVAL_350;
  wire  _EVAL_355;
  wire  _EVAL_360;
  wire  _EVAL_362;
  wire [31:0] monitor_1__EVAL;
  wire  monitor_1__EVAL_0;
  wire  monitor_1__EVAL_1;
  wire  monitor_1__EVAL_2;
  wire [2:0] monitor_1__EVAL_3;
  wire  monitor_1__EVAL_4;
  wire  monitor_1__EVAL_5;
  wire [3:0] monitor_1__EVAL_6;
  wire [3:0] monitor_1__EVAL_7;
  wire  monitor_1__EVAL_8;
  wire  monitor_1__EVAL_9;
  wire [3:0] monitor_1__EVAL_10;
  wire [1:0] monitor_1__EVAL_11;
  wire  monitor_1__EVAL_12;
  wire  monitor_1__EVAL_13;
  wire [3:0] monitor_1__EVAL_14;
  wire [3:0] monitor_1__EVAL_15;
  wire [2:0] monitor_1__EVAL_16;
  wire  monitor_1__EVAL_17;
  wire [2:0] monitor_1__EVAL_18;
  wire  _EVAL_387;
  wire  _EVAL_390;
  wire  _EVAL_393;
  wire  _EVAL_404;
  wire  _EVAL_410;
  wire  _EVAL_411;
  wire  _EVAL_420;
  wire  _EVAL_432;
  wire  _EVAL_442;
  wire  _EVAL_446;
  wire  _EVAL_464;
  wire  _EVAL_494;
  wire  _EVAL_495;
  wire  _EVAL_497;
  _EVAL_1_assert monitor (
    ._EVAL(monitor__EVAL),
    ._EVAL_0(monitor__EVAL_0),
    ._EVAL_1(monitor__EVAL_1),
    ._EVAL_2(monitor__EVAL_2),
    ._EVAL_3(monitor__EVAL_3),
    ._EVAL_4(monitor__EVAL_4),
    ._EVAL_5(monitor__EVAL_5),
    ._EVAL_6(monitor__EVAL_6),
    ._EVAL_7(monitor__EVAL_7),
    ._EVAL_8(monitor__EVAL_8),
    ._EVAL_9(monitor__EVAL_9),
    ._EVAL_10(monitor__EVAL_10),
    ._EVAL_11(monitor__EVAL_11),
    ._EVAL_12(monitor__EVAL_12),
    ._EVAL_13(monitor__EVAL_13),
    ._EVAL_14(monitor__EVAL_14),
    ._EVAL_15(monitor__EVAL_15),
    ._EVAL_16(monitor__EVAL_16),
    ._EVAL_17(monitor__EVAL_17),
    ._EVAL_18(monitor__EVAL_18)
  );
  _EVAL_2_assert monitor_1 (
    ._EVAL(monitor_1__EVAL),
    ._EVAL_0(monitor_1__EVAL_0),
    ._EVAL_1(monitor_1__EVAL_1),
    ._EVAL_2(monitor_1__EVAL_2),
    ._EVAL_3(monitor_1__EVAL_3),
    ._EVAL_4(monitor_1__EVAL_4),
    ._EVAL_5(monitor_1__EVAL_5),
    ._EVAL_6(monitor_1__EVAL_6),
    ._EVAL_7(monitor_1__EVAL_7),
    ._EVAL_8(monitor_1__EVAL_8),
    ._EVAL_9(monitor_1__EVAL_9),
    ._EVAL_10(monitor_1__EVAL_10),
    ._EVAL_11(monitor_1__EVAL_11),
    ._EVAL_12(monitor_1__EVAL_12),
    ._EVAL_13(monitor_1__EVAL_13),
    ._EVAL_14(monitor_1__EVAL_14),
    ._EVAL_15(monitor_1__EVAL_15),
    ._EVAL_16(monitor_1__EVAL_16),
    ._EVAL_17(monitor_1__EVAL_17),
    ._EVAL_18(monitor_1__EVAL_18)
  );
  assign monitor_1__EVAL_4 = _EVAL_258 | _EVAL_153;
  assign _EVAL_154 = ~_EVAL_290;
  assign monitor_1__EVAL = _EVAL_18;
  assign _EVAL_280 = ~_EVAL_134;
  assign _EVAL_108 = ~_EVAL_125;
  assign _EVAL_404 = ~_EVAL_264;
  assign _EVAL_350 = _EVAL_387 | _EVAL_138;
  assign monitor__EVAL_1 = _EVAL_374 | _EVAL_135;
  assign _EVAL_293 = _EVAL_228 | _EVAL_278;
  assign monitor_1__EVAL_12 = _EVAL;
  assign _EVAL_155 = _EVAL_257 | _EVAL;
  assign _EVAL_289 = ~_EVAL_506;
  assign _EVAL_104 = ~_EVAL_382;
  assign monitor__EVAL_2 = _EVAL_9;
  assign _EVAL_253 = _EVAL_344 | _EVAL;
  assign monitor__EVAL_7 = _EVAL_308 | _EVAL_493;
  assign monitor_1__EVAL_8 = _EVAL_307 | _EVAL_197;
  assign _EVAL_420 = _EVAL_212 | _EVAL_384;
  assign monitor_1__EVAL_1 = _EVAL_220 ? _EVAL_264 : _EVAL_330;
  assign _EVAL_209 = _EVAL_293 | _EVAL;
  assign monitor__EVAL_12 = _EVAL_58;
  assign monitor__EVAL_15 = _EVAL_315[0];
  assign _EVAL_432 = _EVAL_210 | _EVAL;
  assign _EVAL_129 = ~_EVAL_274;
  assign _EVAL_302 = _EVAL_387 | _EVAL_114;
  assign monitor__EVAL_8 = _EVAL;
  assign monitor_1__EVAL_15 = _EVAL_6;
  assign _EVAL_210 = _EVAL_328 | _EVAL_390;
  assign monitor_1__EVAL_14 = _EVAL_224 | _EVAL_316;
  assign _EVAL_390 = ~_EVAL_492;
  assign _EVAL_207 = _EVAL_332 | _EVAL_290;
  assign _EVAL_295 = ~_EVAL_253;
  assign _EVAL_98 = ~_EVAL_155;
  assign monitor_1__EVAL_6 = _EVAL_91;
  assign monitor__EVAL_13 = _EVAL_64;
  assign _EVAL_497 = _EVAL_355 | _EVAL_286;
  assign monitor__EVAL_11 = _EVAL_366 | _EVAL_178;
  assign _EVAL_235 = _EVAL_204 | _EVAL_154;
  assign _EVAL_226 = ~_EVAL_209;
  assign monitor_1__EVAL_16 = _EVAL_11;
  assign _EVAL_182 = ~_EVAL_432;
  assign _EVAL_360 = ~_EVAL_261;
  assign _EVAL_387 = ~_EVAL_114;
  assign monitor__EVAL_0 = _EVAL_89;
  assign _EVAL_344 = _EVAL_404 | _EVAL_264;
  assign _EVAL_261 = _EVAL_302 | _EVAL;
  assign monitor_1__EVAL_7 = _EVAL_326[3:0];
  assign _EVAL_101 = _EVAL_497 | _EVAL;
  assign _EVAL_204 = ~_EVAL_332;
  assign monitor__EVAL_16 = _EVAL_74;
  assign _EVAL_228 = ~_EVAL_232;
  assign _EVAL_278 = _EVAL_506 | _EVAL_206;
  assign monitor_1__EVAL_11 = _EVAL_498 | _EVAL_282;
  assign _EVAL_495 = ~_EVAL_411;
  assign monitor__EVAL_3 = _EVAL_61;
  assign _EVAL_411 = _EVAL_285 | _EVAL;
  assign _EVAL_125 = _EVAL_350 | _EVAL;
  assign monitor_1__EVAL_13 = _EVAL_75;
  assign _EVAL_446 = _EVAL_404 | _EVAL_207;
  assign _EVAL_286 = ~_EVAL_384;
  assign monitor_1__EVAL_9 = _EVAL_10;
  assign _EVAL_274 = _EVAL_464 | _EVAL;
  assign monitor__EVAL_14 = _EVAL_392 | _EVAL_301;
  assign _EVAL_494 = ~_EVAL_137;
  assign monitor_1__EVAL_2 = _EVAL_297 | _EVAL_268;
  assign monitor__EVAL_17 = _EVAL_70;
  assign monitor__EVAL = _EVAL_284 ? _EVAL_232 : _EVAL_429;
  assign monitor_1__EVAL_3 = _EVAL_142 | _EVAL_265;
  assign _EVAL_464 = _EVAL_289 | _EVAL_410;
  assign monitor_1__EVAL_10 = _EVAL_29;
  assign monitor__EVAL_4 = _EVAL_380 | _EVAL_123;
  assign _EVAL_355 = ~_EVAL_212;
  assign _EVAL_410 = ~_EVAL_206;
  assign _EVAL_134 = _EVAL_235 | _EVAL;
  assign monitor_1__EVAL_5 = _EVAL_39;
  assign monitor__EVAL_6 = _EVAL_16;
  assign monitor__EVAL_18 = _EVAL_157 | _EVAL_122;
  assign _EVAL_442 = ~_EVAL_101;
  assign _EVAL_138 = _EVAL_177 | _EVAL_492;
  assign _EVAL_393 = ~_EVAL_362;
  assign _EVAL_285 = _EVAL_104 | _EVAL_420;
  assign _EVAL_328 = ~_EVAL_177;
  assign monitor__EVAL_5 = _EVAL_5;
  assign _EVAL_137 = _EVAL_446 | _EVAL;
  assign _EVAL_362 = _EVAL_327 | _EVAL;
  assign monitor_1__EVAL_0 = _EVAL_424 | _EVAL_368;
  assign _EVAL_257 = _EVAL_104 | _EVAL_382;
  assign monitor_1__EVAL_18 = _EVAL_54;
  assign monitor_1__EVAL_17 = _EVAL_30;
  assign monitor__EVAL_10 = _EVAL_488 | _EVAL_296;
  assign monitor__EVAL_9 = _EVAL_10;
  assign _EVAL_327 = _EVAL_228 | _EVAL_232;
  always @(posedge _EVAL_10) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f1ee53f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2af9277)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_360) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_495) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_393) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_360) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63a93300)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f1ee53f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_393) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63a93300)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63a93300)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63a93300)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_442) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2af9277)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_494) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f1ee53f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2af9277)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2af9277)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_442) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_494) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_495) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f1ee53f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
