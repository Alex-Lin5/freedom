//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_64_assert(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  input         _EVAL_4,
  input  [4:0]  _EVAL_5,
  input  [25:0] _EVAL_6,
  input  [2:0]  _EVAL_7,
  input  [4:0]  _EVAL_8,
  input         _EVAL_9,
  input  [2:0]  _EVAL_10,
  input  [2:0]  _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  input  [3:0]  _EVAL_14
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_15;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire [25:0] _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire [17:0] _EVAL_32;
  wire  _EVAL_33;
  reg [3:0] _EVAL_34;
  reg [2:0] _EVAL_35;
  wire  _EVAL_36;
  wire [32:0] _EVAL_37;
  wire [17:0] _EVAL_38;
  reg [17:0] _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire [3:0] _EVAL_43;
  wire [3:0] _EVAL_44;
  wire [5:0] _EVAL_45;
  wire  _EVAL_46;
  wire [17:0] _EVAL_47;
  wire [3:0] _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire [3:0] _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  reg [4:0] _EVAL_61;
  wire [17:0] _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  reg [3:0] _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire [3:0] _EVAL_75;
  wire  _EVAL_76;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire [4:0] _EVAL_79;
  wire [17:0] _EVAL_80;
  wire  _EVAL_81;
  wire [12:0] _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire [2:0] _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire [12:0] _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_98;
  wire [17:0] _EVAL_99;
  wire  _EVAL_100;
  wire [31:0] _EVAL_101;
  wire  _EVAL_102;
  wire [31:0] _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire [26:0] _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire [1:0] _EVAL_117;
  wire  _EVAL_118;
  wire [5:0] _EVAL_119;
  wire [26:0] _EVAL_121;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire [4:0] _EVAL_130;
  reg [31:0] _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire [1:0] _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire [17:0] _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  reg [2:0] _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire [5:0] _EVAL_156;
  wire  _EVAL_157;
  wire [31:0] _EVAL_158;
  reg [2:0] _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  reg [2:0] _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire [3:0] _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire [17:0] _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire [5:0] _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire [3:0] _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire [2:0] _EVAL_208;
  wire  _EVAL_209;
  wire [26:0] _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire [25:0] _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire [3:0] _EVAL_221;
  wire [25:0] _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire [1:0] _EVAL_231;
  wire [4:0] _EVAL_233;
  reg [2:0] _EVAL_234;
  wire  _EVAL_235;
  wire [3:0] _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  reg [3:0] _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  reg [4:0] _EVAL_247;
  wire  _EVAL_248;
  wire [3:0] _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  reg [3:0] _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire [31:0] _EVAL_260;
  wire  _EVAL_261;
  wire [1:0] _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire [31:0] _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire [4:0] _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  reg [25:0] _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_43 = _EVAL_45[5:2];
  assign _EVAL_219 = _EVAL_229 | _EVAL_1;
  assign _EVAL_99 = _EVAL_184 & _EVAL_150;
  assign _EVAL_77 = _EVAL & _EVAL_181;
  assign _EVAL_215 = _EVAL_23 & _EVAL_72;
  assign _EVAL_125 = _EVAL_8 == 5'h10;
  assign _EVAL_174 = _EVAL_66 & _EVAL_146;
  assign _EVAL_202 = _EVAL_14 & _EVAL_44;
  assign _EVAL_145 = _EVAL_231 | 2'h1;
  assign _EVAL_147 = _EVAL_62[0];
  assign _EVAL_89 = _EVAL_145[0];
  assign _EVAL_222 = _EVAL_6 & _EVAL_22;
  assign _EVAL_138 = _EVAL_23 & _EVAL_84;
  assign _EVAL_95 = 13'h3f << _EVAL_11;
  assign _EVAL_140 = _EVAL_5 == _EVAL_61;
  assign _EVAL_263 = _EVAL_253 == 4'h0;
  assign _EVAL_230 = _EVAL & _EVAL_191;
  assign _EVAL_56 = _EVAL_202 == 4'h0;
  assign _EVAL_245 = _EVAL_252 | _EVAL_1;
  assign _EVAL_165 = _EVAL_10 <= 3'h2;
  assign _EVAL_18 = _EVAL_137 | _EVAL_174;
  assign _EVAL_107 = $signed(_EVAL_210) & -27'sh10000;
  assign _EVAL_132 = _EVAL_3 == _EVAL_173;
  assign _EVAL_129 = ~_EVAL_186;
  assign _EVAL_65 = _EVAL_4 & _EVAL_118;
  assign _EVAL_226 = _EVAL_224 | _EVAL_1;
  assign _EVAL_22 = {{20'd0}, _EVAL_45};
  assign _EVAL_47 = _EVAL_39 >> _EVAL_5;
  assign _EVAL_118 = _EVAL_7 == 3'h4;
  assign _EVAL_149 = _EVAL_155 | _EVAL_1;
  assign _EVAL_36 = _EVAL_85 <= 3'h6;
  assign _EVAL_46 = _EVAL_146 & _EVAL_72;
  assign _EVAL_206 = _EVAL_111 | _EVAL_171;
  assign _EVAL_175 = _EVAL_131 < plusarg_reader_out;
  assign _EVAL_229 = _EVAL_8 == _EVAL_247;
  assign _EVAL_203 = _EVAL_7 == 3'h2;
  assign _EVAL_198 = _EVAL_91 | _EVAL_139;
  assign _EVAL_258 = _EVAL_117 == 2'h0;
  assign _EVAL_268 = ~_EVAL_114;
  assign _EVAL_170 = _EVAL_3 == 3'h2;
  assign _EVAL_63 = _EVAL_212 | _EVAL_59;
  assign _EVAL_40 = 3'h6 == _EVAL_11;
  assign _EVAL_167 = _EVAL_180 | _EVAL_175;
  assign _EVAL_50 = _EVAL_201 | _EVAL_26;
  assign _EVAL_19 = _EVAL_161 | _EVAL_102;
  assign _EVAL_52 = _EVAL_0 & _EVAL;
  assign _EVAL_200 = _EVAL_52 | _EVAL_33;
  assign _EVAL_117 = _EVAL_8[4:3];
  assign _EVAL_259 = ~_EVAL_176;
  assign _EVAL_207 = _EVAL_24 | _EVAL_1;
  assign _EVAL_221 = _EVAL_270[3:0];
  assign _EVAL_109 = _EVAL & _EVAL_259;
  assign _EVAL_169 = ~_EVAL_219;
  assign _EVAL_112 = _EVAL_12 >= 3'h2;
  assign _EVAL_135 = _EVAL_111 & _EVAL_237;
  assign _EVAL_237 = _EVAL_127 & _EVAL_193;
  assign _EVAL_62 = _EVAL_80 >> _EVAL_8;
  assign _EVAL_157 = ~_EVAL_235;
  assign _EVAL_66 = _EVAL_145[1];
  assign _EVAL_261 = ~_EVAL_207;
  assign _EVAL_193 = $signed(_EVAL_121) == 27'sh0;
  assign _EVAL_189 = ~_EVAL_271;
  assign _EVAL_270 = _EVAL_253 - 4'h1;
  assign _EVAL_128 = _EVAL_167 | _EVAL_1;
  assign _EVAL_103 = _EVAL_124 ? _EVAL_158 : 32'h0;
  assign _EVAL_186 = _EVAL_214 | _EVAL_1;
  assign _EVAL_242 = _EVAL & _EVAL_243;
  assign _EVAL_262 = _EVAL_5[4:3];
  assign _EVAL_209 = _EVAL_197 | _EVAL_1;
  assign _EVAL_233 = _EVAL_34 - 4'h1;
  assign _EVAL_166 = _EVAL_161 | _EVAL_76;
  assign _EVAL_30 = _EVAL_134 | _EVAL_1;
  assign _EVAL_177 = _EVAL_3 == 3'h7;
  assign _EVAL_81 = ~_EVAL_136;
  assign _EVAL_181 = _EVAL_3 == 3'h5;
  assign _EVAL_228 = _EVAL_258 & _EVAL_246;
  assign _EVAL_216 = _EVAL_7 == 3'h6;
  assign _EVAL_213 = ~_EVAL_209;
  assign _EVAL_224 = _EVAL_7 <= 3'h6;
  assign _EVAL_53 = _EVAL_3 == 3'h3;
  assign _EVAL_199 = _EVAL_7 == 3'h1;
  assign _EVAL_96 = _EVAL_204 & _EVAL_166;
  assign _EVAL_269 = ~_EVAL_78;
  assign _EVAL_121 = _EVAL_107;
  assign _EVAL_69 = _EVAL & _EVAL_172;
  assign _EVAL_141 = _EVAL & _EVAL_42;
  assign _EVAL_208 = _EVAL_8[2:0];
  assign _EVAL_83 = _EVAL_146 & _EVAL_84;
  assign _EVAL_17 = ~_EVAL_149;
  assign _EVAL_156 = ~_EVAL_192;
  assign _EVAL_250 = _EVAL_6 == _EVAL_273;
  assign _EVAL_191 = _EVAL_3 == 3'h0;
  assign _EVAL_146 = ~_EVAL_23;
  assign _EVAL_88 = ~_EVAL_216;
  assign _EVAL_266 = 32'h1 << _EVAL_5;
  assign _EVAL_27 = _EVAL_89 & _EVAL_46;
  assign _EVAL_42 = _EVAL_3 == 3'h4;
  assign _EVAL_58 = ~_EVAL_14;
  assign _EVAL_86 = _EVAL_211 | _EVAL_1;
  assign _EVAL_244 = |_EVAL_39;
  assign _EVAL_92 = _EVAL_4 & _EVAL_49;
  assign _EVAL_158 = 32'h1 << _EVAL_8;
  assign _EVAL_133 = _EVAL_132 | _EVAL_1;
  assign _EVAL_110 = _EVAL_33 & _EVAL_263;
  assign _EVAL_79 = _EVAL_67 - 4'h1;
  assign _EVAL_74 = ~_EVAL_179;
  assign _EVAL_243 = _EVAL_3 == 3'h6;
  assign _EVAL_20 = ~_EVAL_226;
  assign _EVAL_41 = ~_EVAL_70;
  assign _EVAL_85 = _EVAL_5[2:0];
  assign _EVAL_154 = _EVAL_4 & _EVAL_216;
  assign _EVAL_155 = _EVAL_58 == 4'h0;
  assign _EVAL_144 = ~_EVAL_240;
  assign _EVAL_227 = _EVAL & _EVAL_53;
  assign _EVAL_91 = _EVAL_19 | _EVAL_76;
  assign _EVAL_235 = _EVAL_274 | _EVAL_1;
  assign _EVAL_94 = _EVAL_206 | _EVAL_1;
  assign _EVAL_267 = plusarg_reader_out == 32'h0;
  assign _EVAL_45 = ~_EVAL_119;
  assign _EVAL_105 = _EVAL_4 & _EVAL_203;
  assign _EVAL_33 = _EVAL_2 & _EVAL_4;
  assign _EVAL_236 = _EVAL_130[3:0];
  assign _EVAL_251 = _EVAL_112 | _EVAL_1;
  assign _EVAL_187 = _EVAL_164 | _EVAL_1;
  assign _EVAL_205 = ~_EVAL_183;
  assign _EVAL_28 = ~_EVAL_128;
  assign _EVAL_276 = _EVAL_93 | _EVAL_1;
  assign _EVAL_80 = _EVAL_38 | _EVAL_39;
  assign _EVAL_32 = _EVAL_103[17:0];
  assign _EVAL_76 = _EVAL_196 & _EVAL_36;
  assign _EVAL_15 = _EVAL_7[0];
  assign _EVAL_126 = _EVAL_7 == 3'h0;
  assign _EVAL_249 = {_EVAL_50,_EVAL_152,_EVAL_223,_EVAL_106};
  assign _EVAL_171 = _EVAL_40 & _EVAL_139;
  assign _EVAL_255 = _EVAL_8 == 5'h11;
  assign _EVAL_123 = ~_EVAL_245;
  assign _EVAL_168 = _EVAL_89 & _EVAL_138;
  assign _EVAL_93 = _EVAL_222 == 26'h0;
  assign _EVAL_21 = _EVAL & _EVAL_177;
  assign _EVAL_220 = ~_EVAL_73;
  assign _EVAL_190 = ~_EVAL_1;
  assign _EVAL_260 = _EVAL_71 ? _EVAL_266 : 32'h0;
  assign _EVAL_44 = ~_EVAL_249;
  assign _EVAL_114 = _EVAL_16 | _EVAL_1;
  assign _EVAL_192 = _EVAL_82[5:0];
  assign _EVAL_223 = _EVAL_18 | _EVAL_27;
  assign _EVAL_23 = _EVAL_6[1];
  assign _EVAL_160 = ~_EVAL_257;
  assign _EVAL_106 = _EVAL_18 | _EVAL_98;
  assign _EVAL_254 = _EVAL_14 == _EVAL_249;
  assign _EVAL_124 = _EVAL_110 & _EVAL_88;
  assign _EVAL_264 = _EVAL_165 | _EVAL_1;
  assign _EVAL_274 = ~_EVAL_13;
  assign _EVAL_150 = ~_EVAL_32;
  assign _EVAL_143 = _EVAL_52 & _EVAL_176;
  assign _EVAL_60 = ~_EVAL_115;
  assign _EVAL_102 = _EVAL_5 == 5'h10;
  assign _EVAL_134 = _EVAL_10 == _EVAL_159;
  assign _EVAL_163 = _EVAL_113 | _EVAL_1;
  assign _EVAL_275 = _EVAL_250 | _EVAL_1;
  assign _EVAL_164 = _EVAL_12 == _EVAL_234;
  assign _EVAL_90 = _EVAL_66 & _EVAL_23;
  assign _EVAL_210 = {1'b0,$signed(_EVAL_218)};
  assign _EVAL_139 = _EVAL_5 == 5'h8;
  assign _EVAL_179 = _EVAL_135 | _EVAL_1;
  assign _EVAL_73 = _EVAL_63 | _EVAL_1;
  assign _EVAL_265 = _EVAL & _EVAL_170;
  assign _EVAL_57 = ~_EVAL_30;
  assign _EVAL_197 = ~_EVAL_31;
  assign _EVAL_101 = _EVAL_37[31:0];
  assign _EVAL_38 = _EVAL_260[17:0];
  assign _EVAL_212 = _EVAL_241 | _EVAL_228;
  assign _EVAL_68 = _EVAL_4 & _EVAL_126;
  assign _EVAL_218 = _EVAL_6 ^ 26'h2000000;
  assign _EVAL_178 = _EVAL_233[3:0];
  assign _EVAL_271 = _EVAL_137 | _EVAL_1;
  assign _EVAL_82 = 13'h3f << _EVAL_12;
  assign _EVAL_115 = _EVAL_3[2];
  assign _EVAL_201 = _EVAL_137 | _EVAL_90;
  assign _EVAL_176 = _EVAL_34 == 4'h0;
  assign _EVAL_59 = _EVAL_8 == 5'h8;
  assign _EVAL_29 = _EVAL_10 <= 3'h4;
  assign _EVAL_148 = ~_EVAL_86;
  assign _EVAL_214 = _EVAL_10 <= 3'h1;
  assign _EVAL_136 = _EVAL_198 | _EVAL_1;
  assign _EVAL_51 = _EVAL_4 & _EVAL_199;
  assign _EVAL_257 = _EVAL_239 == 4'h0;
  assign _EVAL_185 = _EVAL_4 & _EVAL_160;
  assign _EVAL_71 = _EVAL_52 & _EVAL_87;
  assign _EVAL_100 = _EVAL_147 | _EVAL_1;
  assign _EVAL_151 = ~_EVAL_94;
  assign _EVAL_277 = ~_EVAL_133;
  assign _EVAL_98 = _EVAL_89 & _EVAL_83;
  assign _EVAL_64 = ~_EVAL_187;
  assign _EVAL_78 = _EVAL_140 | _EVAL_1;
  assign _EVAL_16 = _EVAL_11 == _EVAL_153;
  assign _EVAL_49 = _EVAL_7 == 3'h5;
  assign _EVAL_75 = _EVAL_79[3:0];
  assign _EVAL_87 = _EVAL_67 == 4'h0;
  assign _EVAL_182 = ~_EVAL_251;
  assign _EVAL_127 = _EVAL_11 <= 3'h6;
  assign _EVAL_217 = _EVAL_237 | _EVAL_1;
  assign _EVAL_231 = 2'h1 << _EVAL_238;
  assign _EVAL_240 = _EVAL_29 | _EVAL_1;
  assign _EVAL_72 = _EVAL_6[0];
  assign _EVAL_48 = _EVAL_156[5:2];
  assign _EVAL_252 = _EVAL_7 == _EVAL_35;
  assign _EVAL_180 = _EVAL_108 | _EVAL_267;
  assign _EVAL_70 = _EVAL_56 | _EVAL_1;
  assign _EVAL_24 = _EVAL_10 != 3'h0;
  assign _EVAL_195 = ~_EVAL_276;
  assign _EVAL_272 = ~_EVAL_275;
  assign _EVAL_183 = _EVAL_254 | _EVAL_1;
  assign _EVAL_184 = _EVAL_39 | _EVAL_38;
  assign _EVAL_104 = ~_EVAL_163;
  assign _EVAL_108 = ~_EVAL_244;
  assign _EVAL_26 = _EVAL_89 & _EVAL_215;
  assign _EVAL_113 = _EVAL_10 == 3'h0;
  assign _EVAL_248 = ~_EVAL_264;
  assign _EVAL_31 = _EVAL_47[0];
  assign _EVAL_196 = _EVAL_262 == 2'h0;
  assign _EVAL_111 = _EVAL_96 | _EVAL_102;
  assign _EVAL_119 = _EVAL_95[5:0];
  assign _EVAL_225 = ~_EVAL_100;
  assign _EVAL_137 = _EVAL_11 >= 3'h2;
  assign _EVAL_238 = _EVAL_11[0];
  assign _EVAL_152 = _EVAL_201 | _EVAL_168;
  assign _EVAL_204 = _EVAL_11 <= 3'h2;
  assign _EVAL_130 = _EVAL_239 - 4'h1;
  assign _EVAL_84 = ~_EVAL_72;
  assign _EVAL_162 = ~_EVAL_217;
  assign _EVAL_211 = _EVAL_10 <= 3'h3;
  assign _EVAL_241 = _EVAL_255 | _EVAL_125;
  assign _EVAL_246 = _EVAL_208 <= 3'h6;
  assign _EVAL_161 = _EVAL_5 == 5'h11;
  assign _EVAL_55 = _EVAL_33 & _EVAL_257;
  assign _EVAL_37 = _EVAL_131 + 32'h1;
  assign _EVAL_172 = _EVAL_3 == 3'h1;
  always @(posedge _EVAL_9) begin
    if (_EVAL_1) begin
      _EVAL_34 <= 4'h0;
    end else if (_EVAL_52) begin
      if (_EVAL_176) begin
        if (_EVAL_60) begin
          _EVAL_34 <= _EVAL_43;
        end else begin
          _EVAL_34 <= 4'h0;
        end
      end else begin
        _EVAL_34 <= _EVAL_178;
      end
    end
    if (_EVAL_55) begin
      _EVAL_35 <= _EVAL_7;
    end
    if (_EVAL_1) begin
      _EVAL_39 <= 18'h0;
    end else begin
      _EVAL_39 <= _EVAL_99;
    end
    if (_EVAL_143) begin
      _EVAL_61 <= _EVAL_5;
    end
    if (_EVAL_1) begin
      _EVAL_67 <= 4'h0;
    end else if (_EVAL_52) begin
      if (_EVAL_87) begin
        if (_EVAL_60) begin
          _EVAL_67 <= _EVAL_43;
        end else begin
          _EVAL_67 <= 4'h0;
        end
      end else begin
        _EVAL_67 <= _EVAL_75;
      end
    end
    if (_EVAL_1) begin
      _EVAL_131 <= 32'h0;
    end else if (_EVAL_200) begin
      _EVAL_131 <= 32'h0;
    end else begin
      _EVAL_131 <= _EVAL_101;
    end
    if (_EVAL_143) begin
      _EVAL_153 <= _EVAL_11;
    end
    if (_EVAL_143) begin
      _EVAL_159 <= _EVAL_10;
    end
    if (_EVAL_143) begin
      _EVAL_173 <= _EVAL_3;
    end
    if (_EVAL_55) begin
      _EVAL_234 <= _EVAL_12;
    end
    if (_EVAL_1) begin
      _EVAL_239 <= 4'h0;
    end else if (_EVAL_33) begin
      if (_EVAL_257) begin
        if (_EVAL_15) begin
          _EVAL_239 <= _EVAL_48;
        end else begin
          _EVAL_239 <= 4'h0;
        end
      end else begin
        _EVAL_239 <= _EVAL_236;
      end
    end
    if (_EVAL_55) begin
      _EVAL_247 <= _EVAL_8;
    end
    if (_EVAL_1) begin
      _EVAL_253 <= 4'h0;
    end else if (_EVAL_33) begin
      if (_EVAL_263) begin
        if (_EVAL_15) begin
          _EVAL_253 <= _EVAL_48;
        end else begin
          _EVAL_253 <= 4'h0;
        end
      end else begin
        _EVAL_253 <= _EVAL_221;
      end
    end
    if (_EVAL_143) begin
      _EVAL_273 <= _EVAL_6;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42f2bc7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a22e055)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4b66a32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb2751f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1f45e4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87a66b89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a622491)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e2e36cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ae8153b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(513d442f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c85f1d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37110eb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12e9f6d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(246436f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf8fb34c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ffe40c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56379e15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abf5b42c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12f05680)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3fbebc24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af69b15f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b818ebcf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef0c6e40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(209964b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(280da9ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a37d95eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf0b76fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81963bb1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec64a1fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1744f86f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(397474d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61556281)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(526a9f4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de9db57b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9380972b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94e81ddc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96800052)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ac5d25f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a2b1eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(893c3a38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a03b0f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5fee555)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58a9b896)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6f071b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5231656a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6406365a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_268) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff26968)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(983678de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d045fc75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8fa2511e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd182fd1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad0c986a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76e96602)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83d373a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d01f9aeb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(779977c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5145c636)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3002833e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28ff3480)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36daaf41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14552f13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4c694b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb56e98a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f04f3b85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(246436f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0610a10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13f57b4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa03bc39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84de2ea6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c7d03a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ae29081)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af1756a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bac927e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e3b05ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(872f6e44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_227 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_34 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_35 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_39 = _RAND_2[17:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_61 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_67 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_131 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_153 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_159 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_173 = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_234 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_239 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_247 = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_253 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_273 = _RAND_13[25:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
