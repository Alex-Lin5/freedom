//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_26_assert(
  input  [2:0]  _EVAL,
  input  [1:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input  [31:0] _EVAL_4,
  input  [3:0]  _EVAL_5,
  input  [2:0]  _EVAL_6,
  input  [2:0]  _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input  [3:0]  _EVAL_16,
  input  [3:0]  _EVAL_17,
  input         _EVAL_18
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  reg [3:0] _EVAL_26;
  reg [1:0] _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  reg  _EVAL_34;
  wire  _EVAL_35;
  wire [6:0] _EVAL_36;
  wire  _EVAL_37;
  wire [3:0] _EVAL_38;
  wire  _EVAL_39;
  wire [1:0] _EVAL_40;
  wire  _EVAL_41;
  wire [5:0] _EVAL_42;
  wire  _EVAL_43;
  wire [1:0] _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire [5:0] _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire [32:0] _EVAL_56;
  wire [1:0] _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire [1:0] _EVAL_64;
  wire [22:0] _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  reg [31:0] _EVAL_69;
  wire [6:0] _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire [32:0] _EVAL_73;
  wire  _EVAL_74;
  reg [3:0] _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire [32:0] _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire [32:0] _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire [5:0] _EVAL_92;
  wire [5:0] _EVAL_93;
  wire  _EVAL_94;
  wire [1:0] _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  reg [2:0] _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire [1:0] _EVAL_109;
  wire  _EVAL_110;
  wire [3:0] _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire [32:0] _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire [32:0] _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire [32:0] _EVAL_122;
  wire  _EVAL_123;
  wire [32:0] _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  reg [2:0] _EVAL_133;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire [7:0] _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire [31:0] _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire [1:0] _EVAL_154;
  wire  _EVAL_155;
  wire [32:0] _EVAL_156;
  wire [31:0] _EVAL_157;
  wire [1:0] _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire [32:0] _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire [31:0] _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire [7:0] _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire [31:0] _EVAL_181;
  wire [32:0] _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire [32:0] _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire [3:0] _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire [32:0] _EVAL_200;
  wire  _EVAL_201;
  wire [1:0] _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  reg [5:0] _EVAL_208;
  wire [32:0] _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  reg [1:0] _EVAL_212;
  wire  _EVAL_213;
  reg  _EVAL_214;
  wire  _EVAL_215;
  wire [31:0] _EVAL_216;
  wire [6:0] _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire [32:0] _EVAL_227;
  wire  _EVAL_228;
  wire [1:0] _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire [31:0] _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_238;
  wire [7:0] _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire [32:0] _EVAL_244;
  wire [31:0] _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  reg [31:0] _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire [32:0] _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  reg [5:0] _EVAL_257;
  wire [32:0] _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire [22:0] _EVAL_262;
  wire  _EVAL_263;
  wire [32:0] _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire [31:0] _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  reg [5:0] _EVAL_273;
  wire [32:0] _EVAL_274;
  wire [1:0] _EVAL_275;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  reg [5:0] _EVAL_282;
  wire [32:0] _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire [32:0] _EVAL_287;
  wire  _EVAL_288;
  reg  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire [32:0] _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_294;
  wire  _EVAL_295;
  wire  _EVAL_296;
  wire  _EVAL_297;
  wire [5:0] _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_307;
  reg [2:0] _EVAL_308;
  reg  _EVAL_309;
  wire  _EVAL_310;
  wire  _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_317;
  wire  _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_320;
  wire [1:0] _EVAL_321;
  wire [32:0] _EVAL_322;
  wire  _EVAL_323;
  wire  _EVAL_324;
  wire [6:0] _EVAL_325;
  wire  _EVAL_326;
  wire [31:0] _EVAL_327;
  wire  _EVAL_328;
  wire  _EVAL_329;
  wire [7:0] _EVAL_330;
  wire [32:0] _EVAL_332;
  wire  _EVAL_333;
  wire  _EVAL_334;
  wire  _EVAL_335;
  wire  _EVAL_336;
  wire  _EVAL_337;
  wire  _EVAL_338;
  wire  _EVAL_339;
  wire [31:0] _EVAL_340;
  wire  _EVAL_341;
  wire  _EVAL_342;
  wire  _EVAL_343;
  wire  _EVAL_344;
  wire [5:0] _EVAL_345;
  wire [3:0] _EVAL_346;
  wire  _EVAL_347;
  wire  _EVAL_348;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_127 = ~_EVAL_300;
  assign _EVAL_228 = ~_EVAL_341;
  assign _EVAL_170 = _EVAL_314 | _EVAL_10;
  assign _EVAL_217 = _EVAL_208 - 6'h1;
  assign _EVAL_203 = ~_EVAL_41;
  assign _EVAL_261 = ~_EVAL_198;
  assign _EVAL_70 = _EVAL_257 - 6'h1;
  assign _EVAL_196 = ~_EVAL_39;
  assign _EVAL_306 = _EVAL_166 | _EVAL_10;
  assign _EVAL_179 = ~_EVAL_170;
  assign _EVAL_177 = _EVAL_262[7:0];
  assign _EVAL_150 = ~_EVAL_218;
  assign _EVAL_321 = 2'h1 << _EVAL_115;
  assign _EVAL_277 = _EVAL_2 & _EVAL_18;
  assign _EVAL_153 = _EVAL_259 | _EVAL_10;
  assign _EVAL_143 = _EVAL_7 != 3'h0;
  assign _EVAL_253 = $signed(_EVAL_73) & -33'sh4000;
  assign _EVAL_42 = _EVAL_239[7:2];
  assign _EVAL_148 = ~_EVAL_113;
  assign _EVAL_22 = _EVAL_311 | _EVAL_240;
  assign _EVAL_87 = _EVAL_11 == _EVAL_34;
  assign _EVAL_152 = ~_EVAL_236;
  assign _EVAL_146 = _EVAL_4 ^ 32'h40000000;
  assign _EVAL_328 = _EVAL == 3'h4;
  assign _EVAL_173 = _EVAL_4 ^ 32'h1800000;
  assign _EVAL_224 = ~_EVAL_104;
  assign _EVAL_188 = _EVAL_0 == _EVAL_27;
  assign _EVAL_58 = _EVAL_69 < plusarg_reader_out;
  assign _EVAL_259 = _EVAL_17 == _EVAL_111;
  assign _EVAL_53 = _EVAL_301 | _EVAL_10;
  assign _EVAL_239 = ~_EVAL_137;
  assign _EVAL_51 = _EVAL == 3'h0;
  assign _EVAL_132 = _EVAL_5 <= 4'h8;
  assign _EVAL_305 = ~_EVAL_334;
  assign _EVAL_154 = ~_EVAL_57;
  assign _EVAL_251 = _EVAL_43 | _EVAL_10;
  assign _EVAL_112 = _EVAL_315 | _EVAL_10;
  assign _EVAL_140 = _EVAL_280 | _EVAL_10;
  assign _EVAL_68 = _EVAL_15 & _EVAL_333;
  assign _EVAL_65 = 23'hff << _EVAL_16;
  assign _EVAL_36 = _EVAL_273 - 6'h1;
  assign _EVAL_263 = _EVAL_255 | _EVAL_277;
  assign _EVAL_44 = 2'h1 << _EVAL_12;
  assign _EVAL_145 = _EVAL_151 | _EVAL_45;
  assign _EVAL_218 = _EVAL_249 | _EVAL_10;
  assign _EVAL_303 = _EVAL_15 & _EVAL_32;
  assign _EVAL_149 = _EVAL_241 | _EVAL_72;
  assign _EVAL_115 = _EVAL_5[0];
  assign _EVAL_192 = _EVAL_253;
  assign _EVAL_320 = _EVAL_5 <= 4'hb;
  assign _EVAL_111 = {_EVAL_119,_EVAL_176,_EVAL_74,_EVAL_266};
  assign _EVAL_252 = _EVAL_347 & _EVAL_8;
  assign _EVAL_155 = _EVAL_174 | _EVAL_10;
  assign _EVAL_39 = _EVAL_4[0];
  assign _EVAL_310 = ~_EVAL_110;
  assign _EVAL_307 = _EVAL_132 & _EVAL_329;
  assign _EVAL_147 = ~_EVAL_84;
  assign _EVAL_317 = _EVAL_125 | _EVAL_10;
  assign _EVAL_118 = _EVAL_6 == 3'h7;
  assign _EVAL_231 = _EVAL_265 | _EVAL_10;
  assign _EVAL_144 = _EVAL_15 & _EVAL_118;
  assign _EVAL_334 = _EVAL_335 | _EVAL_10;
  assign _EVAL_79 = _EVAL_15 & _EVAL_296;
  assign _EVAL_73 = {1'b0,$signed(_EVAL_173)};
  assign _EVAL_258 = {1'b0,$signed(_EVAL_327)};
  assign _EVAL_195 = _EVAL_109[1];
  assign _EVAL_122 = _EVAL_69 + 32'h1;
  assign _EVAL_345 = _EVAL_325[5:0];
  assign _EVAL_91 = _EVAL_5 <= 4'h6;
  assign _EVAL_287 = $signed(_EVAL_322) & -33'sh10000;
  assign _EVAL_85 = _EVAL_12 == _EVAL_214;
  assign _EVAL_32 = _EVAL_6 == 3'h6;
  assign _EVAL_78 = _EVAL_171 | _EVAL_10;
  assign _EVAL_181 = _EVAL_4 & _EVAL_216;
  assign _EVAL_57 = _EVAL_24 ? _EVAL_44 : 2'h0;
  assign _EVAL_211 = _EVAL == _EVAL_133;
  assign _EVAL_120 = _EVAL_60 | _EVAL_10;
  assign _EVAL_201 = ~_EVAL_46;
  assign _EVAL_157 = _EVAL_4 ^ 32'hc000000;
  assign _EVAL_339 = _EVAL_145 | _EVAL_121;
  assign _EVAL_247 = ~_EVAL_306;
  assign _EVAL_243 = _EVAL_6 == 3'h3;
  assign _EVAL_46 = _EVAL_160 | _EVAL_10;
  assign _EVAL_137 = _EVAL_65[7:0];
  assign _EVAL_123 = _EVAL_7 <= 3'h3;
  assign _EVAL_255 = _EVAL_13 & _EVAL_15;
  assign _EVAL_61 = ~_EVAL_159;
  assign _EVAL_92 = _EVAL_217[5:0];
  assign _EVAL_43 = _EVAL_6 == _EVAL_308;
  assign _EVAL_104 = _EVAL_4[1];
  assign _EVAL_23 = ~_EVAL_140;
  assign _EVAL_116 = _EVAL_91 & _EVAL_260;
  assign _EVAL_299 = ~_EVAL_278;
  assign _EVAL_129 = _EVAL_0 <= 2'h2;
  assign _EVAL_98 = _EVAL_5 == _EVAL_75;
  assign _EVAL_159 = _EVAL_48 | _EVAL_10;
  assign _EVAL_119 = _EVAL_22 | _EVAL_225;
  assign _EVAL_74 = _EVAL_80 | _EVAL_77;
  assign _EVAL_241 = ~_EVAL_206;
  assign _EVAL_139 = _EVAL_109[0];
  assign _EVAL_319 = _EVAL_15 & _EVAL_164;
  assign _EVAL_298 = _EVAL_330[7:2];
  assign _EVAL_163 = _EVAL_139 & _EVAL_167;
  assign _EVAL_175 = _EVAL_91 & _EVAL_288;
  assign _EVAL_185 = ~_EVAL_66;
  assign _EVAL_190 = _EVAL_282 == 6'h0;
  assign _EVAL_174 = _EVAL_16 == _EVAL_26;
  assign _EVAL_89 = _EVAL_6 == 3'h0;
  assign _EVAL_271 = _EVAL_31 | _EVAL_10;
  assign _EVAL_76 = ~_EVAL_316;
  assign _EVAL_234 = ~_EVAL_1;
  assign _EVAL_330 = ~_EVAL_177;
  assign _EVAL_77 = _EVAL_139 & _EVAL_242;
  assign _EVAL_59 = _EVAL_255 & _EVAL_189;
  assign _EVAL_290 = ~_EVAL_153;
  assign _EVAL_340 = _EVAL_4 ^ 32'h3000;
  assign _EVAL_227 = _EVAL_274;
  assign _EVAL_62 = _EVAL_129 | _EVAL_10;
  assign _EVAL_186 = _EVAL_307 | _EVAL_55;
  assign _EVAL_107 = _EVAL_301 & _EVAL_160;
  assign _EVAL_269 = _EVAL_226 | _EVAL_10;
  assign _EVAL_301 = _EVAL_252 | _EVAL_254;
  assign _EVAL_295 = ~_EVAL_53;
  assign _EVAL_332 = _EVAL_124;
  assign _EVAL_109 = _EVAL_321 | 2'h1;
  assign _EVAL_286 = _EVAL_211 | _EVAL_10;
  assign _EVAL_278 = _EVAL_143 | _EVAL_10;
  assign _EVAL_165 = {1'b0,$signed(_EVAL_157)};
  assign _EVAL_88 = _EVAL_114;
  assign _EVAL_191 = ~_EVAL_62;
  assign _EVAL_274 = $signed(_EVAL_56) & -33'sh2000;
  assign _EVAL_347 = _EVAL_5 <= 4'h2;
  assign _EVAL_169 = ~_EVAL_112;
  assign _EVAL_96 = _EVAL_273 == 6'h0;
  assign _EVAL_229 = _EVAL_158 >> _EVAL_12;
  assign _EVAL_294 = _EVAL_15 & _EVAL_205;
  assign _EVAL_230 = ~_EVAL_12;
  assign _EVAL_156 = {1'b0,$signed(_EVAL_340)};
  assign _EVAL_124 = $signed(_EVAL_292) & -33'sh2000;
  assign _EVAL_67 = ~_EVAL_63;
  assign _EVAL_184 = _EVAL_270 | _EVAL_10;
  assign _EVAL_198 = _EVAL_186 | _EVAL_10;
  assign _EVAL_158 = _EVAL_64 | _EVAL_212;
  assign _EVAL_95 = 2'h1 << _EVAL_8;
  assign _EVAL_242 = _EVAL_224 & _EVAL_39;
  assign _EVAL_244 = $signed(_EVAL_258) & -33'sh4000;
  assign _EVAL_180 = _EVAL_104 & _EVAL_196;
  assign _EVAL_281 = ~_EVAL_219;
  assign _EVAL_279 = ~_EVAL_25;
  assign _EVAL_102 = ~_EVAL_155;
  assign _EVAL_205 = _EVAL_6 == 3'h2;
  assign _EVAL_246 = $signed(_EVAL_82) == 33'sh0;
  assign _EVAL_93 = _EVAL_70[5:0];
  assign _EVAL_216 = {{24'd0}, _EVAL_330};
  assign _EVAL_292 = {1'b0,$signed(_EVAL_245)};
  assign _EVAL_215 = _EVAL_7 == _EVAL_100;
  assign _EVAL_72 = plusarg_reader_out == 32'h0;
  assign _EVAL_66 = _EVAL_215 | _EVAL_10;
  assign _EVAL_197 = ~_EVAL_17;
  assign _EVAL_117 = _EVAL_287;
  assign _EVAL_41 = _EVAL_204 | _EVAL_10;
  assign _EVAL_225 = _EVAL_139 & _EVAL_94;
  assign _EVAL_90 = _EVAL_202[0];
  assign _EVAL_280 = _EVAL_0 != 2'h2;
  assign _EVAL_128 = _EVAL_213 | _EVAL_10;
  assign _EVAL_291 = ~_EVAL_142;
  assign _EVAL_204 = _EVAL_149 | _EVAL_58;
  assign _EVAL_136 = _EVAL_318 | _EVAL_10;
  assign _EVAL_24 = _EVAL_161 & _EVAL_310;
  assign _EVAL_220 = _EVAL_233 | _EVAL_10;
  assign _EVAL_324 = _EVAL_37 | _EVAL_10;
  assign _EVAL_240 = _EVAL_195 & _EVAL_104;
  assign _EVAL_83 = $signed(_EVAL_227) == 33'sh0;
  assign _EVAL_56 = {1'b0,$signed(_EVAL_146)};
  assign _EVAL_202 = _EVAL_212 >> _EVAL_8;
  assign _EVAL_55 = _EVAL_91 & _EVAL_248;
  assign _EVAL_342 = _EVAL_64 != _EVAL_57;
  assign _EVAL_245 = _EVAL_4 ^ 32'h20000000;
  assign _EVAL_141 = ~_EVAL_21;
  assign _EVAL_209 = _EVAL_200;
  assign _EVAL_200 = $signed(_EVAL_182) & -33'sh5000;
  assign _EVAL_126 = _EVAL_18 & _EVAL_33;
  assign _EVAL_99 = _EVAL_337 | _EVAL_348;
  assign _EVAL_19 = _EVAL_307 | _EVAL_116;
  assign _EVAL_213 = _EVAL_181 == 32'h0;
  assign _EVAL_232 = ~_EVAL_120;
  assign _EVAL_97 = _EVAL == 3'h5;
  assign _EVAL_297 = _EVAL_106 | _EVAL_10;
  assign _EVAL_142 = _EVAL_234 | _EVAL_10;
  assign _EVAL_264 = $signed(_EVAL_156) & -33'sh1000;
  assign _EVAL_322 = {1'b0,$signed(_EVAL_235)};
  assign _EVAL_37 = _EVAL_12 | _EVAL_230;
  assign _EVAL_341 = _EVAL_188 | _EVAL_10;
  assign _EVAL_131 = _EVAL_18 & _EVAL_51;
  assign _EVAL_189 = _EVAL_257 == 6'h0;
  assign _EVAL_45 = $signed(_EVAL_192) == 33'sh0;
  assign _EVAL_235 = _EVAL_4 ^ 32'h2000000;
  assign _EVAL_348 = $signed(_EVAL_332) == 33'sh0;
  assign _EVAL_108 = ~_EVAL_184;
  assign _EVAL_82 = _EVAL_244;
  assign _EVAL_130 = ~_EVAL_10;
  assign _EVAL_178 = ~_EVAL_8;
  assign _EVAL_226 = _EVAL_0 == 2'h0;
  assign _EVAL_101 = _EVAL_7 <= 3'h4;
  assign _EVAL_49 = _EVAL_99 | _EVAL_83;
  assign _EVAL_327 = _EVAL_4 ^ 32'h80000000;
  assign _EVAL_335 = _EVAL_7 <= 3'h1;
  assign _EVAL_80 = _EVAL_311 | _EVAL_29;
  assign _EVAL_25 = _EVAL_6[2];
  assign _EVAL_266 = _EVAL_80 | _EVAL_163;
  assign _EVAL_193 = ~_EVAL_128;
  assign _EVAL_166 = ~_EVAL_11;
  assign _EVAL_21 = _EVAL_311 | _EVAL_10;
  assign _EVAL_161 = _EVAL_277 & _EVAL_86;
  assign _EVAL_249 = _EVAL_342 | _EVAL_76;
  assign _EVAL_270 = ~_EVAL_90;
  assign _EVAL_105 = ~_EVAL_297;
  assign _EVAL_313 = _EVAL_18 & _EVAL_328;
  assign _EVAL_35 = ~_EVAL_231;
  assign _EVAL_338 = ~_EVAL_256;
  assign _EVAL_38 = _EVAL_17 & _EVAL_346;
  assign _EVAL_265 = _EVAL_38 == 4'h0;
  assign _EVAL_304 = ~_EVAL_96;
  assign _EVAL_47 = ~_EVAL_269;
  assign _EVAL_316 = |_EVAL_64;
  assign _EVAL_337 = _EVAL_339 | _EVAL_343;
  assign _EVAL_260 = _EVAL_337 | _EVAL_246;
  assign _EVAL_314 = _EVAL_4 == _EVAL_250;
  assign _EVAL_296 = _EVAL_6 == 3'h5;
  assign _EVAL_121 = $signed(_EVAL_117) == 33'sh0;
  assign _EVAL_50 = _EVAL_36[5:0];
  assign _EVAL_323 = _EVAL_123 | _EVAL_10;
  assign _EVAL_84 = _EVAL_107 | _EVAL_10;
  assign _EVAL_254 = _EVAL_320 & _EVAL_178;
  assign _EVAL_343 = $signed(_EVAL_88) == 33'sh0;
  assign _EVAL_29 = _EVAL_195 & _EVAL_224;
  assign _EVAL_182 = {1'b0,$signed(_EVAL_4)};
  assign _EVAL_207 = _EVAL == 3'h1;
  assign _EVAL_288 = _EVAL_49 | _EVAL_246;
  assign _EVAL_325 = _EVAL_282 - 6'h1;
  assign _EVAL_176 = _EVAL_22 | _EVAL_199;
  assign _EVAL_206 = |_EVAL_212;
  assign _EVAL_329 = $signed(_EVAL_284) == 33'sh0;
  assign _EVAL_160 = _EVAL_307 | _EVAL_175;
  assign _EVAL_293 = _EVAL_18 & _EVAL_223;
  assign _EVAL_151 = $signed(_EVAL_209) == 33'sh0;
  assign _EVAL_48 = _EVAL_7 <= 3'h2;
  assign _EVAL_248 = _EVAL_348 | _EVAL_83;
  assign _EVAL_272 = _EVAL_18 & _EVAL_110;
  assign _EVAL_210 = _EVAL_18 & _EVAL_207;
  assign _EVAL_318 = ~_EVAL_9;
  assign _EVAL_64 = _EVAL_59 ? _EVAL_95 : 2'h0;
  assign _EVAL_326 = ~_EVAL_136;
  assign _EVAL_275 = _EVAL_40 & _EVAL_154;
  assign _EVAL_194 = ~_EVAL_317;
  assign _EVAL_222 = ~_EVAL_220;
  assign _EVAL_233 = _EVAL <= 3'h6;
  assign _EVAL_54 = ~_EVAL_286;
  assign _EVAL_114 = $signed(_EVAL_165) & -33'sh400000;
  assign _EVAL_113 = _EVAL_85 | _EVAL_10;
  assign _EVAL_219 = _EVAL_98 | _EVAL_10;
  assign _EVAL_71 = _EVAL_19 | _EVAL_10;
  assign _EVAL_40 = _EVAL_212 | _EVAL_64;
  assign _EVAL_315 = _EVAL_229[0];
  assign _EVAL_106 = _EVAL_7 == 3'h0;
  assign _EVAL_125 = _EVAL_14 == _EVAL_289;
  assign _EVAL_172 = _EVAL_15 & _EVAL_243;
  assign _EVAL_168 = _EVAL_15 & _EVAL_89;
  assign _EVAL_63 = _EVAL_87 | _EVAL_10;
  assign _EVAL_94 = _EVAL_104 & _EVAL_39;
  assign _EVAL_262 = 23'hff << _EVAL_5;
  assign _EVAL_162 = _EVAL_197 == 4'h0;
  assign _EVAL_221 = _EVAL_277 & _EVAL_190;
  assign _EVAL_183 = _EVAL_255 & _EVAL_96;
  assign _EVAL_344 = _EVAL_18 & _EVAL_97;
  assign _EVAL_135 = ~_EVAL_324;
  assign _EVAL_86 = _EVAL_208 == 6'h0;
  assign _EVAL_110 = _EVAL == 3'h6;
  assign _EVAL_223 = ~_EVAL_190;
  assign _EVAL_284 = _EVAL_264;
  assign _EVAL_268 = _EVAL_122[31:0];
  assign _EVAL_285 = ~_EVAL_71;
  assign _EVAL_346 = ~_EVAL_111;
  assign _EVAL_311 = _EVAL_5 >= 4'h2;
  assign _EVAL_256 = _EVAL_101 | _EVAL_10;
  assign _EVAL_236 = _EVAL_162 | _EVAL_10;
  assign _EVAL_300 = _EVAL_138 | _EVAL_10;
  assign _EVAL_164 = _EVAL_6 == 3'h1;
  assign _EVAL_333 = _EVAL_6 == 3'h4;
  assign _EVAL_171 = _EVAL_8 == _EVAL_309;
  assign _EVAL_31 = _EVAL_16 >= 4'h2;
  assign _EVAL_302 = _EVAL_15 & _EVAL_304;
  assign _EVAL_199 = _EVAL_139 & _EVAL_180;
  assign _EVAL_138 = _EVAL_8 | _EVAL_178;
  assign _EVAL_20 = ~_EVAL_251;
  assign _EVAL_167 = _EVAL_224 & _EVAL_196;
  assign _EVAL_28 = ~_EVAL_323;
  assign _EVAL_33 = _EVAL == 3'h2;
  assign _EVAL_312 = ~_EVAL_271;
  assign _EVAL_238 = ~_EVAL_78;
  assign _EVAL_60 = _EVAL_166 | _EVAL_1;
  assign _EVAL_336 = _EVAL[0];
  always @(posedge _EVAL_3) begin
    if (_EVAL_221) begin
      _EVAL_26 <= _EVAL_16;
    end
    if (_EVAL_221) begin
      _EVAL_27 <= _EVAL_0;
    end
    if (_EVAL_221) begin
      _EVAL_34 <= _EVAL_11;
    end
    if (_EVAL_10) begin
      _EVAL_69 <= 32'h0;
    end else if (_EVAL_263) begin
      _EVAL_69 <= 32'h0;
    end else begin
      _EVAL_69 <= _EVAL_268;
    end
    if (_EVAL_183) begin
      _EVAL_75 <= _EVAL_5;
    end
    if (_EVAL_183) begin
      _EVAL_100 <= _EVAL_7;
    end
    if (_EVAL_221) begin
      _EVAL_133 <= _EVAL;
    end
    if (_EVAL_10) begin
      _EVAL_208 <= 6'h0;
    end else if (_EVAL_277) begin
      if (_EVAL_86) begin
        if (_EVAL_336) begin
          _EVAL_208 <= _EVAL_42;
        end else begin
          _EVAL_208 <= 6'h0;
        end
      end else begin
        _EVAL_208 <= _EVAL_92;
      end
    end
    if (_EVAL_10) begin
      _EVAL_212 <= 2'h0;
    end else begin
      _EVAL_212 <= _EVAL_275;
    end
    if (_EVAL_221) begin
      _EVAL_214 <= _EVAL_12;
    end
    if (_EVAL_183) begin
      _EVAL_250 <= _EVAL_4;
    end
    if (_EVAL_10) begin
      _EVAL_257 <= 6'h0;
    end else if (_EVAL_255) begin
      if (_EVAL_189) begin
        if (_EVAL_279) begin
          _EVAL_257 <= _EVAL_298;
        end else begin
          _EVAL_257 <= 6'h0;
        end
      end else begin
        _EVAL_257 <= _EVAL_93;
      end
    end
    if (_EVAL_10) begin
      _EVAL_273 <= 6'h0;
    end else if (_EVAL_255) begin
      if (_EVAL_96) begin
        if (_EVAL_279) begin
          _EVAL_273 <= _EVAL_298;
        end else begin
          _EVAL_273 <= 6'h0;
        end
      end else begin
        _EVAL_273 <= _EVAL_50;
      end
    end
    if (_EVAL_10) begin
      _EVAL_282 <= 6'h0;
    end else if (_EVAL_277) begin
      if (_EVAL_190) begin
        if (_EVAL_336) begin
          _EVAL_282 <= _EVAL_42;
        end else begin
          _EVAL_282 <= 6'h0;
        end
      end else begin
        _EVAL_282 <= _EVAL_345;
      end
    end
    if (_EVAL_221) begin
      _EVAL_289 <= _EVAL_14;
    end
    if (_EVAL_183) begin
      _EVAL_308 <= _EVAL_6;
    end
    if (_EVAL_183) begin
      _EVAL_309 <= _EVAL_8;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d09e6875)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc26eb47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_102) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5831e9b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47dfe604)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e1d5b81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5c6a36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6af4ce00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da5f4774)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8301f39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0f93bfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27caa4c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_326) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb7d5048)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db9fd575)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_326) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(995b77b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5c74cc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4bf1d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1663bfeb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb2dd8e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a542a8d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b66c1f0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f676f0ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd5625e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(495c5485)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_326) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7249881)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46fc0c0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72c9c590)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f5146e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_285) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92dc1807)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8bf2afd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65db9035)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53f926c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e06360a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df0dbbeb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8802e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78d2527d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(885b8a42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2aaff6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_299) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(191bdce6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_305) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8301f39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bb0d946)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(590c2ad4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_281) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b3702b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b5c26a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad0cafc8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6dae5fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bc96a46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_338) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(326b7cb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93db0e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(894ce389)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ddd7914)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14129d3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dff2e521)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_326) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a74f4061)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fa430b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9898805a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45c4cc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8157b586)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_326) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac5d4ec0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c23bc7f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13a37980)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a7c947a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf5d5a1c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d69e218)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d6df305)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(344ad383)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8fda8d8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_285) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53ea79e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2f88d66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f14d10c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_326) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82194cbf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5691d13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9e0dc1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de3ee9c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15e25643)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2bbf582)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb0a5ba6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_326) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ae10853)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_305) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ba5553b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_281) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(915c274c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7dff342)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bf6ef90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(794b52cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_102) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d298625)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_299) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d7ca90d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c075d5d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d78485d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_294 & _EVAL_338) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2110283)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_326) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c60bfd27)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22518968)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(988158fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_79 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_272 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9c2898e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_68 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce5f320d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73980745)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88d8b5b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_26 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_27 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_34 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_69 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_75 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_100 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_133 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_208 = _RAND_7[5:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_212 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_214 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_250 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_257 = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_273 = _RAND_12[5:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_282 = _RAND_13[5:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_289 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_308 = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_309 = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
