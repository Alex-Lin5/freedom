//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_100(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input  [3:0]  _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  output [2:0]  _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18,
  output        _EVAL_19,
  input         _EVAL_20,
  input         _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  input         _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  input         _EVAL_30,
  input  [31:0] _EVAL_31,
  input         _EVAL_32,
  input         _EVAL_33,
  input         _EVAL_34,
  input         _EVAL_35,
  input         _EVAL_36,
  input         _EVAL_37,
  input         _EVAL_38,
  input         _EVAL_39,
  input         _EVAL_40,
  input         _EVAL_41,
  input         _EVAL_42,
  input  [27:0] _EVAL_43,
  output [9:0]  _EVAL_44,
  input         _EVAL_45,
  input         _EVAL_46,
  input         _EVAL_47,
  input         _EVAL_48,
  input         _EVAL_49,
  input         _EVAL_50,
  input         _EVAL_51,
  input         _EVAL_52,
  input         _EVAL_53,
  input         _EVAL_54,
  input         _EVAL_55,
  input         _EVAL_56,
  input         _EVAL_57,
  input         _EVAL_58,
  input         _EVAL_59,
  input         _EVAL_60,
  input         _EVAL_61,
  input         _EVAL_62,
  input         _EVAL_63,
  input         _EVAL_64,
  input         _EVAL_65,
  input         _EVAL_66,
  input         _EVAL_67,
  input         _EVAL_68,
  input         _EVAL_69,
  input         _EVAL_70,
  input         _EVAL_71,
  input         _EVAL_72,
  input         _EVAL_73,
  input         _EVAL_74,
  input         _EVAL_75,
  input         _EVAL_76,
  input         _EVAL_77,
  input         _EVAL_78,
  input         _EVAL_79,
  input  [2:0]  _EVAL_80,
  input         _EVAL_81,
  input         _EVAL_82,
  input         _EVAL_83,
  input         _EVAL_84,
  input         _EVAL_85,
  input         _EVAL_86,
  input         _EVAL_87,
  input         _EVAL_88,
  input         _EVAL_89,
  input         _EVAL_90,
  input         _EVAL_91,
  input         _EVAL_92,
  input         _EVAL_93,
  input         _EVAL_94,
  input         _EVAL_95,
  input         _EVAL_96,
  input         _EVAL_97,
  input         _EVAL_98,
  input         _EVAL_99,
  input         _EVAL_100,
  input         _EVAL_101,
  input  [2:0]  _EVAL_102,
  input         _EVAL_103,
  input         _EVAL_104,
  input         _EVAL_105,
  input         _EVAL_106,
  input         _EVAL_107,
  output        _EVAL_108,
  input         _EVAL_109,
  input         _EVAL_110,
  input         _EVAL_111,
  input         _EVAL_112,
  input         _EVAL_113,
  input         _EVAL_114,
  input         _EVAL_115,
  input         _EVAL_116,
  input  [9:0]  _EVAL_117,
  input         _EVAL_118,
  input         _EVAL_119,
  input         _EVAL_120,
  input         _EVAL_121,
  input         _EVAL_122,
  input         _EVAL_123,
  input         _EVAL_124,
  input         _EVAL_125,
  output        _EVAL_126,
  input         _EVAL_127,
  output [1:0]  _EVAL_128,
  input         _EVAL_129,
  input         _EVAL_130,
  input         _EVAL_131,
  input         _EVAL_132,
  input         _EVAL_133,
  input         _EVAL_134,
  input         _EVAL_135,
  input         _EVAL_136,
  input         _EVAL_137,
  input         _EVAL_138,
  input         _EVAL_139,
  output [31:0] _EVAL_140,
  input  [1:0]  _EVAL_141,
  input         _EVAL_142,
  input         _EVAL_143,
  input         _EVAL_144
);
  wire  plic__EVAL;
  wire  plic__EVAL_0;
  wire  plic__EVAL_1;
  wire  plic__EVAL_2;
  wire  plic__EVAL_3;
  wire  plic__EVAL_4;
  wire  plic__EVAL_5;
  wire [2:0] plic__EVAL_6;
  wire  plic__EVAL_7;
  wire  plic__EVAL_8;
  wire  plic__EVAL_9;
  wire  plic__EVAL_10;
  wire  plic__EVAL_11;
  wire  plic__EVAL_12;
  wire  plic__EVAL_13;
  wire  plic__EVAL_14;
  wire  plic__EVAL_15;
  wire  plic__EVAL_16;
  wire [1:0] plic__EVAL_17;
  wire  plic__EVAL_18;
  wire  plic__EVAL_19;
  wire  plic__EVAL_20;
  wire  plic__EVAL_21;
  wire  plic__EVAL_22;
  wire  plic__EVAL_23;
  wire  plic__EVAL_24;
  wire  plic__EVAL_25;
  wire  plic__EVAL_26;
  wire  plic__EVAL_27;
  wire  plic__EVAL_28;
  wire  plic__EVAL_29;
  wire  plic__EVAL_30;
  wire  plic__EVAL_31;
  wire [2:0] plic__EVAL_32;
  wire  plic__EVAL_33;
  wire  plic__EVAL_34;
  wire  plic__EVAL_35;
  wire  plic__EVAL_36;
  wire  plic__EVAL_37;
  wire  plic__EVAL_38;
  wire  plic__EVAL_39;
  wire  plic__EVAL_40;
  wire  plic__EVAL_41;
  wire  plic__EVAL_42;
  wire  plic__EVAL_43;
  wire  plic__EVAL_44;
  wire  plic__EVAL_45;
  wire  plic__EVAL_46;
  wire  plic__EVAL_47;
  wire  plic__EVAL_48;
  wire  plic__EVAL_49;
  wire  plic__EVAL_50;
  wire  plic__EVAL_51;
  wire  plic__EVAL_52;
  wire  plic__EVAL_53;
  wire  plic__EVAL_54;
  wire  plic__EVAL_55;
  wire  plic__EVAL_56;
  wire  plic__EVAL_57;
  wire  plic__EVAL_58;
  wire  plic__EVAL_59;
  wire  plic__EVAL_60;
  wire  plic__EVAL_61;
  wire  plic__EVAL_62;
  wire  plic__EVAL_63;
  wire  plic__EVAL_64;
  wire  plic__EVAL_65;
  wire  plic__EVAL_66;
  wire  plic__EVAL_67;
  wire  plic__EVAL_68;
  wire  plic__EVAL_69;
  wire [2:0] plic__EVAL_70;
  wire  plic__EVAL_71;
  wire  plic__EVAL_72;
  wire [9:0] plic__EVAL_73;
  wire  plic__EVAL_74;
  wire  plic__EVAL_75;
  wire  plic__EVAL_76;
  wire  plic__EVAL_77;
  wire  plic__EVAL_78;
  wire  plic__EVAL_79;
  wire  plic__EVAL_80;
  wire  plic__EVAL_81;
  wire  plic__EVAL_82;
  wire  plic__EVAL_83;
  wire [3:0] plic__EVAL_84;
  wire  plic__EVAL_85;
  wire  plic__EVAL_86;
  wire  plic__EVAL_87;
  wire  plic__EVAL_88;
  wire  plic__EVAL_89;
  wire  plic__EVAL_90;
  wire  plic__EVAL_91;
  wire  plic__EVAL_92;
  wire  plic__EVAL_93;
  wire  plic__EVAL_94;
  wire  plic__EVAL_95;
  wire  plic__EVAL_96;
  wire [31:0] plic__EVAL_97;
  wire  plic__EVAL_98;
  wire  plic__EVAL_99;
  wire  plic__EVAL_100;
  wire [31:0] plic__EVAL_101;
  wire  plic__EVAL_102;
  wire  plic__EVAL_103;
  wire  plic__EVAL_104;
  wire  plic__EVAL_105;
  wire  plic__EVAL_106;
  wire  plic__EVAL_107;
  wire  plic__EVAL_108;
  wire  plic__EVAL_109;
  wire  plic__EVAL_110;
  wire  plic__EVAL_111;
  wire  plic__EVAL_112;
  wire  plic__EVAL_113;
  wire  plic__EVAL_114;
  wire  plic__EVAL_115;
  wire  plic__EVAL_116;
  wire  plic__EVAL_117;
  wire  plic__EVAL_118;
  wire  plic__EVAL_119;
  wire  plic__EVAL_120;
  wire  plic__EVAL_121;
  wire  plic__EVAL_122;
  wire  plic__EVAL_123;
  wire [9:0] plic__EVAL_124;
  wire  plic__EVAL_125;
  wire [1:0] plic__EVAL_126;
  wire  plic__EVAL_127;
  wire  plic__EVAL_128;
  wire  plic__EVAL_129;
  wire [27:0] plic__EVAL_130;
  wire  plic__EVAL_131;
  wire  plic__EVAL_132;
  wire  plic__EVAL_133;
  wire  plic__EVAL_134;
  wire  plic__EVAL_135;
  wire  plic__EVAL_136;
  wire  plic__EVAL_137;
  wire  plic__EVAL_138;
  wire  plic__EVAL_139;
  wire  plic__EVAL_140;
  wire  plic__EVAL_141;
  wire  plic__EVAL_142;
  wire  plic__EVAL_143;
  wire  plic__EVAL_144;
  _EVAL_99 plic (
    ._EVAL(plic__EVAL),
    ._EVAL_0(plic__EVAL_0),
    ._EVAL_1(plic__EVAL_1),
    ._EVAL_2(plic__EVAL_2),
    ._EVAL_3(plic__EVAL_3),
    ._EVAL_4(plic__EVAL_4),
    ._EVAL_5(plic__EVAL_5),
    ._EVAL_6(plic__EVAL_6),
    ._EVAL_7(plic__EVAL_7),
    ._EVAL_8(plic__EVAL_8),
    ._EVAL_9(plic__EVAL_9),
    ._EVAL_10(plic__EVAL_10),
    ._EVAL_11(plic__EVAL_11),
    ._EVAL_12(plic__EVAL_12),
    ._EVAL_13(plic__EVAL_13),
    ._EVAL_14(plic__EVAL_14),
    ._EVAL_15(plic__EVAL_15),
    ._EVAL_16(plic__EVAL_16),
    ._EVAL_17(plic__EVAL_17),
    ._EVAL_18(plic__EVAL_18),
    ._EVAL_19(plic__EVAL_19),
    ._EVAL_20(plic__EVAL_20),
    ._EVAL_21(plic__EVAL_21),
    ._EVAL_22(plic__EVAL_22),
    ._EVAL_23(plic__EVAL_23),
    ._EVAL_24(plic__EVAL_24),
    ._EVAL_25(plic__EVAL_25),
    ._EVAL_26(plic__EVAL_26),
    ._EVAL_27(plic__EVAL_27),
    ._EVAL_28(plic__EVAL_28),
    ._EVAL_29(plic__EVAL_29),
    ._EVAL_30(plic__EVAL_30),
    ._EVAL_31(plic__EVAL_31),
    ._EVAL_32(plic__EVAL_32),
    ._EVAL_33(plic__EVAL_33),
    ._EVAL_34(plic__EVAL_34),
    ._EVAL_35(plic__EVAL_35),
    ._EVAL_36(plic__EVAL_36),
    ._EVAL_37(plic__EVAL_37),
    ._EVAL_38(plic__EVAL_38),
    ._EVAL_39(plic__EVAL_39),
    ._EVAL_40(plic__EVAL_40),
    ._EVAL_41(plic__EVAL_41),
    ._EVAL_42(plic__EVAL_42),
    ._EVAL_43(plic__EVAL_43),
    ._EVAL_44(plic__EVAL_44),
    ._EVAL_45(plic__EVAL_45),
    ._EVAL_46(plic__EVAL_46),
    ._EVAL_47(plic__EVAL_47),
    ._EVAL_48(plic__EVAL_48),
    ._EVAL_49(plic__EVAL_49),
    ._EVAL_50(plic__EVAL_50),
    ._EVAL_51(plic__EVAL_51),
    ._EVAL_52(plic__EVAL_52),
    ._EVAL_53(plic__EVAL_53),
    ._EVAL_54(plic__EVAL_54),
    ._EVAL_55(plic__EVAL_55),
    ._EVAL_56(plic__EVAL_56),
    ._EVAL_57(plic__EVAL_57),
    ._EVAL_58(plic__EVAL_58),
    ._EVAL_59(plic__EVAL_59),
    ._EVAL_60(plic__EVAL_60),
    ._EVAL_61(plic__EVAL_61),
    ._EVAL_62(plic__EVAL_62),
    ._EVAL_63(plic__EVAL_63),
    ._EVAL_64(plic__EVAL_64),
    ._EVAL_65(plic__EVAL_65),
    ._EVAL_66(plic__EVAL_66),
    ._EVAL_67(plic__EVAL_67),
    ._EVAL_68(plic__EVAL_68),
    ._EVAL_69(plic__EVAL_69),
    ._EVAL_70(plic__EVAL_70),
    ._EVAL_71(plic__EVAL_71),
    ._EVAL_72(plic__EVAL_72),
    ._EVAL_73(plic__EVAL_73),
    ._EVAL_74(plic__EVAL_74),
    ._EVAL_75(plic__EVAL_75),
    ._EVAL_76(plic__EVAL_76),
    ._EVAL_77(plic__EVAL_77),
    ._EVAL_78(plic__EVAL_78),
    ._EVAL_79(plic__EVAL_79),
    ._EVAL_80(plic__EVAL_80),
    ._EVAL_81(plic__EVAL_81),
    ._EVAL_82(plic__EVAL_82),
    ._EVAL_83(plic__EVAL_83),
    ._EVAL_84(plic__EVAL_84),
    ._EVAL_85(plic__EVAL_85),
    ._EVAL_86(plic__EVAL_86),
    ._EVAL_87(plic__EVAL_87),
    ._EVAL_88(plic__EVAL_88),
    ._EVAL_89(plic__EVAL_89),
    ._EVAL_90(plic__EVAL_90),
    ._EVAL_91(plic__EVAL_91),
    ._EVAL_92(plic__EVAL_92),
    ._EVAL_93(plic__EVAL_93),
    ._EVAL_94(plic__EVAL_94),
    ._EVAL_95(plic__EVAL_95),
    ._EVAL_96(plic__EVAL_96),
    ._EVAL_97(plic__EVAL_97),
    ._EVAL_98(plic__EVAL_98),
    ._EVAL_99(plic__EVAL_99),
    ._EVAL_100(plic__EVAL_100),
    ._EVAL_101(plic__EVAL_101),
    ._EVAL_102(plic__EVAL_102),
    ._EVAL_103(plic__EVAL_103),
    ._EVAL_104(plic__EVAL_104),
    ._EVAL_105(plic__EVAL_105),
    ._EVAL_106(plic__EVAL_106),
    ._EVAL_107(plic__EVAL_107),
    ._EVAL_108(plic__EVAL_108),
    ._EVAL_109(plic__EVAL_109),
    ._EVAL_110(plic__EVAL_110),
    ._EVAL_111(plic__EVAL_111),
    ._EVAL_112(plic__EVAL_112),
    ._EVAL_113(plic__EVAL_113),
    ._EVAL_114(plic__EVAL_114),
    ._EVAL_115(plic__EVAL_115),
    ._EVAL_116(plic__EVAL_116),
    ._EVAL_117(plic__EVAL_117),
    ._EVAL_118(plic__EVAL_118),
    ._EVAL_119(plic__EVAL_119),
    ._EVAL_120(plic__EVAL_120),
    ._EVAL_121(plic__EVAL_121),
    ._EVAL_122(plic__EVAL_122),
    ._EVAL_123(plic__EVAL_123),
    ._EVAL_124(plic__EVAL_124),
    ._EVAL_125(plic__EVAL_125),
    ._EVAL_126(plic__EVAL_126),
    ._EVAL_127(plic__EVAL_127),
    ._EVAL_128(plic__EVAL_128),
    ._EVAL_129(plic__EVAL_129),
    ._EVAL_130(plic__EVAL_130),
    ._EVAL_131(plic__EVAL_131),
    ._EVAL_132(plic__EVAL_132),
    ._EVAL_133(plic__EVAL_133),
    ._EVAL_134(plic__EVAL_134),
    ._EVAL_135(plic__EVAL_135),
    ._EVAL_136(plic__EVAL_136),
    ._EVAL_137(plic__EVAL_137),
    ._EVAL_138(plic__EVAL_138),
    ._EVAL_139(plic__EVAL_139),
    ._EVAL_140(plic__EVAL_140),
    ._EVAL_141(plic__EVAL_141),
    ._EVAL_142(plic__EVAL_142),
    ._EVAL_143(plic__EVAL_143),
    ._EVAL_144(plic__EVAL_144)
  );
  assign plic__EVAL_96 = _EVAL_129;
  assign plic__EVAL_33 = _EVAL_2;
  assign plic__EVAL_4 = _EVAL_7;
  assign plic__EVAL_31 = _EVAL_12;
  assign plic__EVAL_114 = _EVAL_79;
  assign plic__EVAL_112 = _EVAL_30;
  assign plic__EVAL_27 = _EVAL_138;
  assign plic__EVAL_38 = _EVAL_87;
  assign plic__EVAL_39 = _EVAL_96;
  assign plic__EVAL = _EVAL_63;
  assign plic__EVAL_109 = _EVAL_89;
  assign plic__EVAL_118 = _EVAL_23;
  assign plic__EVAL_2 = _EVAL_134;
  assign plic__EVAL_53 = _EVAL_29;
  assign plic__EVAL_95 = _EVAL_131;
  assign _EVAL_108 = plic__EVAL_47;
  assign plic__EVAL_75 = _EVAL_45;
  assign plic__EVAL_23 = _EVAL_92;
  assign plic__EVAL_43 = _EVAL_106;
  assign plic__EVAL_9 = _EVAL_38;
  assign plic__EVAL_80 = _EVAL_143;
  assign plic__EVAL_3 = _EVAL_57;
  assign _EVAL_44 = plic__EVAL_124;
  assign plic__EVAL_136 = _EVAL_5;
  assign plic__EVAL_72 = _EVAL_73;
  assign plic__EVAL_107 = _EVAL_90;
  assign plic__EVAL_125 = _EVAL_10;
  assign plic__EVAL_12 = _EVAL_113;
  assign plic__EVAL_111 = _EVAL_95;
  assign plic__EVAL_59 = _EVAL_115;
  assign plic__EVAL_115 = _EVAL_88;
  assign plic__EVAL_92 = _EVAL_35;
  assign plic__EVAL_58 = _EVAL_15;
  assign plic__EVAL_10 = _EVAL_25;
  assign plic__EVAL_117 = _EVAL_137;
  assign plic__EVAL_113 = _EVAL_33;
  assign plic__EVAL_105 = _EVAL_68;
  assign plic__EVAL_94 = _EVAL_54;
  assign plic__EVAL_98 = _EVAL_74;
  assign plic__EVAL_141 = _EVAL_110;
  assign plic__EVAL_14 = _EVAL_17;
  assign _EVAL_11 = plic__EVAL_32;
  assign plic__EVAL_101 = _EVAL_31;
  assign plic__EVAL_120 = _EVAL_123;
  assign plic__EVAL_122 = _EVAL_21;
  assign plic__EVAL_62 = _EVAL_104;
  assign plic__EVAL_55 = _EVAL_72;
  assign plic__EVAL_16 = _EVAL_70;
  assign plic__EVAL_93 = _EVAL_39;
  assign plic__EVAL_99 = _EVAL_94;
  assign plic__EVAL_91 = _EVAL_50;
  assign plic__EVAL_83 = _EVAL_107;
  assign plic__EVAL_87 = _EVAL_28;
  assign plic__EVAL_135 = _EVAL_55;
  assign plic__EVAL_129 = _EVAL_142;
  assign plic__EVAL_139 = _EVAL_16;
  assign plic__EVAL_79 = _EVAL_112;
  assign plic__EVAL_85 = _EVAL_36;
  assign plic__EVAL_45 = _EVAL_85;
  assign plic__EVAL_41 = _EVAL;
  assign plic__EVAL_77 = _EVAL_60;
  assign plic__EVAL_29 = _EVAL_51;
  assign _EVAL_126 = plic__EVAL_19;
  assign plic__EVAL_128 = _EVAL_62;
  assign plic__EVAL_108 = _EVAL_26;
  assign plic__EVAL_65 = _EVAL_139;
  assign plic__EVAL_88 = _EVAL_13;
  assign plic__EVAL_5 = _EVAL_37;
  assign plic__EVAL_0 = _EVAL_56;
  assign plic__EVAL_18 = _EVAL_52;
  assign plic__EVAL_7 = _EVAL_144;
  assign plic__EVAL_34 = _EVAL_101;
  assign plic__EVAL_46 = _EVAL_99;
  assign plic__EVAL_86 = _EVAL_84;
  assign plic__EVAL_25 = _EVAL_22;
  assign _EVAL_128 = plic__EVAL_126;
  assign plic__EVAL_44 = _EVAL_69;
  assign plic__EVAL_89 = _EVAL_111;
  assign plic__EVAL_49 = _EVAL_86;
  assign plic__EVAL_143 = _EVAL_124;
  assign plic__EVAL_40 = _EVAL_78;
  assign plic__EVAL_71 = _EVAL_49;
  assign plic__EVAL_84 = _EVAL_3;
  assign plic__EVAL_70 = _EVAL_102;
  assign plic__EVAL_28 = _EVAL_6;
  assign plic__EVAL_110 = _EVAL_59;
  assign plic__EVAL_104 = _EVAL_41;
  assign plic__EVAL_66 = _EVAL_83;
  assign plic__EVAL_56 = _EVAL_93;
  assign plic__EVAL_140 = _EVAL_4;
  assign plic__EVAL_133 = _EVAL_67;
  assign plic__EVAL_123 = _EVAL_64;
  assign plic__EVAL_57 = _EVAL_77;
  assign plic__EVAL_42 = _EVAL_81;
  assign plic__EVAL_13 = _EVAL_98;
  assign plic__EVAL_6 = _EVAL_80;
  assign plic__EVAL_137 = _EVAL_125;
  assign plic__EVAL_76 = _EVAL_105;
  assign plic__EVAL_54 = _EVAL_47;
  assign plic__EVAL_24 = _EVAL_122;
  assign plic__EVAL_132 = _EVAL_97;
  assign plic__EVAL_134 = _EVAL_75;
  assign plic__EVAL_37 = _EVAL_8;
  assign plic__EVAL_106 = _EVAL_118;
  assign plic__EVAL_11 = _EVAL_135;
  assign plic__EVAL_48 = _EVAL_136;
  assign plic__EVAL_144 = _EVAL_27;
  assign plic__EVAL_73 = _EVAL_117;
  assign _EVAL_140 = plic__EVAL_97;
  assign plic__EVAL_22 = _EVAL_65;
  assign plic__EVAL_131 = _EVAL_127;
  assign plic__EVAL_30 = _EVAL_40;
  assign plic__EVAL_63 = _EVAL_71;
  assign plic__EVAL_52 = _EVAL_66;
  assign plic__EVAL_69 = _EVAL_82;
  assign plic__EVAL_119 = _EVAL_121;
  assign plic__EVAL_1 = _EVAL_103;
  assign plic__EVAL_74 = _EVAL_46;
  assign plic__EVAL_102 = _EVAL_42;
  assign plic__EVAL_90 = _EVAL_1;
  assign plic__EVAL_26 = _EVAL_58;
  assign plic__EVAL_127 = _EVAL_14;
  assign plic__EVAL_67 = _EVAL_119;
  assign plic__EVAL_68 = _EVAL_9;
  assign plic__EVAL_138 = _EVAL_61;
  assign plic__EVAL_8 = _EVAL_32;
  assign plic__EVAL_103 = _EVAL_114;
  assign plic__EVAL_78 = _EVAL_116;
  assign plic__EVAL_82 = _EVAL_18;
  assign plic__EVAL_35 = _EVAL_0;
  assign plic__EVAL_121 = _EVAL_76;
  assign plic__EVAL_50 = _EVAL_130;
  assign plic__EVAL_130 = _EVAL_43;
  assign plic__EVAL_116 = _EVAL_34;
  assign plic__EVAL_100 = _EVAL_100;
  assign plic__EVAL_21 = _EVAL_132;
  assign plic__EVAL_81 = _EVAL_48;
  assign plic__EVAL_61 = _EVAL_120;
  assign _EVAL_19 = plic__EVAL_60;
  assign plic__EVAL_64 = _EVAL_109;
  assign plic__EVAL_36 = _EVAL_91;
  assign plic__EVAL_15 = _EVAL_24;
  assign plic__EVAL_142 = _EVAL_133;
  assign plic__EVAL_17 = _EVAL_141;
  assign plic__EVAL_20 = _EVAL_20;
  assign plic__EVAL_51 = _EVAL_53;
endmodule
