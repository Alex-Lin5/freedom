//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_192(
  output  _EVAL,
  output  _EVAL_0,
  input   _EVAL_1,
  output  _EVAL_2,
  input   _EVAL_3,
  input   _EVAL_4,
  input   _EVAL_5,
  input   _EVAL_6,
  input   _EVAL_7,
  output  _EVAL_8,
  output  _EVAL_9,
  output  _EVAL_10,
  input   _EVAL_11,
  output  _EVAL_12,
  output  _EVAL_13,
  input   _EVAL_14,
  output  _EVAL_15,
  output  _EVAL_16,
  output  _EVAL_17,
  input   _EVAL_18,
  input   _EVAL_19,
  output  _EVAL_20,
  output  _EVAL_21,
  output  _EVAL_22,
  output  _EVAL_23,
  input   _EVAL_24,
  input   _EVAL_25,
  output  _EVAL_26,
  input   _EVAL_27,
  input   _EVAL_28,
  input   _EVAL_29,
  input   _EVAL_30
);
  assign _EVAL_26 = _EVAL_11;
  assign _EVAL_17 = _EVAL_27;
  assign _EVAL = _EVAL_1;
  assign _EVAL_9 = _EVAL_30;
  assign _EVAL_13 = _EVAL_19;
  assign _EVAL_12 = _EVAL_6;
  assign _EVAL_20 = _EVAL_5;
  assign _EVAL_0 = _EVAL_18;
  assign _EVAL_10 = _EVAL_24;
  assign _EVAL_23 = _EVAL_3;
  assign _EVAL_22 = _EVAL_14;
  assign _EVAL_2 = _EVAL_29;
  assign _EVAL_8 = _EVAL_25;
  assign _EVAL_15 = _EVAL_4;
  assign _EVAL_21 = _EVAL_28;
  assign _EVAL_16 = _EVAL_7;
endmodule
