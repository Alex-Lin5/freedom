//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_129(
  output [31:0] _EVAL,
  input  [31:0] _EVAL_0,
  output        _EVAL_1,
  input  [31:0] _EVAL_2,
  input  [3:0]  _EVAL_3,
  output [31:0] _EVAL_4
);
  wire [31:0] _EVAL_5;
  wire  _EVAL_6;
  wire [23:0] _EVAL_7;
  wire [31:0] _EVAL_8;
  wire [31:0] _EVAL_9;
  wire [31:0] _EVAL_10;
  wire [29:0] _EVAL_11;
  wire [31:0] _EVAL_12;
  wire  _EVAL_13;
  wire [31:0] _EVAL_14;
  wire [30:0] _EVAL_15;
  wire  _EVAL_16;
  wire [31:0] _EVAL_17;
  wire [31:0] _EVAL_18;
  wire  _EVAL_19;
  wire [31:0] _EVAL_20;
  wire [29:0] _EVAL_21;
  wire [31:0] _EVAL_22;
  wire [29:0] _EVAL_23;
  wire [31:0] _EVAL_24;
  wire  _EVAL_25;
  wire [31:0] _EVAL_26;
  wire [32:0] _EVAL_27;
  wire [31:0] _EVAL_28;
  wire  _EVAL_29;
  wire [32:0] _EVAL_30;
  wire [31:0] _EVAL_31;
  wire [31:0] _EVAL_32;
  wire [31:0] _EVAL_33;
  wire [31:0] _EVAL_34;
  wire [31:0] _EVAL_35;
  wire [23:0] _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire [4:0] _EVAL_39;
  wire  _EVAL_40;
  wire [31:0] _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire [31:0] _EVAL_44;
  wire [31:0] _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire [31:0] _EVAL_48;
  wire [31:0] _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire [27:0] _EVAL_52;
  wire [31:0] _EVAL_53;
  wire [31:0] _EVAL_54;
  wire [31:0] _EVAL_55;
  wire [31:0] _EVAL_56;
  wire [31:0] _EVAL_57;
  wire [31:0] _EVAL_58;
  wire [31:0] _EVAL_59;
  wire [31:0] _EVAL_60;
  wire  _EVAL_61;
  wire [31:0] _EVAL_62;
  wire [15:0] _EVAL_63;
  wire [31:0] _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire [31:0] _EVAL_67;
  wire [31:0] _EVAL_68;
  wire [23:0] _EVAL_69;
  wire [30:0] _EVAL_70;
  wire [31:0] _EVAL_71;
  wire [15:0] _EVAL_72;
  wire [31:0] _EVAL_73;
  wire [31:0] _EVAL_74;
  wire  _EVAL_75;
  wire [31:0] _EVAL_76;
  wire [31:0] _EVAL_77;
  wire [31:0] _EVAL_78;
  wire  _EVAL_79;
  wire [32:0] _EVAL_80;
  wire [31:0] _EVAL_81;
  wire [31:0] _EVAL_82;
  wire [27:0] _EVAL_83;
  wire [31:0] _EVAL_84;
  wire [15:0] _EVAL_85;
  wire [30:0] _EVAL_86;
  wire [31:0] _EVAL_87;
  wire  _EVAL_88;
  wire [30:0] _EVAL_89;
  wire [31:0] _EVAL_90;
  wire [31:0] _EVAL_91;
  wire [31:0] _EVAL_92;
  wire [31:0] _EVAL_93;
  wire [31:0] _EVAL_94;
  wire [29:0] _EVAL_95;
  wire [27:0] _EVAL_96;
  wire [27:0] _EVAL_97;
  wire [31:0] _EVAL_98;
  wire [32:0] _EVAL_99;
  wire  _EVAL_100;
  wire [31:0] _EVAL_101;
  wire [31:0] _EVAL_102;
  wire [31:0] _EVAL_103;
  wire  _EVAL_104;
  wire [15:0] _EVAL_105;
  wire  _EVAL_106;
  wire [31:0] _EVAL_107;
  wire [31:0] _EVAL_108;
  wire  _EVAL_109;
  wire [23:0] _EVAL_110;
  wire  _EVAL_111;
  wire [31:0] _EVAL_112;
  wire [31:0] _EVAL_113;
  wire [31:0] _EVAL_114;
  wire [31:0] _EVAL_115;
  wire [31:0] _EVAL_116;
  wire  _EVAL_117;
  wire [31:0] _EVAL_118;
  wire  _EVAL_119;
  wire [31:0] _EVAL_120;
  wire [32:0] _EVAL_121;
  wire [31:0] _EVAL_122;
  wire [31:0] _EVAL_123;
  assign _EVAL_116 = _EVAL_102 | _EVAL_67;
  assign _EVAL_4 = _EVAL_27[31:0];
  assign _EVAL_120 = {{8'd0}, _EVAL_110};
  assign _EVAL_70 = _EVAL_107[30:0];
  assign _EVAL_106 = _EVAL_109 & _EVAL_75;
  assign _EVAL_68 = {{8'd0}, _EVAL_7};
  assign _EVAL_40 = _EVAL_3 == 4'h5;
  assign _EVAL_45 = _EVAL_59 | _EVAL_73;
  assign _EVAL_98 = {_EVAL_70, 1'h0};
  assign _EVAL_60 = _EVAL_34 & 32'hf0f0f0f0;
  assign _EVAL_59 = {{16'd0}, _EVAL_85};
  assign _EVAL_53 = _EVAL_92 & 32'hffff0000;
  assign _EVAL_94 = {_EVAL_36, 8'h0};
  assign _EVAL_44 = _EVAL_68 & 32'hff00ff;
  assign _EVAL_73 = _EVAL_91 & 32'hffff0000;
  assign _EVAL_87 = _EVAL_13 ? _EVAL_2 : _EVAL_77;
  assign _EVAL_84 = {_EVAL_69, 8'h0};
  assign _EVAL_74 = _EVAL_12 | _EVAL_49;
  assign _EVAL_77 = _EVAL_35 | _EVAL_18;
  assign _EVAL_71 = _EVAL_120 & 32'hff00ff;
  assign _EVAL_93 = {{31'd0}, _EVAL_42};
  assign _EVAL_101 = {{1'd0}, _EVAL_89};
  assign _EVAL_123 = _EVAL_38 ? _EVAL_74 : 32'h0;
  assign _EVAL_91 = {_EVAL_105, 16'h0};
  assign _EVAL_21 = _EVAL_14[29:0];
  assign _EVAL_24 = _EVAL_108 | _EVAL_114;
  assign _EVAL_28 = _EVAL_122 & 32'hcccccccc;
  assign _EVAL_111 = ~_EVAL_42;
  assign _EVAL_16 = _EVAL_46 | _EVAL_119;
  assign _EVAL_48 = _EVAL_9 | _EVAL_60;
  assign _EVAL_34 = {_EVAL_97, 4'h0};
  assign _EVAL = _EVAL_47 ? _EVAL_4 : _EVAL_116;
  assign _EVAL_12 = _EVAL_5 & 32'h55555555;
  assign _EVAL_90 = _EVAL_78 & 32'h33333333;
  assign _EVAL_27 = _EVAL_32 + _EVAL_93;
  assign _EVAL_51 = _EVAL_87[31];
  assign _EVAL_5 = {{1'd0}, _EVAL_86};
  assign _EVAL_25 = _EVAL_3[1];
  assign _EVAL_58 = {{2'd0}, _EVAL_23};
  assign _EVAL_114 = _EVAL_16 ? _EVAL_103 : 32'h0;
  assign _EVAL_97 = _EVAL_31[27:0];
  assign _EVAL_82 = {_EVAL_21, 2'h0};
  assign _EVAL_107 = _EVAL_90 | _EVAL_28;
  assign _EVAL_11 = _EVAL_48[29:0];
  assign _EVAL_61 = _EVAL_25 ? _EVAL_6 : _EVAL_29;
  assign _EVAL_42 = _EVAL_3[3];
  assign _EVAL_118 = _EVAL_13 ? _EVAL_55 : 32'h0;
  assign _EVAL_15 = _EVAL_41[30:0];
  assign _EVAL_22 = _EVAL_42 ? _EVAL_10 : _EVAL_0;
  assign _EVAL_43 = _EVAL_3 == 4'h4;
  assign _EVAL_96 = _EVAL_64[31:4];
  assign _EVAL_33 = _EVAL_58 & 32'h33333333;
  assign _EVAL_17 = {{16'd0}, _EVAL_63};
  assign _EVAL_69 = _EVAL_56[23:0];
  assign _EVAL_7 = _EVAL_45[31:8];
  assign _EVAL_10 = ~_EVAL_0;
  assign _EVAL_13 = _EVAL_40 | _EVAL_65;
  assign _EVAL_19 = _EVAL_29 == _EVAL_6;
  assign _EVAL_121 = _EVAL_30;
  assign _EVAL_102 = _EVAL_112 | _EVAL_24;
  assign _EVAL_52 = _EVAL_64[27:0];
  assign _EVAL_39 = _EVAL_0[4:0];
  assign _EVAL_6 = _EVAL_0[31];
  assign _EVAL_8 = {{4'd0}, _EVAL_96};
  assign _EVAL_110 = _EVAL_56[31:8];
  assign _EVAL_23 = _EVAL_14[31:2];
  assign _EVAL_92 = {_EVAL_72, 16'h0};
  assign _EVAL_112 = {{31'd0}, _EVAL_106};
  assign _EVAL_56 = _EVAL_17 | _EVAL_53;
  assign _EVAL_85 = _EVAL_55[31:16];
  assign _EVAL_99 = $signed(_EVAL_121) >>> _EVAL_39;
  assign _EVAL_20 = _EVAL_82 & 32'hcccccccc;
  assign _EVAL_81 = _EVAL_84 & 32'hff00ff00;
  assign _EVAL_117 = _EVAL_113 == 32'h0;
  assign _EVAL_54 = {_EVAL_52, 4'h0};
  assign _EVAL_72 = _EVAL_2[15:0];
  assign _EVAL_31 = _EVAL_71 | _EVAL_81;
  assign _EVAL_104 = _EVAL_3 == 4'h0;
  assign _EVAL_32 = _EVAL_80[31:0];
  assign _EVAL_38 = _EVAL_3 == 4'h1;
  assign _EVAL_64 = _EVAL_44 | _EVAL_115;
  assign _EVAL_26 = _EVAL_54 & 32'hf0f0f0f0;
  assign _EVAL_9 = _EVAL_57 & 32'hf0f0f0f;
  assign _EVAL_105 = _EVAL_55[15:0];
  assign _EVAL_113 = _EVAL_2 ^ _EVAL_22;
  assign _EVAL_109 = _EVAL_3 >= 4'hc;
  assign _EVAL_47 = _EVAL_104 | _EVAL_79;
  assign _EVAL_79 = _EVAL_3 == 4'ha;
  assign _EVAL_30 = {_EVAL_66,_EVAL_87};
  assign _EVAL_76 = _EVAL_8 & 32'hf0f0f0f;
  assign _EVAL_115 = _EVAL_94 & 32'hff00ff00;
  assign _EVAL_86 = _EVAL_41[31:1];
  assign _EVAL_119 = _EVAL_3 == 4'h7;
  assign _EVAL_95 = _EVAL_48[31:2];
  assign _EVAL_55 = _EVAL_99[31:0];
  assign _EVAL_14 = _EVAL_76 | _EVAL_26;
  assign _EVAL_49 = _EVAL_62 & 32'haaaaaaaa;
  assign _EVAL_80 = _EVAL_2 + _EVAL_22;
  assign _EVAL_18 = _EVAL_98 & 32'haaaaaaaa;
  assign _EVAL_78 = {{2'd0}, _EVAL_95};
  assign _EVAL_66 = _EVAL_42 & _EVAL_51;
  assign _EVAL_63 = _EVAL_2[31:16];
  assign _EVAL_103 = _EVAL_2 & _EVAL_0;
  assign _EVAL_122 = {_EVAL_11, 2'h0};
  assign _EVAL_75 = _EVAL_19 ? _EVAL_100 : _EVAL_61;
  assign _EVAL_37 = _EVAL_43 | _EVAL_46;
  assign _EVAL_35 = _EVAL_101 & 32'h55555555;
  assign _EVAL_83 = _EVAL_31[31:4];
  assign _EVAL_36 = _EVAL_45[23:0];
  assign _EVAL_89 = _EVAL_107[31:1];
  assign _EVAL_57 = {{4'd0}, _EVAL_83};
  assign _EVAL_50 = _EVAL_111 ? _EVAL_117 : _EVAL_75;
  assign _EVAL_41 = _EVAL_33 | _EVAL_20;
  assign _EVAL_108 = _EVAL_37 ? _EVAL_113 : 32'h0;
  assign _EVAL_67 = _EVAL_118 | _EVAL_123;
  assign _EVAL_88 = _EVAL_3[0];
  assign _EVAL_29 = _EVAL_2[31];
  assign _EVAL_65 = _EVAL_3 == 4'hb;
  assign _EVAL_100 = _EVAL_4[31];
  assign _EVAL_1 = _EVAL_88 ^ _EVAL_50;
  assign _EVAL_46 = _EVAL_3 == 4'h6;
  assign _EVAL_62 = {_EVAL_15, 1'h0};
endmodule
