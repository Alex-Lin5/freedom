//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_53_assert(
  input  [2:0]  _EVAL,
  input  [3:0]  _EVAL_0,
  input         _EVAL_1,
  input  [4:0]  _EVAL_2,
  input  [3:0]  _EVAL_3,
  input  [4:0]  _EVAL_4,
  input  [13:0] _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input  [3:0]  _EVAL_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_16;
  wire [1:0] _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  reg [13:0] _EVAL_23;
  wire  _EVAL_24;
  wire [5:0] _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire [17:0] _EVAL_28;
  wire [5:0] _EVAL_29;
  wire  _EVAL_30;
  wire [17:0] _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire [32:0] _EVAL_43;
  wire [6:0] _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire [3:0] _EVAL_49;
  wire [31:0] _EVAL_50;
  wire  _EVAL_51;
  reg [3:0] _EVAL_52;
  wire [17:0] _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire [6:0] _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire [17:0] _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  reg [5:0] _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire [13:0] _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire [7:0] _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_104;
  wire  _EVAL_106;
  wire [5:0] _EVAL_107;
  wire [2:0] _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  reg [17:0] _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire [7:0] _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  reg [5:0] _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire [17:0] _EVAL_131;
  wire [2:0] _EVAL_132;
  wire  _EVAL_133;
  wire [13:0] _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  reg [2:0] _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire [22:0] _EVAL_145;
  wire  _EVAL_146;
  wire [7:0] _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire [17:0] _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire [31:0] _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_164;
  wire [3:0] _EVAL_165;
  wire [14:0] _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire [3:0] _EVAL_172;
  wire  _EVAL_173;
  wire [5:0] _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire [13:0] _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire [5:0] _EVAL_192;
  reg [5:0] _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  reg [31:0] _EVAL_197;
  wire [31:0] _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire [31:0] _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  reg [2:0] _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  reg [5:0] _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  reg [4:0] _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire [1:0] _EVAL_230;
  wire [7:0] _EVAL_231;
  wire [1:0] _EVAL_232;
  wire  _EVAL_234;
  wire [14:0] _EVAL_235;
  wire [14:0] _EVAL_236;
  wire [17:0] _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire [17:0] _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire [31:0] _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  reg [4:0] _EVAL_256;
  wire  _EVAL_257;
  wire [22:0] _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire [1:0] _EVAL_262;
  wire  _EVAL_263;
  reg [3:0] _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire [5:0] _EVAL_267;
  wire  _EVAL_268;
  wire [3:0] _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire [6:0] _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  reg [2:0] _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire [6:0] _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_294;
  wire  _EVAL_295;
  wire  _EVAL_296;
  wire  _EVAL_297;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_56 = ~_EVAL_61;
  assign _EVAL_142 = _EVAL_189 | _EVAL_14;
  assign _EVAL_95 = _EVAL_109 | _EVAL_213;
  assign _EVAL_271 = _EVAL_208 & _EVAL_290;
  assign _EVAL_34 = _EVAL == 3'h0;
  assign _EVAL_106 = _EVAL_263 & _EVAL_58;
  assign _EVAL_203 = _EVAL_12 == _EVAL_139;
  assign _EVAL_192 = _EVAL_100[7:2];
  assign _EVAL_269 = ~_EVAL_49;
  assign _EVAL_170 = ~_EVAL_292;
  assign _EVAL_258 = 23'hff << _EVAL_0;
  assign _EVAL_159 = _EVAL_214 ? _EVAL_198 : 32'h0;
  assign _EVAL_20 = _EVAL_162 & _EVAL_124;
  assign _EVAL_132 = _EVAL_2[2:0];
  assign _EVAL_126 = _EVAL_7 & _EVAL_259;
  assign _EVAL_251 = _EVAL_12 != 3'h0;
  assign _EVAL_204 = ~_EVAL_69;
  assign _EVAL_64 = _EVAL_75[0];
  assign _EVAL_18 = ~_EVAL_58;
  assign _EVAL_211 = ~_EVAL_73;
  assign _EVAL_37 = _EVAL_271 | _EVAL_14;
  assign _EVAL_155 = _EVAL_9 & _EVAL_156;
  assign _EVAL_111 = _EVAL_172 == 4'h0;
  assign _EVAL_88 = _EVAL == 3'h4;
  assign _EVAL_287 = ~_EVAL_37;
  assign _EVAL_169 = ~_EVAL_137;
  assign _EVAL_240 = _EVAL_50[17:0];
  assign _EVAL_99 = ~_EVAL_19;
  assign _EVAL_280 = _EVAL_41 & _EVAL_290;
  assign _EVAL_172 = _EVAL_15 & _EVAL_269;
  assign _EVAL_104 = _EVAL_289 & _EVAL_221;
  assign _EVAL_109 = _EVAL_81 | _EVAL_114;
  assign _EVAL_77 = _EVAL_4 == 5'h11;
  assign _EVAL_51 = _EVAL_0 == _EVAL_52;
  assign _EVAL_174 = _EVAL_276[5:0];
  assign _EVAL_221 = _EVAL_5[1];
  assign _EVAL_260 = _EVAL_6 == 3'h4;
  assign _EVAL_214 = _EVAL_171 & _EVAL_46;
  assign _EVAL_101 = ~_EVAL_221;
  assign _EVAL_178 = _EVAL_295 | _EVAL_14;
  assign _EVAL_219 = _EVAL_221 & _EVAL_283;
  assign _EVAL_207 = _EVAL_101 & _EVAL_239;
  assign _EVAL_153 = _EVAL_8 | _EVAL_14;
  assign _EVAL_96 = _EVAL_5 ^ 14'h3000;
  assign _EVAL_179 = _EVAL_7 & _EVAL_82;
  assign _EVAL_78 = ~_EVAL_22;
  assign _EVAL_86 = ~_EVAL_120;
  assign _EVAL_141 = _EVAL_81 | _EVAL_104;
  assign _EVAL_32 = ~_EVAL_248;
  assign _EVAL_35 = _EVAL == 3'h5;
  assign _EVAL_206 = _EVAL_263 & _EVAL_254;
  assign _EVAL_165 = ~_EVAL_15;
  assign _EVAL_196 = _EVAL_2 == 5'h8;
  assign _EVAL_156 = _EVAL == 3'h6;
  assign _EVAL_85 = _EVAL_141 | _EVAL_20;
  assign _EVAL_175 = ~_EVAL_65;
  assign _EVAL_87 = _EVAL_188 | _EVAL_14;
  assign _EVAL_27 = _EVAL_41 & _EVAL_113;
  assign _EVAL_255 = _EVAL_27 | _EVAL_117;
  assign _EVAL_276 = _EVAL_125 - 6'h1;
  assign _EVAL_31 = _EVAL_115 >> _EVAL_2;
  assign _EVAL_183 = _EVAL_17 == 2'h0;
  assign _EVAL_149 = _EVAL_111 | _EVAL_14;
  assign _EVAL_296 = ~_EVAL_26;
  assign _EVAL_222 = ~_EVAL_8;
  assign _EVAL_55 = _EVAL_12 <= 3'h2;
  assign _EVAL_152 = _EVAL_162 & _EVAL_219;
  assign _EVAL_75 = _EVAL_131 >> _EVAL_4;
  assign _EVAL_44 = _EVAL_193 - 6'h1;
  assign _EVAL_92 = _EVAL_251 | _EVAL_14;
  assign _EVAL_133 = ~_EVAL_187;
  assign _EVAL_261 = _EVAL_3 == _EVAL_264;
  assign _EVAL_268 = _EVAL_277 | _EVAL_14;
  assign _EVAL_124 = _EVAL_221 & _EVAL_239;
  assign _EVAL_213 = _EVAL_162 & _EVAL_207;
  assign _EVAL_123 = _EVAL_7 & _EVAL_84;
  assign _EVAL_297 = _EVAL_230 == 2'h0;
  assign _EVAL_129 = _EVAL_228 | _EVAL_14;
  assign _EVAL_70 = _EVAL_0 <= 4'hb;
  assign _EVAL_43 = _EVAL_197 + 32'h1;
  assign _EVAL_263 = _EVAL_1 & _EVAL_9;
  assign _EVAL_89 = ~_EVAL_288;
  assign _EVAL_102 = _EVAL_240 != _EVAL_53;
  assign _EVAL_121 = _EVAL_4 == 5'h10;
  assign _EVAL_194 = 4'h6 == _EVAL_0;
  assign _EVAL_108 = _EVAL_4[2:0];
  assign _EVAL_281 = _EVAL_6 <= 3'h6;
  assign _EVAL_184 = _EVAL_6 == 3'h0;
  assign _EVAL_116 = _EVAL_294 & _EVAL_176;
  assign _EVAL_229 = |_EVAL_115;
  assign _EVAL_290 = $signed(_EVAL_235) == 15'sh0;
  assign _EVAL_145 = 23'hff << _EVAL_3;
  assign _EVAL_138 = _EVAL_6 == 3'h5;
  assign _EVAL_26 = _EVAL_272 | _EVAL_14;
  assign _EVAL_91 = ~_EVAL_185;
  assign _EVAL_270 = ~_EVAL_142;
  assign _EVAL_173 = _EVAL == _EVAL_279;
  assign _EVAL_273 = _EVAL_101 & _EVAL_283;
  assign _EVAL_46 = ~_EVAL_202;
  assign _EVAL_228 = _EVAL_167 | _EVAL_196;
  assign _EVAL_16 = ~_EVAL_130;
  assign _EVAL_278 = _EVAL == 3'h3;
  assign _EVAL_154 = _EVAL_109 | _EVAL_54;
  assign _EVAL_234 = _EVAL_220 == 6'h0;
  assign _EVAL_41 = _EVAL_0 <= 4'h2;
  assign _EVAL_47 = ~_EVAL_178;
  assign _EVAL_160 = _EVAL_7 & _EVAL_184;
  assign _EVAL_49 = {_EVAL_85,_EVAL_93,_EVAL_95,_EVAL_154};
  assign _EVAL_71 = plusarg_reader_out == 32'h0;
  assign _EVAL_200 = _EVAL_6[0];
  assign _EVAL_198 = 32'h1 << _EVAL_4;
  assign _EVAL_62 = _EVAL_5 == _EVAL_23;
  assign _EVAL_243 = ~_EVAL_87;
  assign _EVAL_199 = ~_EVAL_67;
  assign _EVAL_50 = _EVAL_206 ? _EVAL_205 : 32'h0;
  assign _EVAL_167 = _EVAL_112 | _EVAL_176;
  assign _EVAL_250 = _EVAL_263 | _EVAL_241;
  assign _EVAL_223 = _EVAL_116 & _EVAL_280;
  assign _EVAL_230 = _EVAL_4[4:3];
  assign _EVAL_171 = _EVAL_241 & _EVAL_234;
  assign _EVAL_24 = ~_EVAL_186;
  assign _EVAL_295 = _EVAL_293 | _EVAL_118;
  assign _EVAL_244 = _EVAL_2 == _EVAL_256;
  assign _EVAL_118 = _EVAL_4 == 5'h8;
  assign _EVAL_74 = _EVAL_110 | _EVAL_14;
  assign _EVAL_210 = _EVAL_12 <= 3'h4;
  assign _EVAL_98 = ~_EVAL_90;
  assign _EVAL_208 = _EVAL_0 <= 4'h8;
  assign _EVAL_117 = _EVAL_70 & _EVAL_195;
  assign _EVAL_266 = _EVAL_7 & _EVAL_260;
  assign _EVAL_128 = _EVAL_9 & _EVAL_88;
  assign _EVAL_286 = ~_EVAL_39;
  assign _EVAL_202 = _EVAL_6 == 3'h6;
  assign _EVAL_274 = _EVAL_102 | _EVAL_217;
  assign _EVAL_212 = _EVAL_7 & _EVAL_202;
  assign _EVAL_275 = _EVAL_291 | _EVAL_238;
  assign _EVAL_42 = _EVAL_2 == 5'h11;
  assign _EVAL_180 = _EVAL_5 & _EVAL_134;
  assign _EVAL_80 = _EVAL_244 | _EVAL_14;
  assign _EVAL_249 = ~_EVAL_21;
  assign _EVAL_191 = _EVAL_194 & _EVAL_196;
  assign _EVAL_110 = _EVAL_255 | _EVAL_191;
  assign _EVAL_224 = _EVAL_297 & _EVAL_168;
  assign _EVAL_61 = _EVAL_275 | _EVAL_14;
  assign _EVAL_127 = _EVAL_165 == 4'h0;
  assign _EVAL_226 = ~_EVAL_97;
  assign _EVAL_231 = _EVAL_258[7:0];
  assign _EVAL_114 = _EVAL_289 & _EVAL_101;
  assign _EVAL_76 = ~_EVAL_74;
  assign _EVAL_38 = ~_EVAL_149;
  assign _EVAL_40 = _EVAL_203 | _EVAL_14;
  assign _EVAL_272 = _EVAL_3 >= 4'h2;
  assign _EVAL_100 = ~_EVAL_231;
  assign _EVAL_282 = ~_EVAL_11;
  assign _EVAL_188 = _EVAL_12 <= 3'h1;
  assign _EVAL_65 = _EVAL_119 | _EVAL_14;
  assign _EVAL_232 = _EVAL_262 | 2'h1;
  assign _EVAL_217 = ~_EVAL_265;
  assign _EVAL_147 = _EVAL_145[7:0];
  assign _EVAL_267 = _EVAL_60[5:0];
  assign _EVAL_158 = ~_EVAL_14;
  assign _EVAL_81 = _EVAL_0 >= 4'h2;
  assign _EVAL_176 = _EVAL_183 & _EVAL_79;
  assign _EVAL_39 = _EVAL_31[0];
  assign _EVAL_135 = ~_EVAL_129;
  assign _EVAL_164 = ~_EVAL_80;
  assign _EVAL_195 = _EVAL_2 == 5'h10;
  assign _EVAL_73 = _EVAL_286 | _EVAL_14;
  assign _EVAL_25 = _EVAL_122[7:2];
  assign _EVAL_148 = ~_EVAL_181;
  assign _EVAL_292 = _EVAL_45 | _EVAL_14;
  assign _EVAL_186 = _EVAL_210 | _EVAL_14;
  assign _EVAL_218 = _EVAL_7 & _EVAL_138;
  assign _EVAL_146 = _EVAL_241 & _EVAL_57;
  assign _EVAL_93 = _EVAL_141 | _EVAL_152;
  assign _EVAL_181 = _EVAL_173 | _EVAL_14;
  assign _EVAL_241 = _EVAL_10 & _EVAL_7;
  assign _EVAL_120 = _EVAL_274 | _EVAL_14;
  assign _EVAL_57 = _EVAL_125 == 6'h0;
  assign _EVAL_119 = _EVAL_180 == 14'h0;
  assign _EVAL_33 = _EVAL == 3'h2;
  assign _EVAL_72 = _EVAL_9 & _EVAL_66;
  assign _EVAL_216 = _EVAL_9 & _EVAL_33;
  assign _EVAL_130 = _EVAL_247 | _EVAL_14;
  assign _EVAL_140 = ~_EVAL_153;
  assign _EVAL_265 = |_EVAL_240;
  assign _EVAL_235 = _EVAL_166;
  assign _EVAL_90 = _EVAL_261 | _EVAL_14;
  assign _EVAL_187 = _EVAL_51 | _EVAL_14;
  assign _EVAL_238 = _EVAL_197 < plusarg_reader_out;
  assign _EVAL_58 = _EVAL_83 == 6'h0;
  assign _EVAL_59 = ~_EVAL_268;
  assign _EVAL_293 = _EVAL_136 | _EVAL_224;
  assign _EVAL_190 = _EVAL_55 | _EVAL_14;
  assign _EVAL_209 = _EVAL_9 & _EVAL_34;
  assign _EVAL_79 = _EVAL_132 <= 3'h6;
  assign _EVAL_285 = _EVAL_83 - 6'h1;
  assign _EVAL_288 = _EVAL_127 | _EVAL_14;
  assign _EVAL_294 = 4'h2 == _EVAL_0;
  assign _EVAL_236 = {1'b0,$signed(_EVAL_96)};
  assign _EVAL_66 = _EVAL == 3'h7;
  assign _EVAL_69 = _EVAL_30 | _EVAL_14;
  assign _EVAL_22 = _EVAL_222 | _EVAL_14;
  assign _EVAL_136 = _EVAL_77 | _EVAL_121;
  assign _EVAL_21 = _EVAL[2];
  assign _EVAL_17 = _EVAL_2[4:3];
  assign _EVAL_150 = ~_EVAL_190;
  assign _EVAL_19 = _EVAL_81 | _EVAL_14;
  assign _EVAL_189 = _EVAL_12 == 3'h0;
  assign _EVAL_262 = 2'h1 << _EVAL_227;
  assign _EVAL_284 = _EVAL_9 & _EVAL_18;
  assign _EVAL_131 = _EVAL_240 | _EVAL_115;
  assign _EVAL_257 = _EVAL_9 & _EVAL_94;
  assign _EVAL_253 = _EVAL_9 & _EVAL_278;
  assign _EVAL_277 = _EVAL_6 == _EVAL_215;
  assign _EVAL_157 = ~_EVAL_63;
  assign _EVAL_254 = _EVAL_193 == 6'h0;
  assign _EVAL_113 = _EVAL_42 | _EVAL_176;
  assign _EVAL_283 = ~_EVAL_239;
  assign _EVAL_30 = _EVAL_4 == _EVAL_225;
  assign _EVAL_122 = ~_EVAL_147;
  assign _EVAL_45 = _EVAL_15 == _EVAL_49;
  assign _EVAL_68 = ~_EVAL_92;
  assign _EVAL_237 = ~_EVAL_53;
  assign _EVAL_248 = _EVAL_282 | _EVAL_14;
  assign _EVAL_161 = _EVAL_9 & _EVAL_35;
  assign _EVAL_259 = ~_EVAL_57;
  assign _EVAL_177 = ~_EVAL_40;
  assign _EVAL_53 = _EVAL_159[17:0];
  assign _EVAL_185 = _EVAL_223 | _EVAL_14;
  assign _EVAL_289 = _EVAL_232[1];
  assign _EVAL_63 = _EVAL_281 | _EVAL_14;
  assign _EVAL_137 = _EVAL_64 | _EVAL_14;
  assign _EVAL_205 = 32'h1 << _EVAL_2;
  assign _EVAL_134 = {{6'd0}, _EVAL_100};
  assign _EVAL_246 = _EVAL_255 & _EVAL_271;
  assign _EVAL_36 = ~_EVAL_229;
  assign _EVAL_94 = _EVAL == 3'h1;
  assign _EVAL_97 = _EVAL_62 | _EVAL_14;
  assign _EVAL_162 = _EVAL_232[0];
  assign _EVAL_29 = _EVAL_44[5:0];
  assign _EVAL_291 = _EVAL_36 | _EVAL_71;
  assign _EVAL_247 = _EVAL_12 <= 3'h3;
  assign _EVAL_151 = _EVAL_115 | _EVAL_240;
  assign _EVAL_84 = _EVAL_6 == 3'h2;
  assign _EVAL_28 = _EVAL_151 & _EVAL_237;
  assign _EVAL_60 = _EVAL_220 - 6'h1;
  assign _EVAL_227 = _EVAL_0[0];
  assign _EVAL_112 = _EVAL_42 | _EVAL_195;
  assign _EVAL_245 = _EVAL_43[31:0];
  assign _EVAL_82 = _EVAL_6 == 3'h1;
  assign _EVAL_166 = $signed(_EVAL_236) & -15'sh1000;
  assign _EVAL_168 = _EVAL_108 <= 3'h6;
  assign _EVAL_67 = _EVAL_246 | _EVAL_14;
  assign _EVAL_54 = _EVAL_162 & _EVAL_273;
  assign _EVAL_107 = _EVAL_285[5:0];
  assign _EVAL_239 = _EVAL_5[0];
  always @(posedge _EVAL_13) begin
    if (_EVAL_106) begin
      _EVAL_23 <= _EVAL_5;
    end
    if (_EVAL_106) begin
      _EVAL_52 <= _EVAL_0;
    end
    if (_EVAL_14) begin
      _EVAL_83 <= 6'h0;
    end else if (_EVAL_263) begin
      if (_EVAL_58) begin
        if (_EVAL_249) begin
          _EVAL_83 <= _EVAL_192;
        end else begin
          _EVAL_83 <= 6'h0;
        end
      end else begin
        _EVAL_83 <= _EVAL_107;
      end
    end
    if (_EVAL_14) begin
      _EVAL_115 <= 18'h0;
    end else begin
      _EVAL_115 <= _EVAL_28;
    end
    if (_EVAL_14) begin
      _EVAL_125 <= 6'h0;
    end else if (_EVAL_241) begin
      if (_EVAL_57) begin
        if (_EVAL_200) begin
          _EVAL_125 <= _EVAL_25;
        end else begin
          _EVAL_125 <= 6'h0;
        end
      end else begin
        _EVAL_125 <= _EVAL_174;
      end
    end
    if (_EVAL_106) begin
      _EVAL_139 <= _EVAL_12;
    end
    if (_EVAL_14) begin
      _EVAL_193 <= 6'h0;
    end else if (_EVAL_263) begin
      if (_EVAL_254) begin
        if (_EVAL_249) begin
          _EVAL_193 <= _EVAL_192;
        end else begin
          _EVAL_193 <= 6'h0;
        end
      end else begin
        _EVAL_193 <= _EVAL_29;
      end
    end
    if (_EVAL_14) begin
      _EVAL_197 <= 32'h0;
    end else if (_EVAL_250) begin
      _EVAL_197 <= 32'h0;
    end else begin
      _EVAL_197 <= _EVAL_245;
    end
    if (_EVAL_146) begin
      _EVAL_215 <= _EVAL_6;
    end
    if (_EVAL_14) begin
      _EVAL_220 <= 6'h0;
    end else if (_EVAL_241) begin
      if (_EVAL_234) begin
        if (_EVAL_200) begin
          _EVAL_220 <= _EVAL_25;
        end else begin
          _EVAL_220 <= 6'h0;
        end
      end else begin
        _EVAL_220 <= _EVAL_267;
      end
    end
    if (_EVAL_146) begin
      _EVAL_225 <= _EVAL_4;
    end
    if (_EVAL_106) begin
      _EVAL_256 <= _EVAL_2;
    end
    if (_EVAL_146) begin
      _EVAL_264 <= _EVAL_3;
    end
    if (_EVAL_106) begin
      _EVAL_279 <= _EVAL;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e0f33ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_211) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(826cecf8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b629a49b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71c39ecd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89a70237)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_287) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1771991a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_287) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3665939)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b8099ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65645413)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1be45b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_287) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a6b9ab7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb678f11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16190f82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee767f72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3cb78501)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32ec0330)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a446ed65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23d30466)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_16) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca302fa5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_7 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6d86346)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10fcdc69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a04bce0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c863aed9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1838bd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98844dc7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_7 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdb613da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd50598)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(389d00df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7e4ecfb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_211) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f0632ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e71f3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f600e79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(779f64b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40394c1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_287) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a55eb4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d482c4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7caf466)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bbcaed52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ac48c7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cf367b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d76159d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b5f582)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aac05ecd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dcd02f16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30c8e430)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_16) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fed7930c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56af9e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28196de8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16038b74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e63e56dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4800cb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a7b646)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ed69334)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d88bdc2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fad9c17b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(603f97b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_287) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e0f33ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6de2c0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83f16ae5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_99) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58ed3ec8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f3fe56a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_99) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9c70f09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b16df594)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fc6389a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d1b5af5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95dda5d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a50d33d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3bea9ce9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b098cf36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f7d1b95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_99) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27a493de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(437751d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_99) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_287) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_216 & _EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e07b5c84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1ef6770)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ce033f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_199) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e73d3d85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d24685e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3ab97d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(47ca2591)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_199) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8802b2c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(711cf76e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a59b2c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae8bfdf1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_23 = _RAND_0[13:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_52 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_83 = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_115 = _RAND_3[17:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_125 = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_139 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_193 = _RAND_6[5:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_197 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_215 = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_220 = _RAND_9[5:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_225 = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_256 = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_264 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_279 = _RAND_13[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
