//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_45_assert(
  input  [3:0]  _EVAL,
  input  [4:0]  _EVAL_0,
  input  [3:0]  _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input  [2:0]  _EVAL_4,
  input         _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  input  [3:0]  _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  input  [31:0] _EVAL_14,
  input         _EVAL_15,
  input  [1:0]  _EVAL_16,
  input         _EVAL_17,
  input  [4:0]  _EVAL_18
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire [1:0] _EVAL_19;
  wire [2:0] _EVAL_20;
  wire [7:0] _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  reg [3:0] _EVAL_29;
  wire  _EVAL_30;
  reg  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire [32:0] _EVAL_38;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire [31:0] _EVAL_41;
  wire [22:0] _EVAL_42;
  wire  _EVAL_43;
  wire [5:0] _EVAL_44;
  wire  _EVAL_45;
  wire [6:0] _EVAL_46;
  wire  _EVAL_47;
  wire [3:0] _EVAL_48;
  wire  _EVAL_49;
  wire [17:0] _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire [31:0] _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire [3:0] _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire [32:0] _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire [32:0] _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire [17:0] _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire [22:0] _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire [32:0] _EVAL_111;
  wire  _EVAL_112;
  wire [5:0] _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire [32:0] _EVAL_120;
  reg [2:0] _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire [32:0] _EVAL_124;
  reg [31:0] _EVAL_125;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire [7:0] _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire [32:0] _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire [31:0] _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire [32:0] _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire [32:0] _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire [17:0] _EVAL_152;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire [1:0] _EVAL_159;
  wire [31:0] _EVAL_160;
  wire [32:0] _EVAL_161;
  wire [32:0] _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire [32:0] _EVAL_168;
  wire [1:0] _EVAL_169;
  reg [5:0] _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire [7:0] _EVAL_175;
  wire [31:0] _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire [32:0] _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire [32:0] _EVAL_195;
  wire [31:0] _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire [5:0] _EVAL_207;
  wire  _EVAL_208;
  wire [31:0] _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire [6:0] _EVAL_215;
  wire  _EVAL_216;
  reg  _EVAL_217;
  wire  _EVAL_218;
  reg [1:0] _EVAL_220;
  wire [32:0] _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire [31:0] _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire [32:0] _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  reg [2:0] _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  reg [3:0] _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire [31:0] _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  reg [4:0] _EVAL_250;
  wire [7:0] _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire [17:0] _EVAL_257;
  wire  _EVAL_258;
  wire [31:0] _EVAL_259;
  wire [32:0] _EVAL_260;
  wire [17:0] _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  reg [31:0] _EVAL_267;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire [5:0] _EVAL_276;
  wire [6:0] _EVAL_277;
  reg [5:0] _EVAL_278;
  wire  _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire [3:0] _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire [32:0] _EVAL_291;
  wire  _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_294;
  wire  _EVAL_295;
  wire [3:0] _EVAL_296;
  wire [31:0] _EVAL_297;
  wire  _EVAL_298;
  reg [17:0] _EVAL_299;
  wire [6:0] _EVAL_300;
  wire [32:0] _EVAL_301;
  wire  _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_307;
  wire  _EVAL_308;
  wire  _EVAL_309;
  wire  _EVAL_310;
  wire  _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire [5:0] _EVAL_314;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_317;
  reg [4:0] _EVAL_318;
  wire  _EVAL_319;
  wire [31:0] _EVAL_320;
  wire  _EVAL_321;
  wire  _EVAL_323;
  reg [5:0] _EVAL_324;
  wire  _EVAL_325;
  wire [17:0] _EVAL_326;
  wire  _EVAL_327;
  wire [17:0] _EVAL_328;
  wire  _EVAL_329;
  wire  _EVAL_330;
  wire  _EVAL_331;
  wire  _EVAL_332;
  wire  _EVAL_333;
  wire  _EVAL_334;
  wire  _EVAL_335;
  wire  _EVAL_336;
  wire  _EVAL_337;
  wire [31:0] _EVAL_338;
  wire  _EVAL_339;
  wire  _EVAL_340;
  wire  _EVAL_341;
  wire [1:0] _EVAL_342;
  wire [17:0] _EVAL_343;
  wire  _EVAL_345;
  wire  _EVAL_346;
  wire  _EVAL_347;
  reg [2:0] _EVAL_348;
  wire  _EVAL_349;
  wire  _EVAL_350;
  wire [32:0] _EVAL_351;
  wire  _EVAL_352;
  wire [5:0] _EVAL_353;
  wire  _EVAL_354;
  wire  _EVAL_355;
  wire  _EVAL_356;
  wire  _EVAL_357;
  wire  _EVAL_358;
  wire [32:0] _EVAL_359;
  wire [2:0] _EVAL_360;
  wire  _EVAL_361;
  wire  _EVAL_362;
  wire  _EVAL_363;
  wire  _EVAL_364;
  wire  _EVAL_365;
  reg [5:0] _EVAL_366;
  wire [32:0] _EVAL_367;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_69 = _EVAL_256 | _EVAL_3;
  assign _EVAL_251 = ~_EVAL_175;
  assign _EVAL_206 = ~_EVAL_47;
  assign _EVAL_187 = _EVAL_159 == 2'h0;
  assign _EVAL_349 = _EVAL_142 | _EVAL_202;
  assign _EVAL_134 = _EVAL_4 == 3'h2;
  assign _EVAL_291 = _EVAL_38;
  assign _EVAL_354 = _EVAL_252 | _EVAL_332;
  assign _EVAL_129 = ~_EVAL_21;
  assign _EVAL_136 = _EVAL_12 == 3'h0;
  assign _EVAL_335 = _EVAL == _EVAL_29;
  assign _EVAL_296 = _EVAL_8 & _EVAL_284;
  assign _EVAL_264 = _EVAL_360 <= 3'h6;
  assign _EVAL_257 = _EVAL_299 >> _EVAL_0;
  assign _EVAL_35 = _EVAL_66 | _EVAL_3;
  assign _EVAL_192 = _EVAL_352 & _EVAL_272;
  assign _EVAL_254 = _EVAL_99 | _EVAL_3;
  assign _EVAL_265 = ~_EVAL_53;
  assign _EVAL_363 = _EVAL_19[0];
  assign _EVAL_49 = ~_EVAL_37;
  assign _EVAL_23 = _EVAL_270 | _EVAL_229;
  assign _EVAL_345 = _EVAL_1 <= 4'hb;
  assign _EVAL_163 = _EVAL_313 | _EVAL_22;
  assign _EVAL_212 = _EVAL_147 | _EVAL_3;
  assign _EVAL_281 = _EVAL_0 == _EVAL_250;
  assign _EVAL_317 = _EVAL_308 | _EVAL_3;
  assign _EVAL_204 = _EVAL_257[0];
  assign _EVAL_140 = _EVAL_269 | _EVAL_3;
  assign _EVAL_359 = {1'b0,$signed(_EVAL_60)};
  assign _EVAL_210 = _EVAL_11 == _EVAL_31;
  assign _EVAL_274 = _EVAL_7 & _EVAL_283;
  assign _EVAL_158 = _EVAL_211 | _EVAL_3;
  assign _EVAL_68 = _EVAL_293 | _EVAL_107;
  assign _EVAL_74 = _EVAL_17 & _EVAL_52;
  assign _EVAL_63 = _EVAL_305 | _EVAL_3;
  assign _EVAL_246 = 32'h1 << _EVAL_0;
  assign _EVAL_293 = _EVAL_99 | _EVAL_192;
  assign _EVAL_64 = ~_EVAL_27;
  assign _EVAL_76 = $signed(_EVAL_124) & -33'sh10000;
  assign _EVAL_301 = _EVAL_260;
  assign _EVAL_215 = _EVAL_324 - 6'h1;
  assign _EVAL_122 = _EVAL_20 <= 3'h6;
  assign _EVAL_186 = _EVAL_2 & _EVAL_7;
  assign _EVAL_197 = ~_EVAL_204;
  assign _EVAL_295 = _EVAL_187 & _EVAL_264;
  assign _EVAL_185 = _EVAL_199 | _EVAL_151;
  assign _EVAL_190 = _EVAL_288 | _EVAL_241;
  assign _EVAL_350 = $signed(_EVAL_143) == 33'sh0;
  assign _EVAL_282 = ~_EVAL_94;
  assign _EVAL_102 = _EVAL_12 == 3'h1;
  assign _EVAL_34 = _EVAL_18 == _EVAL_318;
  assign _EVAL_253 = _EVAL_216 | _EVAL_327;
  assign _EVAL_61 = _EVAL_7 & _EVAL_325;
  assign _EVAL_161 = _EVAL_267 + 32'h1;
  assign _EVAL_237 = 4'h6 == _EVAL_1;
  assign _EVAL_95 = ~_EVAL_321;
  assign _EVAL_201 = _EVAL_248 | _EVAL_77;
  assign _EVAL_171 = $signed(_EVAL_79) == 33'sh0;
  assign _EVAL_224 = ~_EVAL_306;
  assign _EVAL_261 = _EVAL_196[17:0];
  assign _EVAL_279 = _EVAL_12 == _EVAL_348;
  assign _EVAL_149 = ~_EVAL_213;
  assign _EVAL_198 = |_EVAL_299;
  assign _EVAL_309 = _EVAL_355 | _EVAL_3;
  assign _EVAL_227 = _EVAL_334 & _EVAL_150;
  assign _EVAL_168 = $signed(_EVAL_359) & -33'sh400000;
  assign _EVAL_145 = plusarg_reader_out == 32'h0;
  assign _EVAL_160 = _EVAL_14 ^ 32'h3000;
  assign _EVAL_321 = _EVAL_34 | _EVAL_3;
  assign _EVAL_273 = _EVAL_89 & _EVAL_22;
  assign _EVAL_166 = _EVAL_252 | _EVAL_273;
  assign _EVAL_156 = _EVAL_154 | _EVAL_3;
  assign _EVAL_203 = _EVAL_363 & _EVAL_292;
  assign _EVAL_88 = _EVAL_169 == 2'h0;
  assign _EVAL_154 = ~_EVAL_11;
  assign _EVAL_110 = _EVAL_137 & _EVAL_115;
  assign _EVAL_258 = _EVAL_266 | _EVAL_329;
  assign _EVAL_142 = _EVAL_172 | _EVAL_341;
  assign _EVAL_255 = _EVAL_330 & _EVAL_114;
  assign _EVAL_143 = _EVAL_135;
  assign _EVAL_162 = {1'b0,$signed(_EVAL_259)};
  assign _EVAL_300 = _EVAL_278 - 6'h1;
  assign _EVAL_141 = ~_EVAL_174;
  assign _EVAL_194 = _EVAL_354 | _EVAL_3;
  assign _EVAL_208 = _EVAL_199 | _EVAL_285;
  assign _EVAL_328 = _EVAL_261 | _EVAL_299;
  assign _EVAL_195 = _EVAL_168;
  assign _EVAL_294 = ~_EVAL_10;
  assign _EVAL_117 = _EVAL_14[1];
  assign _EVAL_355 = _EVAL_16 == 2'h0;
  assign _EVAL_107 = _EVAL_363 & _EVAL_245;
  assign _EVAL_132 = _EVAL_6 == 3'h0;
  assign _EVAL_176 = _EVAL_14 & _EVAL_297;
  assign _EVAL_242 = ~_EVAL_336;
  assign _EVAL_137 = _EVAL_255 | _EVAL_103;
  assign _EVAL_144 = _EVAL_39 | _EVAL_3;
  assign _EVAL_223 = _EVAL_331 & _EVAL_190;
  assign _EVAL_316 = _EVAL_186 & _EVAL_312;
  assign _EVAL_116 = _EVAL_16 <= 2'h2;
  assign _EVAL_275 = _EVAL_12[0];
  assign _EVAL_218 = ~_EVAL_140;
  assign _EVAL_272 = ~_EVAL_117;
  assign _EVAL_313 = _EVAL_201 | _EVAL_127;
  assign _EVAL_58 = ~_EVAL_319;
  assign _EVAL_106 = _EVAL_4 == 3'h6;
  assign _EVAL_303 = _EVAL_48 == 4'h0;
  assign _EVAL_37 = _EVAL_179 | _EVAL_3;
  assign _EVAL_290 = _EVAL_4 == 3'h1;
  assign _EVAL_42 = 23'hff << _EVAL_1;
  assign _EVAL_108 = 23'hff << _EVAL;
  assign _EVAL_214 = _EVAL_210 | _EVAL_3;
  assign _EVAL_342 = 2'h1 << _EVAL_138;
  assign _EVAL_38 = $signed(_EVAL_234) & -33'sh2000;
  assign _EVAL_337 = _EVAL_17 & _EVAL_62;
  assign _EVAL_306 = _EVAL_110 | _EVAL_3;
  assign _EVAL_285 = _EVAL_363 & _EVAL_78;
  assign _EVAL_307 = _EVAL_18 == 5'h8;
  assign _EVAL_43 = ~_EVAL_214;
  assign _EVAL_269 = _EVAL_12 <= 3'h6;
  assign _EVAL_120 = $signed(_EVAL_162) & -33'sh4000;
  assign _EVAL_70 = _EVAL_197 | _EVAL_3;
  assign _EVAL_216 = _EVAL_0 == 5'h11;
  assign _EVAL_59 = _EVAL_154 | _EVAL_10;
  assign _EVAL_367 = {1'b0,$signed(_EVAL_14)};
  assign _EVAL_191 = ~_EVAL_62;
  assign _EVAL_292 = _EVAL_272 & _EVAL_54;
  assign _EVAL_280 = ~_EVAL_346;
  assign _EVAL_181 = _EVAL_1 <= 4'h8;
  assign _EVAL_305 = _EVAL_176 == 32'h0;
  assign _EVAL_286 = _EVAL_4 == 3'h7;
  assign _EVAL_32 = ~_EVAL_86;
  assign _EVAL_26 = _EVAL_98 | _EVAL_3;
  assign _EVAL_225 = _EVAL_339 ? _EVAL_41 : 32'h0;
  assign _EVAL_252 = _EVAL_181 & _EVAL_87;
  assign _EVAL_196 = _EVAL_316 ? _EVAL_246 : 32'h0;
  assign _EVAL_364 = ~_EVAL_226;
  assign _EVAL_249 = _EVAL_170 == 6'h0;
  assign _EVAL_130 = ~_EVAL_133;
  assign _EVAL_235 = ~_EVAL_194;
  assign _EVAL_297 = {{24'd0}, _EVAL_251};
  assign _EVAL_30 = _EVAL_349 | _EVAL_307;
  assign _EVAL_131 = _EVAL_12 == 3'h4;
  assign _EVAL_50 = _EVAL_152 & _EVAL_326;
  assign _EVAL_351 = {1'b0,$signed(_EVAL_209)};
  assign _EVAL_202 = _EVAL_88 & _EVAL_122;
  assign _EVAL_232 = ~_EVAL_92;
  assign _EVAL_28 = _EVAL_14 == _EVAL_125;
  assign _EVAL_83 = ~_EVAL_323;
  assign _EVAL_276 = _EVAL_46[5:0];
  assign _EVAL_213 = _EVAL_4[2];
  assign _EVAL_205 = ~_EVAL_26;
  assign _EVAL_94 = _EVAL_258 | _EVAL_3;
  assign _EVAL_179 = _EVAL_13 == _EVAL_217;
  assign _EVAL_333 = _EVAL_137 | _EVAL_340;
  assign _EVAL_199 = _EVAL_99 | _EVAL_56;
  assign _EVAL_256 = ~_EVAL_15;
  assign _EVAL_229 = _EVAL_267 < plusarg_reader_out;
  assign _EVAL_175 = _EVAL_42[7:0];
  assign _EVAL_310 = _EVAL_334 & _EVAL_249;
  assign _EVAL_184 = ~_EVAL_165;
  assign _EVAL_334 = _EVAL_5 & _EVAL_17;
  assign _EVAL_356 = _EVAL_6 != 3'h0;
  assign _EVAL_60 = _EVAL_14 ^ 32'hc000000;
  assign _EVAL_343 = _EVAL_328 >> _EVAL_18;
  assign _EVAL_304 = _EVAL_6 <= 3'h2;
  assign _EVAL_51 = _EVAL_59 | _EVAL_3;
  assign _EVAL_89 = _EVAL_1 <= 4'h6;
  assign _EVAL_39 = _EVAL_8 == _EVAL_71;
  assign _EVAL_233 = ~_EVAL_69;
  assign _EVAL_277 = _EVAL_366 - 6'h1;
  assign _EVAL_67 = _EVAL_186 & _EVAL_123;
  assign _EVAL_341 = _EVAL_18 == 5'h10;
  assign _EVAL_55 = _EVAL_4 == _EVAL_121;
  assign _EVAL_146 = _EVAL_186 | _EVAL_334;
  assign _EVAL_157 = _EVAL_16 != 2'h2;
  assign _EVAL_66 = _EVAL_6 <= 3'h4;
  assign _EVAL_148 = {1'b0,$signed(_EVAL_160)};
  assign _EVAL_234 = {1'b0,$signed(_EVAL_139)};
  assign _EVAL_239 = ~_EVAL_63;
  assign _EVAL_221 = $signed(_EVAL_148) & -33'sh1000;
  assign _EVAL_352 = _EVAL_19[1];
  assign _EVAL_159 = _EVAL_0[4:3];
  assign _EVAL_331 = _EVAL_40 & _EVAL_295;
  assign _EVAL_323 = _EVAL_157 | _EVAL_3;
  assign _EVAL_147 = _EVAL_343[0];
  assign _EVAL_302 = _EVAL_1 == _EVAL_243;
  assign _EVAL_128 = _EVAL_17 & _EVAL_102;
  assign _EVAL_222 = _EVAL >= 4'h2;
  assign _EVAL_118 = ~_EVAL_311;
  assign _EVAL_327 = _EVAL_0 == 5'h10;
  assign _EVAL_320 = _EVAL_161[31:0];
  assign _EVAL_99 = _EVAL_1 >= 4'h2;
  assign _EVAL_20 = _EVAL_18[2:0];
  assign _EVAL_332 = _EVAL_89 & _EVAL_85;
  assign _EVAL_100 = _EVAL_89 & _EVAL_180;
  assign _EVAL_101 = _EVAL_225[17:0];
  assign _EVAL_211 = _EVAL_6 == _EVAL_238;
  assign _EVAL_314 = _EVAL_251[7:2];
  assign _EVAL_105 = _EVAL_12 == 3'h2;
  assign _EVAL_361 = _EVAL_7 & _EVAL_289;
  assign _EVAL_247 = _EVAL_7 & _EVAL_286;
  assign _EVAL_357 = _EVAL_4 == 3'h0;
  assign _EVAL_113 = _EVAL_277[5:0];
  assign _EVAL_57 = ~_EVAL_70;
  assign _EVAL_139 = _EVAL_14 ^ 32'h20000000;
  assign _EVAL_97 = ~_EVAL_244;
  assign _EVAL_271 = ~_EVAL_317;
  assign _EVAL_365 = ~_EVAL_144;
  assign _EVAL_92 = _EVAL_223 | _EVAL_3;
  assign _EVAL_104 = ~_EVAL_254;
  assign _EVAL_33 = $signed(_EVAL_301) == 33'sh0;
  assign _EVAL_287 = _EVAL_7 & _EVAL_106;
  assign _EVAL_36 = _EVAL_117 & _EVAL_119;
  assign _EVAL_270 = _EVAL_81 | _EVAL_145;
  assign _EVAL_228 = _EVAL_4 == 3'h5;
  assign _EVAL_330 = _EVAL_1 <= 4'h2;
  assign _EVAL_262 = _EVAL_166 | _EVAL_3;
  assign _EVAL_346 = _EVAL_335 | _EVAL_3;
  assign _EVAL_347 = ~_EVAL_212;
  assign _EVAL_56 = _EVAL_352 & _EVAL_117;
  assign _EVAL_155 = ~_EVAL_35;
  assign _EVAL_98 = _EVAL_16 == _EVAL_220;
  assign _EVAL_173 = _EVAL_93 | _EVAL_3;
  assign _EVAL_78 = _EVAL_117 & _EVAL_54;
  assign _EVAL_123 = _EVAL_366 == 6'h0;
  assign _EVAL_114 = _EVAL_216 | _EVAL_295;
  assign _EVAL_25 = _EVAL_7 & _EVAL_228;
  assign _EVAL_165 = _EVAL_303 | _EVAL_3;
  assign _EVAL_248 = _EVAL_350 | _EVAL_33;
  assign _EVAL_124 = {1'b0,$signed(_EVAL_338)};
  assign _EVAL_127 = $signed(_EVAL_195) == 33'sh0;
  assign _EVAL_72 = ~_EVAL_262;
  assign _EVAL_312 = _EVAL_278 == 6'h0;
  assign _EVAL_47 = _EVAL_23 | _EVAL_3;
  assign _EVAL_62 = _EVAL_12 == 3'h6;
  assign _EVAL_135 = $signed(_EVAL_367) & -33'sh5000;
  assign _EVAL_85 = _EVAL_313 | _EVAL_171;
  assign _EVAL_231 = ~_EVAL_3;
  assign _EVAL_46 = _EVAL_170 - 6'h1;
  assign _EVAL_188 = _EVAL_221;
  assign _EVAL_45 = ~_EVAL_109;
  assign _EVAL_338 = _EVAL_14 ^ 32'h2000000;
  assign _EVAL_172 = _EVAL_18 == 5'h11;
  assign _EVAL_48 = ~_EVAL_8;
  assign _EVAL_44 = _EVAL_129[7:2];
  assign _EVAL_82 = ~_EVAL_158;
  assign _EVAL_169 = _EVAL_18[4:3];
  assign _EVAL_19 = _EVAL_342 | 2'h1;
  assign _EVAL_71 = {_EVAL_208,_EVAL_185,_EVAL_298,_EVAL_68};
  assign _EVAL_151 = _EVAL_363 & _EVAL_36;
  assign _EVAL_21 = _EVAL_108[7:0];
  assign _EVAL_230 = ~_EVAL_236;
  assign _EVAL_22 = $signed(_EVAL_291) == 33'sh0;
  assign _EVAL_41 = 32'h1 << _EVAL_18;
  assign _EVAL_193 = _EVAL_17 & _EVAL_105;
  assign _EVAL_87 = $signed(_EVAL_188) == 33'sh0;
  assign _EVAL_53 = _EVAL_281 | _EVAL_3;
  assign _EVAL_289 = ~_EVAL_123;
  assign _EVAL_178 = ~_EVAL_51;
  assign _EVAL_77 = $signed(_EVAL_111) == 33'sh0;
  assign _EVAL_111 = _EVAL_76;
  assign _EVAL_245 = _EVAL_272 & _EVAL_119;
  assign _EVAL_54 = _EVAL_14[0];
  assign _EVAL_80 = ~_EVAL_84;
  assign _EVAL_133 = _EVAL_356 | _EVAL_3;
  assign _EVAL_189 = _EVAL_17 & _EVAL_136;
  assign _EVAL_207 = _EVAL_300[5:0];
  assign _EVAL_283 = _EVAL_4 == 3'h4;
  assign _EVAL_236 = _EVAL_333 | _EVAL_3;
  assign _EVAL_52 = _EVAL_12 == 3'h5;
  assign _EVAL_90 = _EVAL_17 & _EVAL_177;
  assign _EVAL_180 = _EVAL_163 | _EVAL_171;
  assign _EVAL_79 = _EVAL_120;
  assign _EVAL_40 = 4'h2 == _EVAL_1;
  assign _EVAL_167 = _EVAL_7 & _EVAL_290;
  assign _EVAL_241 = _EVAL_40 & _EVAL_171;
  assign _EVAL_353 = _EVAL_215[5:0];
  assign _EVAL_84 = _EVAL_30 | _EVAL_3;
  assign _EVAL_260 = $signed(_EVAL_351) & -33'sh4000;
  assign _EVAL_150 = _EVAL_324 == 6'h0;
  assign _EVAL_93 = _EVAL_6 <= 3'h3;
  assign _EVAL_174 = _EVAL_222 | _EVAL_3;
  assign _EVAL_325 = _EVAL_4 == 3'h3;
  assign _EVAL_152 = _EVAL_299 | _EVAL_261;
  assign _EVAL_266 = _EVAL_253 | _EVAL_295;
  assign _EVAL_65 = _EVAL_304 | _EVAL_3;
  assign _EVAL_183 = ~_EVAL_173;
  assign _EVAL_326 = ~_EVAL_101;
  assign _EVAL_308 = _EVAL_6 <= 3'h1;
  assign _EVAL_86 = _EVAL_294 | _EVAL_3;
  assign _EVAL_112 = _EVAL_7 & _EVAL_357;
  assign _EVAL_315 = _EVAL_7 & _EVAL_134;
  assign _EVAL_340 = _EVAL_237 & _EVAL_329;
  assign _EVAL_284 = ~_EVAL_71;
  assign _EVAL_164 = _EVAL_296 == 4'h0;
  assign _EVAL_27 = _EVAL_302 | _EVAL_3;
  assign _EVAL_240 = _EVAL_17 & _EVAL_131;
  assign _EVAL_298 = _EVAL_293 | _EVAL_203;
  assign _EVAL_138 = _EVAL_1[0];
  assign _EVAL_339 = _EVAL_227 & _EVAL_191;
  assign _EVAL_319 = _EVAL_164 | _EVAL_3;
  assign _EVAL_244 = _EVAL_116 | _EVAL_3;
  assign _EVAL_177 = ~_EVAL_249;
  assign _EVAL_329 = _EVAL_0 == 5'h8;
  assign _EVAL_81 = ~_EVAL_198;
  assign _EVAL_360 = _EVAL_0[2:0];
  assign _EVAL_103 = _EVAL_345 & _EVAL_327;
  assign _EVAL_115 = _EVAL_252 | _EVAL_100;
  assign _EVAL_358 = _EVAL_115 | _EVAL_3;
  assign _EVAL_200 = ~_EVAL_309;
  assign _EVAL_109 = _EVAL_279 | _EVAL_3;
  assign _EVAL_259 = _EVAL_14 ^ 32'h80000000;
  assign _EVAL_119 = ~_EVAL_54;
  assign _EVAL_288 = _EVAL_330 & _EVAL_87;
  assign _EVAL_362 = ~_EVAL_156;
  assign _EVAL_75 = ~_EVAL_358;
  assign _EVAL_209 = _EVAL_14 ^ 32'h1800000;
  assign _EVAL_226 = _EVAL_132 | _EVAL_3;
  assign _EVAL_311 = _EVAL_55 | _EVAL_3;
  assign _EVAL_336 = _EVAL_28 | _EVAL_3;
  assign _EVAL_263 = ~_EVAL_65;
  always @(posedge _EVAL_9) begin
    if (_EVAL_310) begin
      _EVAL_29 <= _EVAL;
    end
    if (_EVAL_310) begin
      _EVAL_31 <= _EVAL_11;
    end
    if (_EVAL_67) begin
      _EVAL_121 <= _EVAL_4;
    end
    if (_EVAL_67) begin
      _EVAL_125 <= _EVAL_14;
    end
    if (_EVAL_3) begin
      _EVAL_170 <= 6'h0;
    end else if (_EVAL_334) begin
      if (_EVAL_249) begin
        if (_EVAL_275) begin
          _EVAL_170 <= _EVAL_44;
        end else begin
          _EVAL_170 <= 6'h0;
        end
      end else begin
        _EVAL_170 <= _EVAL_276;
      end
    end
    if (_EVAL_310) begin
      _EVAL_217 <= _EVAL_13;
    end
    if (_EVAL_310) begin
      _EVAL_220 <= _EVAL_16;
    end
    if (_EVAL_67) begin
      _EVAL_238 <= _EVAL_6;
    end
    if (_EVAL_67) begin
      _EVAL_243 <= _EVAL_1;
    end
    if (_EVAL_67) begin
      _EVAL_250 <= _EVAL_0;
    end
    if (_EVAL_3) begin
      _EVAL_267 <= 32'h0;
    end else if (_EVAL_146) begin
      _EVAL_267 <= 32'h0;
    end else begin
      _EVAL_267 <= _EVAL_320;
    end
    if (_EVAL_3) begin
      _EVAL_278 <= 6'h0;
    end else if (_EVAL_186) begin
      if (_EVAL_312) begin
        if (_EVAL_149) begin
          _EVAL_278 <= _EVAL_314;
        end else begin
          _EVAL_278 <= 6'h0;
        end
      end else begin
        _EVAL_278 <= _EVAL_207;
      end
    end
    if (_EVAL_3) begin
      _EVAL_299 <= 18'h0;
    end else begin
      _EVAL_299 <= _EVAL_50;
    end
    if (_EVAL_310) begin
      _EVAL_318 <= _EVAL_18;
    end
    if (_EVAL_3) begin
      _EVAL_324 <= 6'h0;
    end else if (_EVAL_334) begin
      if (_EVAL_150) begin
        if (_EVAL_275) begin
          _EVAL_324 <= _EVAL_44;
        end else begin
          _EVAL_324 <= 6'h0;
        end
      end else begin
        _EVAL_324 <= _EVAL_353;
      end
    end
    if (_EVAL_310) begin
      _EVAL_348 <= _EVAL_12;
    end
    if (_EVAL_3) begin
      _EVAL_366 <= 6'h0;
    end else if (_EVAL_186) begin
      if (_EVAL_123) begin
        if (_EVAL_149) begin
          _EVAL_366 <= _EVAL_314;
        end else begin
          _EVAL_366 <= 6'h0;
        end
      end else begin
        _EVAL_366 <= _EVAL_113;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_337 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ace3de25)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_337 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b620c18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_364) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a234bff9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_337 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c3e7e04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_365) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1b9d27e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33c31c55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ddd503f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7a0bd31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3fab353)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_265) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34c8d9bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21724172)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce40d9f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f20b6aeb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39dd47e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4af5038e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_316 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16c8c43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_337 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9aaea86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_265) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(906d45ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db121fc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1b62431)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d821114)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af72db1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_364) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed2d2648)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(893d4a82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52cf224a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b2fe7c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61c21412)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ecd7bba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1eda06b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52c7135b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_364) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5429b8ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf714f84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13904059)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_337 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69a1c2e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d54cc28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39382b76)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(216246a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_365) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_365) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f46aa84a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_364) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17b50b7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5102a618)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13f7170)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2676aea9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_347) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39464ffb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d821114)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbcdde23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53f6fbe0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_365) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e445a1db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f5f7d7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f15b4e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa599725)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_130) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20556b58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b5bdb2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e29f21f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2137b313)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10fa5fa0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccb5c706)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82f1e0e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_364) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(238ca0f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c30fc22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_337 & _EVAL_362) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b422ca09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9717cd10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5a2c80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_337 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b17633ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_316 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b68b2fe0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_232) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2950036c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(baf0b601)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_365) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb347e8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92f3958e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(896b1edd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_232) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afb38415)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25ceaa52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(591478fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a539ebe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e12be32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50c6959d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_365) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccfe40cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45f4131d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_364) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36a9504b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_365) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_365) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa121135)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_274 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27bcf7c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1c952f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_337 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37afda6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_347) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(767d086f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_247 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a35893e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2de7807)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_365) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92dd537a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_337 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9dcc350)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3111ce12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d766562)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_337 & _EVAL_362) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7189bf24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_365) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(add5f6f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_189 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(147cc354)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df27b669)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_29 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_31 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_121 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_125 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_170 = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_217 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_220 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_238 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_243 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_250 = _RAND_9[4:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_267 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_278 = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_299 = _RAND_12[17:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_318 = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_324 = _RAND_14[5:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_348 = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_366 = _RAND_16[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
