//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_15(
  input         _EVAL,
  output        _EVAL_0,
  input  [30:0] _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  output [2:0]  _EVAL_4,
  output        _EVAL_5,
  output [1:0]  _EVAL_6,
  output [3:0]  _EVAL_7,
  input         _EVAL_8,
  input  [31:0] _EVAL_9,
  input         _EVAL_10,
  output [31:0] _EVAL_11,
  output        _EVAL_12,
  input         _EVAL_13,
  output [2:0]  _EVAL_14,
  input  [2:0]  _EVAL_15,
  input         _EVAL_16,
  input  [3:0]  _EVAL_17,
  output [2:0]  _EVAL_18,
  output        _EVAL_19,
  input  [2:0]  _EVAL_20,
  input  [2:0]  _EVAL_21,
  output [31:0] _EVAL_22,
  input  [4:0]  _EVAL_23,
  output        _EVAL_24,
  output [30:0] _EVAL_25,
  output        _EVAL_26,
  input         _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  input  [31:0] _EVAL_30,
  output [1:0]  _EVAL_31,
  input         _EVAL_32,
  output [2:0]  _EVAL_33,
  output [4:0]  _EVAL_34
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire [5:0] _EVAL_39;
  wire [1:0] _EVAL_40;
  reg [2:0] _EVAL_41;
  wire  _EVAL_42;
  wire [1:0] _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire [2:0] q__EVAL;
  wire  q__EVAL_0;
  wire [2:0] q__EVAL_1;
  wire  q__EVAL_2;
  wire  q__EVAL_3;
  wire [31:0] q__EVAL_4;
  wire [4:0] q__EVAL_5;
  wire [31:0] q__EVAL_6;
  wire  q__EVAL_7;
  wire [4:0] q__EVAL_8;
  wire  q__EVAL_9;
  wire  q__EVAL_10;
  wire  q__EVAL_11;
  wire [2:0] q__EVAL_12;
  wire  q__EVAL_13;
  wire [1:0] q__EVAL_14;
  wire  q__EVAL_15;
  wire  q__EVAL_16;
  wire [2:0] q__EVAL_17;
  wire  q__EVAL_18;
  wire  _EVAL_47;
  wire  _EVAL_49;
  wire  _EVAL_50;
  reg  _EVAL_51;
  wire  _EVAL_52;
  reg  _EVAL_53;
  wire [3:0] _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire [3:0] _EVAL_57;
  reg  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_64;
  wire [24:0] _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire [2:0] _EVAL_71;
  wire  _EVAL_73;
  wire  _EVAL_75;
  wire [30:0] _EVAL_76;
  reg [31:0] _EVAL_77;
  wire  _EVAL_78;
  wire [5:0] _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_85;
  wire [30:0] _EVAL_86;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire [12:0] _EVAL_90;
  reg  _EVAL_91;
  reg  _EVAL_92;
  wire  _EVAL_93;
  wire [3:0] _EVAL_94;
  wire  _EVAL_95;
  wire [1:0] _EVAL_96;
  wire  _EVAL_98;
  reg [2:0] _EVAL_101;
  wire [3:0] _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire [1:0] _EVAL_105;
  wire  _EVAL_107;
  wire  _EVAL_108;
  reg  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_116;
  wire [30:0] _EVAL_117;
  wire  _EVAL_119;
  wire  _EVAL_122;
  wire [2:0] _EVAL_125;
  wire [1:0] _EVAL_127;
  wire [3:0] _EVAL_129;
  wire [30:0] _EVAL_130;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire [30:0] _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire [1:0] _EVAL_137;
  wire  _EVAL_139;
  wire [3:0] _EVAL_140;
  reg  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  reg  _EVAL_146;
  wire [1:0] _EVAL_148;
  wire [2:0] _EVAL_149;
  wire [3:0] _EVAL_150;
  reg [2:0] _EVAL_151;
  reg  _EVAL_152;
  reg  _EVAL_153;
  wire  _EVAL_156;
  wire [5:0] _EVAL_157;
  wire [30:0] _EVAL_158;
  reg [2:0] _EVAL_159;
  wire [30:0] _EVAL_160;
  wire [4:0] _EVAL_161;
  wire [1:0] _EVAL_162;
  wire [2:0] _EVAL_166;
  wire  _EVAL_167;
  reg  _EVAL_168;
  reg  _EVAL_169;
  wire [1:0] _EVAL_170;
  wire [27:0] _EVAL_172;
  wire [2:0] _EVAL_174;
  reg [1:0] _EVAL_175;
  reg [4:0] _EVAL_176;
  wire  _EVAL_177;
  wire [5:0] _EVAL_178;
  reg [30:0] _EVAL_179;
  reg  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  reg [4:0] _EVAL_184;
  wire  _EVAL_187;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  reg [31:0] _EVAL_192;
  reg  _EVAL_195;
  wire [3:0] _EVAL_196;
  wire  _EVAL_198;
  wire  _EVAL_200;
  wire [6:0] _EVAL_201;
  _EVAL_14 q (
    ._EVAL(q__EVAL),
    ._EVAL_0(q__EVAL_0),
    ._EVAL_1(q__EVAL_1),
    ._EVAL_2(q__EVAL_2),
    ._EVAL_3(q__EVAL_3),
    ._EVAL_4(q__EVAL_4),
    ._EVAL_5(q__EVAL_5),
    ._EVAL_6(q__EVAL_6),
    ._EVAL_7(q__EVAL_7),
    ._EVAL_8(q__EVAL_8),
    ._EVAL_9(q__EVAL_9),
    ._EVAL_10(q__EVAL_10),
    ._EVAL_11(q__EVAL_11),
    ._EVAL_12(q__EVAL_12),
    ._EVAL_13(q__EVAL_13),
    ._EVAL_14(q__EVAL_14),
    ._EVAL_15(q__EVAL_15),
    ._EVAL_16(q__EVAL_16),
    ._EVAL_17(q__EVAL_17),
    ._EVAL_18(q__EVAL_18)
  );
  assign _EVAL_80 = _EVAL_135 & _EVAL_144;
  assign _EVAL_52 = _EVAL_45 | _EVAL_183;
  assign _EVAL_125 = _EVAL_116 ? _EVAL_15 : 3'h2;
  assign q__EVAL_1 = {{1'd0}, _EVAL_137};
  assign _EVAL_172 = _EVAL_76[30:3];
  assign q__EVAL_8 = _EVAL_184;
  assign _EVAL_107 = |_EVAL_172;
  assign _EVAL_25 = _EVAL_179;
  assign _EVAL_64 = ~_EVAL_169;
  assign _EVAL_47 = ~_EVAL_181;
  assign _EVAL_68 = _EVAL_21 == 3'h5;
  assign _EVAL_59 = _EVAL_27 | _EVAL_145;
  assign _EVAL_50 = _EVAL_45 ? _EVAL_153 : _EVAL_93;
  assign _EVAL_78 = ~_EVAL_153;
  assign _EVAL_156 = _EVAL_146 & _EVAL_55;
  assign _EVAL_140 = _EVAL_104 ? {{1'd0}, _EVAL_101} : _EVAL_57;
  assign _EVAL_170 = _EVAL_195 ? 2'h2 : 2'h3;
  assign _EVAL_178 = _EVAL_201[5:0];
  assign _EVAL_69 = _EVAL_104 ? _EVAL_153 : _EVAL_50;
  assign _EVAL_88 = ~_EVAL_187;
  assign _EVAL_39 = _EVAL_179[5:0];
  assign _EVAL_24 = q__EVAL_10;
  assign _EVAL_162 = {{1'd0}, _EVAL_89};
  assign _EVAL_187 = _EVAL_21[2];
  assign _EVAL_26 = q__EVAL_2;
  assign _EVAL_104 = _EVAL_146 & _EVAL_42;
  assign _EVAL_67 = _EVAL_179[30:6];
  assign _EVAL_160 = {{25'd0}, _EVAL_157};
  assign _EVAL_46 = _EVAL_45 ? _EVAL_195 : _EVAL_119;
  assign _EVAL_148 = _EVAL_174[1:0];
  assign _EVAL_95 = _EVAL_144 | _EVAL;
  assign _EVAL_98 = _EVAL_146 & _EVAL_113;
  assign _EVAL_6 = _EVAL_156 ? _EVAL_170 : _EVAL_44;
  assign _EVAL_11 = _EVAL_192;
  assign _EVAL_177 = _EVAL_104 | _EVAL_52;
  assign _EVAL_4 = q__EVAL_12;
  assign _EVAL_110 = _EVAL_94[3];
  assign _EVAL_174 = _EVAL_175 + _EVAL_162;
  assign _EVAL_166 = _EVAL_140[2:0];
  assign _EVAL_108 = _EVAL_16 | _EVAL_141;
  assign q__EVAL_4 = _EVAL_9;
  assign _EVAL_36 = _EVAL_191 & _EVAL_182;
  assign _EVAL_129 = {1'h0,_EVAL_15};
  assign _EVAL_76 = _EVAL_160 & _EVAL_86;
  assign _EVAL_136 = _EVAL_175 >= 2'h3;
  assign _EVAL_135 = ~_EVAL_136;
  assign _EVAL_70 = ~_EVAL_107;
  assign _EVAL_96 = {_EVAL_92,_EVAL_198};
  assign _EVAL_142 = _EVAL_191 | _EVAL_177;
  assign _EVAL_75 = _EVAL_98 & _EVAL_59;
  assign _EVAL_143 = _EVAL_177 ? _EVAL_200 : _EVAL_135;
  assign _EVAL_31 = q__EVAL_14;
  assign _EVAL_71 = _EVAL_94[2:0];
  assign _EVAL_40 = {_EVAL_109,_EVAL_53};
  assign _EVAL_157 = ~_EVAL_79;
  assign _EVAL_55 = ~_EVAL_91;
  assign _EVAL_144 = ~_EVAL_168;
  assign _EVAL_5 = _EVAL_168;
  assign _EVAL_161 = _EVAL_129 - 4'h3;
  assign q__EVAL_3 = _EVAL_103 & _EVAL_47;
  assign _EVAL_201 = _EVAL_39 + 6'h4;
  assign _EVAL_19 = _EVAL_104 ? 1'h0 : _EVAL_143;
  assign _EVAL_85 = _EVAL_27 | _EVAL_181;
  assign _EVAL_196 = _EVAL_116 ? 4'h0 : _EVAL_102;
  assign _EVAL_133 = _EVAL_104 ? 1'h0 : _EVAL_143;
  assign _EVAL_117 = {_EVAL_67,_EVAL_178};
  assign _EVAL_33 = _EVAL_101;
  assign q__EVAL_18 = _EVAL_10;
  assign _EVAL_150 = {_EVAL_71, 1'h0};
  assign _EVAL_60 = _EVAL_169 ? 1'h0 : 1'h1;
  assign _EVAL_89 = _EVAL_104 ? 1'h0 : _EVAL_35;
  assign _EVAL_18 = _EVAL_41;
  assign _EVAL_183 = _EVAL_152 & _EVAL_78;
  assign _EVAL_130 = _EVAL_104 ? _EVAL_179 : _EVAL_134;
  assign _EVAL_102 = _EVAL_150 | 4'h1;
  assign _EVAL_54 = _EVAL_36 ? _EVAL_196 : {{1'd0}, _EVAL_101};
  assign _EVAL_119 = _EVAL_183 ? 1'h0 : 1'h1;
  assign q__EVAL_11 = _EVAL_8;
  assign _EVAL_200 = _EVAL_135 & _EVAL_168;
  assign _EVAL_12 = q__EVAL_9;
  assign _EVAL_14 = q__EVAL_17;
  assign _EVAL_182 = ~_EVAL_68;
  assign _EVAL_134 = _EVAL_45 ? _EVAL_179 : _EVAL_158;
  assign _EVAL_56 = _EVAL_49 | _EVAL_181;
  assign _EVAL_158 = _EVAL_183 ? _EVAL_117 : _EVAL_179;
  assign q__EVAL_7 = _EVAL_122 & _EVAL_47;
  assign _EVAL_57 = _EVAL_177 ? {{1'd0}, _EVAL_101} : _EVAL_54;
  assign _EVAL_0 = q__EVAL_0;
  assign _EVAL_79 = _EVAL_90[5:0];
  assign _EVAL_94 = _EVAL_161[3:0];
  assign _EVAL_116 = _EVAL_68 | _EVAL_110;
  assign _EVAL_42 = ~_EVAL_59;
  assign _EVAL_198 = ~_EVAL_58;
  assign _EVAL_73 = q__EVAL_10;
  assign _EVAL_190 = _EVAL_104 ? _EVAL_195 : _EVAL_46;
  assign _EVAL_113 = _EVAL_153 | _EVAL_144;
  assign _EVAL_103 = _EVAL_16 & _EVAL_64;
  assign _EVAL_44 = _EVAL_195 ? 2'h0 : 2'h1;
  assign _EVAL_93 = _EVAL_183 ? _EVAL_70 : _EVAL_153;
  assign _EVAL_35 = _EVAL_177 ? _EVAL_80 : _EVAL_191;
  assign _EVAL_149 = _EVAL_148 - _EVAL_105;
  assign _EVAL_127 = _EVAL_149[1:0];
  assign _EVAL_137 = _EVAL_181 ? 2'h2 : {{1'd0}, _EVAL_60};
  assign _EVAL_34 = q__EVAL_5;
  assign _EVAL_139 = _EVAL_191 | _EVAL_104;
  assign q__EVAL_15 = _EVAL_51 & _EVAL_85;
  assign _EVAL_22 = q__EVAL_6;
  assign _EVAL_122 = _EVAL_108 & _EVAL_169;
  assign _EVAL_45 = _EVAL_152 & _EVAL_167;
  assign _EVAL_112 = _EVAL_59 & _EVAL_146;
  assign _EVAL_167 = ~_EVAL_146;
  assign q__EVAL_16 = _EVAL_28;
  assign q__EVAL = _EVAL_151;
  assign _EVAL_105 = {{1'd0}, _EVAL_189};
  assign _EVAL_7 = {_EVAL_40,_EVAL_96};
  assign _EVAL_49 = ~_EVAL_51;
  assign _EVAL_86 = ~_EVAL_179;
  assign _EVAL_90 = 13'h3f << _EVAL_159;
  assign _EVAL_132 = _EVAL_135 & _EVAL_95;
  assign _EVAL_191 = _EVAL_133 & _EVAL;
  assign _EVAL_189 = _EVAL_8 & _EVAL_73;
  assign _EVAL_145 = _EVAL_91 & _EVAL_56;
  always @(posedge _EVAL_28) begin
    if (_EVAL_10) begin
      _EVAL_41 <= 3'h0;
    end else if (!(_EVAL_104)) begin
      if (!(_EVAL_177)) begin
        if (_EVAL_36) begin
          _EVAL_41 <= _EVAL_125;
        end
      end
    end
    if (_EVAL_10) begin
      _EVAL_51 <= 1'h0;
    end else if (_EVAL_85) begin
      _EVAL_51 <= _EVAL_75;
    end
    if (_EVAL_10) begin
      _EVAL_53 <= 1'h0;
    end else if (!(_EVAL_104)) begin
      if (!(_EVAL_177)) begin
        if (_EVAL_191) begin
          _EVAL_53 <= _EVAL_2;
        end
      end
    end
    if (_EVAL_10) begin
      _EVAL_58 <= 1'h0;
    end else if (!(_EVAL_104)) begin
      if (!(_EVAL_177)) begin
        if (_EVAL_191) begin
          _EVAL_58 <= _EVAL_3;
        end
      end
    end
    if (!(_EVAL_104)) begin
      if (_EVAL_177) begin
        _EVAL_77 <= _EVAL_30;
      end else if (_EVAL_36) begin
        _EVAL_77 <= _EVAL_30;
      end
    end
    if (!(_EVAL_104)) begin
      if (!(_EVAL_177)) begin
        if (_EVAL_191) begin
          _EVAL_91 <= _EVAL_68;
        end
      end
    end
    if (_EVAL_10) begin
      _EVAL_92 <= 1'h0;
    end else if (!(_EVAL_104)) begin
      if (!(_EVAL_177)) begin
        if (_EVAL_191) begin
          _EVAL_92 <= _EVAL_29;
        end
      end
    end
    if (_EVAL_10) begin
      _EVAL_101 <= 3'h0;
    end else begin
      _EVAL_101 <= _EVAL_166;
    end
    if (_EVAL_10) begin
      _EVAL_109 <= 1'h0;
    end else if (!(_EVAL_104)) begin
      if (!(_EVAL_177)) begin
        if (_EVAL_191) begin
          _EVAL_109 <= _EVAL_13;
        end
      end
    end
    if (_EVAL_85) begin
      if (_EVAL_195) begin
        _EVAL_141 <= 1'h0;
      end else begin
        _EVAL_141 <= _EVAL_108;
      end
    end
    if (_EVAL_10) begin
      _EVAL_146 <= 1'h0;
    end else if (_EVAL_104) begin
      _EVAL_146 <= _EVAL_104;
    end else if (_EVAL_177) begin
      _EVAL_146 <= _EVAL_132;
    end else begin
      _EVAL_146 <= _EVAL_139;
    end
    if (_EVAL_112) begin
      _EVAL_151 <= _EVAL_159;
    end
    if (_EVAL_10) begin
      _EVAL_152 <= 1'h0;
    end else if (_EVAL_104) begin
      _EVAL_152 <= _EVAL_177;
    end else if (_EVAL_177) begin
      _EVAL_152 <= _EVAL_177;
    end else begin
      _EVAL_152 <= _EVAL_142;
    end
    if (_EVAL_104) begin
      _EVAL_153 <= _EVAL_69;
    end else if (_EVAL_177) begin
      _EVAL_153 <= _EVAL_69;
    end else if (_EVAL_191) begin
      _EVAL_153 <= _EVAL_116;
    end else begin
      _EVAL_153 <= _EVAL_69;
    end
    if (!(_EVAL_104)) begin
      if (!(_EVAL_177)) begin
        if (_EVAL_191) begin
          _EVAL_159 <= _EVAL_15;
        end
      end
    end
    if (_EVAL_10) begin
      _EVAL_168 <= 1'h0;
    end else if (!(_EVAL_104)) begin
      if (!(_EVAL_177)) begin
        if (_EVAL_36) begin
          _EVAL_168 <= _EVAL_88;
        end
      end
    end
    if (_EVAL_10) begin
      _EVAL_169 <= 1'h0;
    end else if (_EVAL_112) begin
      _EVAL_169 <= _EVAL_168;
    end
    if (_EVAL_10) begin
      _EVAL_175 <= 2'h0;
    end else begin
      _EVAL_175 <= _EVAL_127;
    end
    if (!(_EVAL_104)) begin
      if (!(_EVAL_177)) begin
        if (_EVAL_191) begin
          _EVAL_176 <= _EVAL_23;
        end
      end
    end
    if (_EVAL_10) begin
      _EVAL_179 <= 31'h0;
    end else if (_EVAL_104) begin
      _EVAL_179 <= _EVAL_130;
    end else if (_EVAL_177) begin
      _EVAL_179 <= _EVAL_130;
    end else if (_EVAL_36) begin
      _EVAL_179 <= _EVAL_1;
    end else begin
      _EVAL_179 <= _EVAL_130;
    end
    if (_EVAL_112) begin
      _EVAL_181 <= _EVAL_91;
    end
    if (_EVAL_112) begin
      _EVAL_184 <= _EVAL_176;
    end
    if (_EVAL_59) begin
      _EVAL_192 <= _EVAL_77;
    end
    _EVAL_195 <= _EVAL_10 | _EVAL_190;
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_41 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_51 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_53 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_58 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_77 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_91 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_92 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_101 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_109 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_141 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_146 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_151 = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_152 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_153 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_159 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_168 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_169 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _EVAL_175 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  _EVAL_176 = _RAND_18[4:0];
  _RAND_19 = {1{`RANDOM}};
  _EVAL_179 = _RAND_19[30:0];
  _RAND_20 = {1{`RANDOM}};
  _EVAL_181 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _EVAL_184 = _RAND_21[4:0];
  _RAND_22 = {1{`RANDOM}};
  _EVAL_192 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  _EVAL_195 = _RAND_23[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
