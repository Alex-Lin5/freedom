//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_51_assert(
  input  [3:0]  _EVAL,
  input         _EVAL_0,
  input  [1:0]  _EVAL_1,
  input  [2:0]  _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input  [31:0] _EVAL_5,
  input  [4:0]  _EVAL_6,
  input  [2:0]  _EVAL_7,
  input         _EVAL_8,
  input  [3:0]  _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [3:0]  _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input  [4:0]  _EVAL_17,
  input         _EVAL_18
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire [32:0] _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire [1:0] _EVAL_23;
  wire [31:0] _EVAL_24;
  wire  _EVAL_25;
  wire [31:0] _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  reg [4:0] _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire [32:0] _EVAL_34;
  reg  _EVAL_35;
  wire  _EVAL_36;
  wire [32:0] _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire [31:0] _EVAL_41;
  wire  _EVAL_42;
  wire [6:0] _EVAL_43;
  reg [2:0] _EVAL_44;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire [32:0] _EVAL_49;
  wire [32:0] _EVAL_50;
  wire  _EVAL_51;
  wire [17:0] _EVAL_52;
  wire  _EVAL_53;
  wire [22:0] _EVAL_54;
  wire  _EVAL_55;
  wire [31:0] _EVAL_56;
  wire [3:0] _EVAL_57;
  wire [7:0] _EVAL_58;
  wire  _EVAL_59;
  wire [32:0] _EVAL_60;
  wire  _EVAL_61;
  wire [6:0] _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire [17:0] _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire [1:0] _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  reg [3:0] _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire [5:0] _EVAL_99;
  wire [31:0] _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire [17:0] _EVAL_108;
  wire  _EVAL_109;
  wire [3:0] _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire [17:0] _EVAL_117;
  wire  _EVAL_118;
  wire [31:0] _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire [32:0] _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  reg [5:0] _EVAL_129;
  wire [32:0] _EVAL_130;
  wire  _EVAL_131;
  wire [3:0] _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire [32:0] _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire [17:0] _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire [5:0] _EVAL_146;
  wire [2:0] _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  reg [5:0] _EVAL_150;
  wire [1:0] _EVAL_151;
  wire  _EVAL_152;
  wire [5:0] _EVAL_153;
  wire [31:0] _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire [32:0] _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  reg [4:0] _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire [3:0] _EVAL_168;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire [32:0] _EVAL_172;
  wire [32:0] _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  reg [31:0] _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire [5:0] _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  reg [2:0] _EVAL_213;
  wire  _EVAL_214;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire [17:0] _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  reg [3:0] _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire [31:0] _EVAL_234;
  wire  _EVAL_235;
  wire [31:0] _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire [32:0] _EVAL_240;
  wire [32:0] _EVAL_241;
  wire  _EVAL_242;
  wire [32:0] _EVAL_243;
  reg [1:0] _EVAL_245;
  wire  _EVAL_246;
  wire [2:0] _EVAL_247;
  wire  _EVAL_248;
  reg [5:0] _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire [31:0] _EVAL_255;
  wire  _EVAL_256;
  reg [17:0] _EVAL_257;
  reg [31:0] _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire [32:0] _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  reg [5:0] _EVAL_278;
  reg [2:0] _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire [5:0] _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_294;
  wire [6:0] _EVAL_295;
  wire  _EVAL_296;
  wire [6:0] _EVAL_297;
  wire  _EVAL_298;
  wire [32:0] _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire [7:0] _EVAL_302;
  wire  _EVAL_303;
  wire [31:0] _EVAL_304;
  wire [32:0] _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_307;
  wire [17:0] _EVAL_308;
  wire  _EVAL_309;
  wire  _EVAL_310;
  wire [7:0] _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_317;
  wire  _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_321;
  wire  _EVAL_322;
  wire  _EVAL_323;
  wire  _EVAL_324;
  wire  _EVAL_325;
  wire  _EVAL_326;
  wire  _EVAL_327;
  wire [31:0] _EVAL_329;
  wire  _EVAL_330;
  wire  _EVAL_331;
  wire  _EVAL_332;
  wire  _EVAL_333;
  wire  _EVAL_334;
  wire  _EVAL_335;
  wire  _EVAL_336;
  wire  _EVAL_337;
  wire [17:0] _EVAL_338;
  wire [22:0] _EVAL_339;
  wire  _EVAL_340;
  wire  _EVAL_341;
  wire [32:0] _EVAL_342;
  wire  _EVAL_343;
  wire  _EVAL_344;
  wire  _EVAL_345;
  wire  _EVAL_346;
  wire  _EVAL_347;
  wire  _EVAL_348;
  wire  _EVAL_349;
  reg  _EVAL_350;
  wire  _EVAL_351;
  wire  _EVAL_352;
  wire  _EVAL_353;
  wire  _EVAL_354;
  wire  _EVAL_355;
  wire  _EVAL_356;
  wire [31:0] _EVAL_357;
  wire  _EVAL_358;
  wire [1:0] _EVAL_359;
  wire [32:0] _EVAL_360;
  wire  _EVAL_361;
  wire  _EVAL_362;
  wire [5:0] _EVAL_364;
  wire  _EVAL_365;
  wire  _EVAL_366;
  wire  _EVAL_367;
  wire [7:0] _EVAL_368;
  wire  _EVAL_369;
  wire  _EVAL_370;
  wire  _EVAL_371;
  wire [32:0] _EVAL_372;
  wire  _EVAL_373;
  wire [32:0] _EVAL_374;
  wire  _EVAL_375;
  wire  _EVAL_376;
  wire  _EVAL_377;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_339 = 23'hff << _EVAL;
  assign _EVAL_98 = ~_EVAL_292;
  assign _EVAL_293 = $signed(_EVAL_49) == 33'sh0;
  assign _EVAL_353 = _EVAL_229 & _EVAL_315;
  assign _EVAL_49 = _EVAL_50;
  assign _EVAL_151 = 2'h1 << _EVAL_319;
  assign _EVAL_292 = _EVAL_202 | _EVAL_4;
  assign _EVAL_333 = _EVAL_277 & _EVAL_88;
  assign _EVAL_20 = _EVAL_77 | _EVAL_4;
  assign _EVAL_234 = {{24'd0}, _EVAL_302};
  assign _EVAL_255 = _EVAL_5 & _EVAL_234;
  assign _EVAL_37 = _EVAL_360;
  assign _EVAL_368 = ~_EVAL_58;
  assign _EVAL_165 = _EVAL_33 | _EVAL_4;
  assign _EVAL_205 = ~_EVAL_69;
  assign _EVAL_370 = ~_EVAL_294;
  assign _EVAL_110 = ~_EVAL_13;
  assign _EVAL_302 = ~_EVAL_311;
  assign _EVAL_259 = _EVAL_367 & _EVAL_334;
  assign _EVAL_104 = _EVAL_12 == _EVAL_213;
  assign _EVAL_194 = _EVAL_224 | _EVAL_4;
  assign _EVAL_268 = _EVAL_201 | _EVAL_322;
  assign _EVAL_63 = _EVAL_84 | _EVAL_4;
  assign _EVAL_22 = _EVAL_218 | _EVAL_309;
  assign _EVAL_308 = _EVAL_329[17:0];
  assign _EVAL_167 = ~_EVAL_349;
  assign _EVAL_192 = _EVAL_287 | _EVAL_4;
  assign _EVAL_229 = _EVAL_359 == 2'h0;
  assign _EVAL_178 = ~_EVAL_291;
  assign _EVAL_337 = _EVAL_327 | _EVAL_4;
  assign _EVAL_270 = _EVAL_156 & _EVAL_185;
  assign _EVAL_152 = _EVAL_17 == 5'h10;
  assign _EVAL_241 = {1'b0,$signed(_EVAL_236)};
  assign _EVAL_133 = _EVAL_14 & _EVAL_10;
  assign _EVAL_323 = ~_EVAL_165;
  assign _EVAL_176 = _EVAL_10 & _EVAL_83;
  assign _EVAL_254 = ~_EVAL_75;
  assign _EVAL_211 = _EVAL_23[1];
  assign _EVAL_48 = _EVAL_318 | _EVAL_267;
  assign _EVAL_64 = _EVAL_280 | _EVAL_267;
  assign _EVAL_215 = _EVAL_10 & _EVAL_212;
  assign _EVAL_347 = ~_EVAL_25;
  assign _EVAL_141 = 4'h6 == _EVAL;
  assign _EVAL_79 = _EVAL_17 == 5'h8;
  assign _EVAL_265 = _EVAL_1 == 2'h0;
  assign _EVAL_371 = _EVAL_0 & _EVAL_51;
  assign _EVAL_43 = _EVAL_129 - 6'h1;
  assign _EVAL_195 = _EVAL_0 & _EVAL_184;
  assign _EVAL_168 = _EVAL_13 & _EVAL_132;
  assign _EVAL_344 = _EVAL_10 & _EVAL_377;
  assign _EVAL_170 = _EVAL_204 | _EVAL_55;
  assign _EVAL_275 = _EVAL_104 | _EVAL_4;
  assign _EVAL_332 = _EVAL_22 | _EVAL_79;
  assign _EVAL_125 = _EVAL_298 | _EVAL_4;
  assign _EVAL_237 = ~_EVAL_301;
  assign _EVAL_281 = _EVAL_7 <= 3'h1;
  assign _EVAL_284 = _EVAL_86 | _EVAL_4;
  assign _EVAL_217 = _EVAL_101 | _EVAL_4;
  assign _EVAL_53 = _EVAL_0 & _EVAL_324;
  assign _EVAL_305 = $signed(_EVAL_241) & -33'sh1000;
  assign _EVAL_298 = ~_EVAL_3;
  assign _EVAL_287 = _EVAL_1 <= 2'h2;
  assign _EVAL_19 = $signed(_EVAL_34) & -33'sh10000;
  assign _EVAL_90 = _EVAL_76 & _EVAL_93;
  assign _EVAL_196 = _EVAL_277 & _EVAL_64;
  assign _EVAL_39 = ~_EVAL_46;
  assign _EVAL_162 = _EVAL_150 == 6'h0;
  assign _EVAL_71 = _EVAL_12 == 3'h4;
  assign _EVAL_224 = _EVAL_110 == 4'h0;
  assign _EVAL_115 = _EVAL_17 == 5'h11;
  assign _EVAL_291 = _EVAL_59 | _EVAL_4;
  assign _EVAL_184 = _EVAL_12 == 3'h6;
  assign _EVAL_321 = _EVAL_228 | _EVAL_142;
  assign _EVAL_166 = _EVAL_133 & _EVAL_25;
  assign _EVAL_55 = _EVAL_141 & _EVAL_79;
  assign _EVAL_36 = _EVAL_116 & _EVAL_309;
  assign _EVAL_218 = _EVAL_115 | _EVAL_152;
  assign _EVAL_87 = _EVAL_5 == _EVAL_182;
  assign _EVAL_106 = _EVAL_10 & _EVAL_197;
  assign _EVAL_334 = _EVAL_91 & _EVAL_193;
  assign _EVAL_263 = _EVAL_332 | _EVAL_4;
  assign _EVAL_362 = _EVAL_73 | _EVAL_4;
  assign _EVAL_283 = _EVAL_330 | _EVAL_346;
  assign _EVAL_318 = _EVAL_219 | _EVAL_88;
  assign _EVAL_160 = _EVAL_19;
  assign _EVAL_103 = ~_EVAL_316;
  assign _EVAL_159 = _EVAL_276 & _EVAL_152;
  assign _EVAL_304 = _EVAL_5 ^ 32'hc000000;
  assign _EVAL_107 = _EVAL_6 == 5'h8;
  assign _EVAL_52 = _EVAL_41[17:0];
  assign _EVAL_342 = _EVAL_258 + 32'h1;
  assign _EVAL_341 = ~_EVAL_343;
  assign _EVAL_161 = _EVAL_3 == _EVAL_35;
  assign _EVAL_289 = _EVAL_368[7:2];
  assign _EVAL_105 = _EVAL_70 == 2'h0;
  assign _EVAL_28 = ~_EVAL_264;
  assign _EVAL_68 = _EVAL_120 | _EVAL_121;
  assign _EVAL_239 = _EVAL_10 & _EVAL_81;
  assign _EVAL_197 = _EVAL_2 == 3'h7;
  assign _EVAL_122 = _EVAL_288 | _EVAL_4;
  assign _EVAL_200 = _EVAL_62[5:0];
  assign _EVAL_139 = _EVAL_355 | _EVAL_4;
  assign _EVAL_144 = _EVAL_129 == 6'h0;
  assign _EVAL_324 = ~_EVAL_144;
  assign _EVAL_232 = _EVAL_1 == _EVAL_245;
  assign _EVAL_119 = _EVAL_5 ^ 32'h2000000;
  assign _EVAL_235 = _EVAL_340 & _EVAL_256;
  assign _EVAL_357 = _EVAL_342[31:0];
  assign _EVAL_21 = ~_EVAL_63;
  assign _EVAL_149 = _EVAL_87 | _EVAL_4;
  assign _EVAL_248 = _EVAL_268 | _EVAL_27;
  assign _EVAL_290 = _EVAL_12 == 3'h1;
  assign _EVAL_124 = {1'b0,$signed(_EVAL_5)};
  assign _EVAL_314 = ~_EVAL_158;
  assign _EVAL_134 = ~_EVAL_131;
  assign _EVAL_367 = _EVAL_23[0];
  assign _EVAL_24 = 32'h1 << _EVAL_17;
  assign _EVAL_118 = $signed(_EVAL_160) == 33'sh0;
  assign _EVAL_366 = ~_EVAL_217;
  assign _EVAL_359 = _EVAL_6[4:3];
  assign _EVAL_296 = _EVAL_250 | _EVAL_4;
  assign _EVAL_111 = _EVAL_373 | _EVAL_4;
  assign _EVAL_210 = _EVAL_7 == 3'h0;
  assign _EVAL_123 = _EVAL_10 & _EVAL_216;
  assign _EVAL_312 = ~_EVAL_199;
  assign _EVAL_209 = _EVAL_138 | _EVAL_4;
  assign _EVAL_201 = _EVAL >= 4'h2;
  assign _EVAL_262 = _EVAL_91 & _EVAL_256;
  assign _EVAL_310 = _EVAL_6 == 5'h10;
  assign _EVAL_135 = $signed(_EVAL_60) & -33'sh2000;
  assign _EVAL_343 = _EVAL_265 | _EVAL_4;
  assign _EVAL_373 = _EVAL_227 | _EVAL_107;
  assign _EVAL_372 = _EVAL_305;
  assign _EVAL_355 = _EVAL_270 | _EVAL_307;
  assign _EVAL_273 = _EVAL_18 & _EVAL_0;
  assign _EVAL_246 = _EVAL_376 | _EVAL_121;
  assign _EVAL_360 = $signed(_EVAL_299) & -33'sh4000;
  assign _EVAL_252 = ~_EVAL_125;
  assign _EVAL_84 = _EVAL_168 == 4'h0;
  assign _EVAL_186 = _EVAL_268 | _EVAL_29;
  assign _EVAL_319 = _EVAL[0];
  assign _EVAL_143 = _EVAL <= 4'h2;
  assign _EVAL_208 = _EVAL_210 | _EVAL_4;
  assign _EVAL_193 = ~_EVAL_256;
  assign _EVAL_214 = ~_EVAL_326;
  assign _EVAL_112 = _EVAL_281 | _EVAL_4;
  assign _EVAL_30 = _EVAL_9 == _EVAL_89;
  assign _EVAL_146 = _EVAL_295[5:0];
  assign _EVAL_128 = _EVAL_66 | _EVAL_4;
  assign _EVAL_307 = _EVAL_277 & _EVAL_358;
  assign _EVAL_300 = ~_EVAL_128;
  assign _EVAL_181 = _EVAL_12 <= 3'h6;
  assign _EVAL_188 = _EVAL_0 & _EVAL_97;
  assign _EVAL_326 = _EVAL_136 | _EVAL_4;
  assign _EVAL_174 = ~_EVAL_40;
  assign _EVAL_27 = _EVAL_367 & _EVAL_72;
  assign _EVAL_354 = ~_EVAL_208;
  assign _EVAL_74 = ~_EVAL_203;
  assign _EVAL_26 = _EVAL_5 ^ 32'h20000000;
  assign _EVAL_330 = _EVAL_308 != _EVAL_52;
  assign _EVAL_207 = _EVAL_181 | _EVAL_4;
  assign _EVAL_101 = _EVAL_9 >= 4'h2;
  assign _EVAL_240 = {1'b0,$signed(_EVAL_304)};
  assign _EVAL_375 = _EVAL_2[2];
  assign _EVAL_202 = _EVAL == _EVAL_231;
  assign _EVAL_325 = _EVAL_143 & _EVAL_48;
  assign _EVAL_51 = _EVAL_12 == 3'h0;
  assign _EVAL_78 = _EVAL_1 != 2'h2;
  assign _EVAL_225 = ~_EVAL_139;
  assign _EVAL_276 = _EVAL <= 4'hb;
  assign _EVAL_377 = _EVAL_2 == 3'h1;
  assign _EVAL_351 = _EVAL_30 | _EVAL_4;
  assign _EVAL_216 = _EVAL_2 == 3'h3;
  assign _EVAL_83 = _EVAL_2 == 3'h4;
  assign _EVAL_108 = _EVAL_338 >> _EVAL_6;
  assign _EVAL_155 = _EVAL_0 & _EVAL_290;
  assign _EVAL_81 = _EVAL_2 == 3'h6;
  assign _EVAL_299 = {1'b0,$signed(_EVAL_100)};
  assign _EVAL_116 = 4'h2 == _EVAL;
  assign _EVAL_82 = _EVAL_175 | _EVAL_310;
  assign _EVAL_120 = $signed(_EVAL_243) == 33'sh0;
  assign _EVAL_153 = _EVAL_297[5:0];
  assign _EVAL_99 = _EVAL_43[5:0];
  assign _EVAL_346 = ~_EVAL_126;
  assign _EVAL_313 = ~_EVAL_272;
  assign _EVAL_336 = ~_EVAL_16;
  assign _EVAL_340 = ~_EVAL_91;
  assign _EVAL_376 = _EVAL_120 | _EVAL_185;
  assign _EVAL_164 = _EVAL_283 | _EVAL_4;
  assign _EVAL_32 = _EVAL_204 & _EVAL_355;
  assign _EVAL_57 = {_EVAL_321,_EVAL_191,_EVAL_186,_EVAL_248};
  assign _EVAL_271 = _EVAL_7 <= 3'h4;
  assign _EVAL_95 = _EVAL_10 & _EVAL_347;
  assign _EVAL_238 = _EVAL_2 == 3'h0;
  assign _EVAL_180 = _EVAL_246 | _EVAL_118;
  assign _EVAL_309 = _EVAL_105 & _EVAL_365;
  assign _EVAL_356 = ~_EVAL_122;
  assign _EVAL_40 = _EVAL_232 | _EVAL_4;
  assign _EVAL_317 = ~_EVAL_209;
  assign _EVAL_349 = _EVAL_345 | _EVAL_4;
  assign _EVAL_250 = _EVAL_17 == _EVAL_31;
  assign _EVAL_288 = _EVAL_2 == _EVAL_279;
  assign _EVAL_365 = _EVAL_247 <= 3'h6;
  assign _EVAL_297 = _EVAL_249 - 6'h1;
  assign _EVAL_130 = _EVAL_135;
  assign _EVAL_69 = _EVAL_206 | _EVAL_4;
  assign _EVAL_274 = _EVAL_161 | _EVAL_4;
  assign _EVAL_138 = _EVAL_255 == 32'h0;
  assign _EVAL_358 = _EVAL_171 | _EVAL_267;
  assign _EVAL_220 = ~_EVAL_296;
  assign _EVAL_303 = _EVAL_12 == 3'h2;
  assign _EVAL_187 = _EVAL_2 == 3'h5;
  assign _EVAL_76 = _EVAL_273 & _EVAL_109;
  assign _EVAL_42 = ~_EVAL_149;
  assign _EVAL_156 = _EVAL <= 4'h8;
  assign _EVAL_264 = _EVAL_170 | _EVAL_4;
  assign _EVAL_261 = _EVAL_115 | _EVAL_309;
  assign _EVAL_171 = _EVAL_280 | _EVAL_88;
  assign _EVAL_73 = _EVAL_36 & _EVAL_325;
  assign _EVAL_60 = {1'b0,$signed(_EVAL_26)};
  assign _EVAL_56 = _EVAL_5 ^ 32'h1800000;
  assign _EVAL_236 = _EVAL_5 ^ 32'h3000;
  assign _EVAL_34 = {1'b0,$signed(_EVAL_119)};
  assign _EVAL_172 = $signed(_EVAL_269) & -33'sh4000;
  assign _EVAL_47 = _EVAL_273 & _EVAL_144;
  assign _EVAL_80 = _EVAL_8 == _EVAL_350;
  assign _EVAL_222 = _EVAL_68 | _EVAL_118;
  assign _EVAL_212 = _EVAL_2 == 3'h2;
  assign _EVAL_285 = _EVAL_12[0];
  assign _EVAL_280 = _EVAL_222 | _EVAL_293;
  assign _EVAL_315 = _EVAL_147 <= 3'h6;
  assign _EVAL_117 = _EVAL_65 & _EVAL_140;
  assign _EVAL_25 = _EVAL_249 == 6'h0;
  assign _EVAL_374 = _EVAL_172;
  assign _EVAL_62 = _EVAL_150 - 6'h1;
  assign _EVAL_260 = _EVAL_211 & _EVAL_91;
  assign _EVAL_277 = _EVAL <= 4'h6;
  assign _EVAL_142 = _EVAL_367 & _EVAL_262;
  assign _EVAL_94 = ~_EVAL_192;
  assign _EVAL_183 = _EVAL_143 & _EVAL_261;
  assign _EVAL_86 = _EVAL_7 == _EVAL_44;
  assign _EVAL_329 = _EVAL_157 ? _EVAL_24 : 32'h0;
  assign _EVAL_97 = _EVAL_12 == 3'h5;
  assign _EVAL_206 = _EVAL_331 | _EVAL_148;
  assign _EVAL_93 = ~_EVAL_184;
  assign _EVAL_75 = _EVAL_78 | _EVAL_4;
  assign _EVAL_140 = ~_EVAL_52;
  assign _EVAL_33 = _EVAL_270 | _EVAL_333;
  assign _EVAL_66 = _EVAL_298 | _EVAL_16;
  assign _EVAL_361 = ~_EVAL_194;
  assign _EVAL_269 = {1'b0,$signed(_EVAL_56)};
  assign _EVAL_113 = ~_EVAL_351;
  assign _EVAL_145 = ~_EVAL_207;
  assign _EVAL_191 = _EVAL_228 | _EVAL_259;
  assign _EVAL_50 = $signed(_EVAL_240) & -33'sh400000;
  assign _EVAL_226 = _EVAL_223 | _EVAL_4;
  assign _EVAL_243 = _EVAL_173;
  assign _EVAL_327 = ~_EVAL_251;
  assign _EVAL_311 = _EVAL_339[7:0];
  assign _EVAL_251 = _EVAL_221[0];
  assign _EVAL_247 = _EVAL_17[2:0];
  assign _EVAL_267 = $signed(_EVAL_37) == 33'sh0;
  assign _EVAL_132 = ~_EVAL_57;
  assign _EVAL_109 = _EVAL_278 == 6'h0;
  assign _EVAL_286 = ~_EVAL_362;
  assign _EVAL_41 = _EVAL_90 ? _EVAL_154 : 32'h0;
  assign _EVAL_199 = _EVAL_102 | _EVAL_4;
  assign _EVAL_77 = ~_EVAL_11;
  assign _EVAL_126 = |_EVAL_308;
  assign _EVAL_38 = _EVAL_0 & _EVAL_71;
  assign _EVAL_233 = _EVAL_10 & _EVAL_238;
  assign _EVAL_91 = _EVAL_5[1];
  assign _EVAL_316 = _EVAL_336 | _EVAL_4;
  assign _EVAL_219 = _EVAL_180 | _EVAL_293;
  assign _EVAL_266 = ~_EVAL_112;
  assign _EVAL_253 = ~_EVAL_375;
  assign _EVAL_198 = _EVAL_133 | _EVAL_273;
  assign _EVAL_158 = _EVAL_189 | _EVAL_4;
  assign _EVAL_173 = $signed(_EVAL_124) & -33'sh5000;
  assign _EVAL_131 = _EVAL_201 | _EVAL_4;
  assign _EVAL_157 = _EVAL_133 & _EVAL_162;
  assign _EVAL_46 = _EVAL_369 | _EVAL_4;
  assign _EVAL_72 = _EVAL_340 & _EVAL_193;
  assign _EVAL_65 = _EVAL_257 | _EVAL_308;
  assign _EVAL_127 = plusarg_reader_out == 32'h0;
  assign _EVAL_338 = _EVAL_308 | _EVAL_257;
  assign _EVAL_137 = ~_EVAL_275;
  assign _EVAL_223 = _EVAL_270 | _EVAL_196;
  assign _EVAL_96 = ~_EVAL_274;
  assign _EVAL_322 = _EVAL_211 & _EVAL_340;
  assign _EVAL_100 = _EVAL_5 ^ 32'h80000000;
  assign _EVAL_59 = _EVAL_7 <= 3'h3;
  assign _EVAL_335 = ~_EVAL_20;
  assign _EVAL_294 = _EVAL_80 | _EVAL_4;
  assign _EVAL_121 = $signed(_EVAL_374) == 33'sh0;
  assign _EVAL_306 = ~_EVAL_226;
  assign _EVAL_348 = ~_EVAL_263;
  assign _EVAL_221 = _EVAL_257 >> _EVAL_17;
  assign _EVAL_179 = _EVAL_10 & _EVAL_187;
  assign _EVAL_148 = _EVAL_258 < plusarg_reader_out;
  assign _EVAL_175 = _EVAL_6 == 5'h11;
  assign _EVAL_364 = _EVAL_302[7:2];
  assign _EVAL_23 = _EVAL_151 | 2'h1;
  assign _EVAL_272 = _EVAL_32 | _EVAL_4;
  assign _EVAL_85 = ~_EVAL_337;
  assign _EVAL_203 = _EVAL_271 | _EVAL_4;
  assign _EVAL_301 = |_EVAL_257;
  assign _EVAL_345 = _EVAL_7 <= 3'h2;
  assign _EVAL_70 = _EVAL_17[4:3];
  assign _EVAL_88 = $signed(_EVAL_130) == 33'sh0;
  assign _EVAL_295 = _EVAL_278 - 6'h1;
  assign _EVAL_242 = _EVAL_0 & _EVAL_303;
  assign _EVAL_369 = _EVAL_6 == _EVAL_163;
  assign _EVAL_92 = ~_EVAL_4;
  assign _EVAL_227 = _EVAL_82 | _EVAL_353;
  assign _EVAL_352 = ~_EVAL_284;
  assign _EVAL_256 = _EVAL_5[0];
  assign _EVAL_185 = $signed(_EVAL_372) == 33'sh0;
  assign _EVAL_61 = ~_EVAL_111;
  assign _EVAL_189 = _EVAL_108[0];
  assign _EVAL_102 = _EVAL_13 == _EVAL_57;
  assign _EVAL_154 = 32'h1 << _EVAL_6;
  assign _EVAL_147 = _EVAL_6[2:0];
  assign _EVAL_54 = 23'hff << _EVAL_9;
  assign _EVAL_228 = _EVAL_201 | _EVAL_260;
  assign _EVAL_282 = ~_EVAL_164;
  assign _EVAL_58 = _EVAL_54[7:0];
  assign _EVAL_331 = _EVAL_237 | _EVAL_127;
  assign _EVAL_136 = _EVAL_7 != 3'h0;
  assign _EVAL_29 = _EVAL_367 & _EVAL_235;
  assign _EVAL_204 = _EVAL_183 | _EVAL_159;
  always @(posedge _EVAL_15) begin
    if (_EVAL_166) begin
      _EVAL_31 <= _EVAL_17;
    end
    if (_EVAL_47) begin
      _EVAL_35 <= _EVAL_3;
    end
    if (_EVAL_166) begin
      _EVAL_44 <= _EVAL_7;
    end
    if (_EVAL_47) begin
      _EVAL_89 <= _EVAL_9;
    end
    if (_EVAL_4) begin
      _EVAL_129 <= 6'h0;
    end else if (_EVAL_273) begin
      if (_EVAL_144) begin
        if (_EVAL_285) begin
          _EVAL_129 <= _EVAL_289;
        end else begin
          _EVAL_129 <= 6'h0;
        end
      end else begin
        _EVAL_129 <= _EVAL_99;
      end
    end
    if (_EVAL_4) begin
      _EVAL_150 <= 6'h0;
    end else if (_EVAL_133) begin
      if (_EVAL_162) begin
        if (_EVAL_253) begin
          _EVAL_150 <= _EVAL_364;
        end else begin
          _EVAL_150 <= 6'h0;
        end
      end else begin
        _EVAL_150 <= _EVAL_200;
      end
    end
    if (_EVAL_47) begin
      _EVAL_163 <= _EVAL_6;
    end
    if (_EVAL_166) begin
      _EVAL_182 <= _EVAL_5;
    end
    if (_EVAL_47) begin
      _EVAL_213 <= _EVAL_12;
    end
    if (_EVAL_166) begin
      _EVAL_231 <= _EVAL;
    end
    if (_EVAL_47) begin
      _EVAL_245 <= _EVAL_1;
    end
    if (_EVAL_4) begin
      _EVAL_249 <= 6'h0;
    end else if (_EVAL_133) begin
      if (_EVAL_25) begin
        if (_EVAL_253) begin
          _EVAL_249 <= _EVAL_364;
        end else begin
          _EVAL_249 <= 6'h0;
        end
      end else begin
        _EVAL_249 <= _EVAL_153;
      end
    end
    if (_EVAL_4) begin
      _EVAL_257 <= 18'h0;
    end else begin
      _EVAL_257 <= _EVAL_117;
    end
    if (_EVAL_4) begin
      _EVAL_258 <= 32'h0;
    end else if (_EVAL_198) begin
      _EVAL_258 <= 32'h0;
    end else begin
      _EVAL_258 <= _EVAL_357;
    end
    if (_EVAL_4) begin
      _EVAL_278 <= 6'h0;
    end else if (_EVAL_273) begin
      if (_EVAL_109) begin
        if (_EVAL_285) begin
          _EVAL_278 <= _EVAL_289;
        end else begin
          _EVAL_278 <= 6'h0;
        end
      end else begin
        _EVAL_278 <= _EVAL_146;
      end
    end
    if (_EVAL_166) begin
      _EVAL_279 <= _EVAL_2;
    end
    if (_EVAL_47) begin
      _EVAL_350 <= _EVAL_8;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_335) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb49beeb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d3a0b43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_300) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ac0623)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_317) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_306) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_370) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29d88919)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_356) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af688b14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_317) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6619f61)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_366) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e92700d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_361) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da070992)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_348) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(161e83c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(934ffa84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_317) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f56b7a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_317) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e53ecede)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(903717fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_352) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9cc76c87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_323) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d78b4056)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_335) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a260b4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a6025e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_341) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_361) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_341) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46a028de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_348) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16f8204b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dac604b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_352) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d06ad17f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_313) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_145) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c0924d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_300) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ade3567)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe452372)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_371 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74acd6ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_348) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(103de570)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a83c4ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69de435c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_317) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_348) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f67f106)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32f0416b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_370) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_314) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93b396df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_354) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4323ef5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_371 & _EVAL_341) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(523a0e4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_348) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f20f8b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_348) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_356) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_341) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9122d124)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_341) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34b24952)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_335) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_348) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_366) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b881dfc7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_348) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_317) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acf2bd79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_317) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_366) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14b53465)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_354) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19aae2ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_341) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5fc0726)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bde244b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_348) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70233777)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c868be6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_348) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c005f2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_317) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d359d25)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_348) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec2deee8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_361) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_348) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_354) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(221e0179)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30b86fc8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e85e45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_371 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_317) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4397085b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_348) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77dc52db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_74) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88098565)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0d97a18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7621b2f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a310a0f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_317) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_335) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_348) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a723bfd8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_371 & _EVAL_341) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9892362b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7607dc35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_306) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7de5edc9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0666687)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_335) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_317) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4bb7c3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae2d5206)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_348) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(210d7e6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89ee33b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41956d35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd3284dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_335) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(120c0fd0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_74) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(537e132e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91b07483)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_317) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60646166)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_348) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbdeffbe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d60c8d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_314) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_317) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_366) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0061540)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_317) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_313) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75433748)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40bf5fc1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(415683ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_300) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c81eb35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_317) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c2caa6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_354) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b511d979)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_354) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_366) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63e4db9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(375e55b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7621b2f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_341) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63d3852f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_335) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff65f95f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_317) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c2c873f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53957f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a941cbb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0cda94)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_366) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_195 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(facefae1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_371 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_354) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_335) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c7a0665)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_361) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2544680)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_323) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_300) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(931950f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_371 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d03d56f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_31 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_35 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_44 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_89 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_129 = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_150 = _RAND_5[5:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_163 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_182 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_213 = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_231 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_245 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_249 = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_257 = _RAND_12[17:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_258 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_278 = _RAND_14[5:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_279 = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_350 = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
