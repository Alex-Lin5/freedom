//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_162(
  output [31:0] _EVAL,
  input  [8:0]  _EVAL_0,
  output [2:0]  _EVAL_1,
  output [2:0]  _EVAL_2,
  output        _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [31:0] _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  output        _EVAL_10,
  input  [2:0]  _EVAL_11,
  input         _EVAL_12,
  output        _EVAL_13,
  output [1:0]  _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input  [1:0]  _EVAL_17,
  input  [2:0]  _EVAL_18,
  output        _EVAL_19,
  input         _EVAL_20,
  input  [1:0]  _EVAL_21,
  input  [31:0] _EVAL_22,
  output        _EVAL_23,
  output [31:0] _EVAL_24,
  output [8:0]  _EVAL_25,
  output        _EVAL_26,
  output        _EVAL_27,
  output [1:0]  _EVAL_28,
  input         _EVAL_29,
  input         _EVAL_30
);
  wire [2:0] error__EVAL;
  wire  error__EVAL_0;
  wire [127:0] error__EVAL_1;
  wire  error__EVAL_2;
  wire  error__EVAL_3;
  wire [2:0] error__EVAL_4;
  wire  error__EVAL_5;
  wire  error__EVAL_6;
  wire  error__EVAL_7;
  wire  error__EVAL_8;
  wire [31:0] bar__EVAL;
  wire  bar__EVAL_0;
  wire  bar__EVAL_1;
  wire [8:0] bar__EVAL_2;
  wire  bar__EVAL_3;
  wire [2:0] bar__EVAL_4;
  wire  bar__EVAL_5;
  wire  bar__EVAL_6;
  wire  bar__EVAL_7;
  wire  bar__EVAL_8;
  wire  bar__EVAL_9;
  wire [8:0] bar__EVAL_10;
  wire  bar__EVAL_11;
  wire [127:0] bar__EVAL_12;
  wire [2:0] bar__EVAL_13;
  wire [2:0] bar__EVAL_14;
  wire [1:0] bar__EVAL_15;
  wire [31:0] bar__EVAL_16;
  wire [31:0] bar__EVAL_17;
  wire  bar__EVAL_18;
  wire  bar__EVAL_19;
  wire  bar__EVAL_20;
  wire [31:0] bar__EVAL_21;
  wire  bar__EVAL_22;
  wire [2:0] bar__EVAL_23;
  wire [1:0] bar__EVAL_24;
  wire  bar__EVAL_25;
  wire  bar__EVAL_26;
  wire  bar__EVAL_27;
  wire  bar__EVAL_28;
  wire  bar__EVAL_29;
  wire  bar__EVAL_30;
  wire [2:0] bar__EVAL_31;
  wire  bar__EVAL_32;
  wire  bar__EVAL_33;
  wire [2:0] bar__EVAL_34;
  wire  bar__EVAL_35;
  wire [1:0] bar__EVAL_36;
  wire  bar__EVAL_37;
  wire [1:0] bar__EVAL_38;
  _EVAL_161 error (
    ._EVAL(error__EVAL),
    ._EVAL_0(error__EVAL_0),
    ._EVAL_1(error__EVAL_1),
    ._EVAL_2(error__EVAL_2),
    ._EVAL_3(error__EVAL_3),
    ._EVAL_4(error__EVAL_4),
    ._EVAL_5(error__EVAL_5),
    ._EVAL_6(error__EVAL_6),
    ._EVAL_7(error__EVAL_7),
    ._EVAL_8(error__EVAL_8)
  );
  _EVAL_159 bar (
    ._EVAL(bar__EVAL),
    ._EVAL_0(bar__EVAL_0),
    ._EVAL_1(bar__EVAL_1),
    ._EVAL_2(bar__EVAL_2),
    ._EVAL_3(bar__EVAL_3),
    ._EVAL_4(bar__EVAL_4),
    ._EVAL_5(bar__EVAL_5),
    ._EVAL_6(bar__EVAL_6),
    ._EVAL_7(bar__EVAL_7),
    ._EVAL_8(bar__EVAL_8),
    ._EVAL_9(bar__EVAL_9),
    ._EVAL_10(bar__EVAL_10),
    ._EVAL_11(bar__EVAL_11),
    ._EVAL_12(bar__EVAL_12),
    ._EVAL_13(bar__EVAL_13),
    ._EVAL_14(bar__EVAL_14),
    ._EVAL_15(bar__EVAL_15),
    ._EVAL_16(bar__EVAL_16),
    ._EVAL_17(bar__EVAL_17),
    ._EVAL_18(bar__EVAL_18),
    ._EVAL_19(bar__EVAL_19),
    ._EVAL_20(bar__EVAL_20),
    ._EVAL_21(bar__EVAL_21),
    ._EVAL_22(bar__EVAL_22),
    ._EVAL_23(bar__EVAL_23),
    ._EVAL_24(bar__EVAL_24),
    ._EVAL_25(bar__EVAL_25),
    ._EVAL_26(bar__EVAL_26),
    ._EVAL_27(bar__EVAL_27),
    ._EVAL_28(bar__EVAL_28),
    ._EVAL_29(bar__EVAL_29),
    ._EVAL_30(bar__EVAL_30),
    ._EVAL_31(bar__EVAL_31),
    ._EVAL_32(bar__EVAL_32),
    ._EVAL_33(bar__EVAL_33),
    ._EVAL_34(bar__EVAL_34),
    ._EVAL_35(bar__EVAL_35),
    ._EVAL_36(bar__EVAL_36),
    ._EVAL_37(bar__EVAL_37),
    ._EVAL_38(bar__EVAL_38)
  );
  assign error__EVAL_4 = bar__EVAL_31;
  assign bar__EVAL_8 = _EVAL_16;
  assign bar__EVAL_4 = _EVAL_11;
  assign _EVAL_14 = bar__EVAL_38;
  assign error__EVAL_1 = bar__EVAL_12;
  assign _EVAL_19 = bar__EVAL_7;
  assign _EVAL_27 = bar__EVAL_5;
  assign bar__EVAL_10 = _EVAL_0;
  assign bar__EVAL_35 = _EVAL_15;
  assign bar__EVAL_17 = _EVAL_22;
  assign _EVAL_23 = bar__EVAL_26;
  assign _EVAL_13 = bar__EVAL_1;
  assign bar__EVAL_29 = error__EVAL_6;
  assign bar__EVAL_11 = _EVAL_9;
  assign error__EVAL_3 = _EVAL_29;
  assign error__EVAL_0 = _EVAL_16;
  assign bar__EVAL_20 = _EVAL_5;
  assign bar__EVAL_22 = error__EVAL_2;
  assign bar__EVAL_28 = _EVAL_12;
  assign _EVAL_26 = bar__EVAL_32;
  assign _EVAL_10 = bar__EVAL_6;
  assign _EVAL_25 = bar__EVAL_2;
  assign bar__EVAL_14 = _EVAL_18;
  assign bar__EVAL_15 = _EVAL_17;
  assign _EVAL_28 = bar__EVAL_24;
  assign bar__EVAL_33 = _EVAL_29;
  assign bar__EVAL_25 = _EVAL_20;
  assign bar__EVAL_27 = _EVAL_6;
  assign error__EVAL_7 = bar__EVAL_9;
  assign bar__EVAL_19 = error__EVAL_5;
  assign bar__EVAL_36 = _EVAL_21;
  assign _EVAL = bar__EVAL_16;
  assign bar__EVAL_37 = _EVAL_4;
  assign bar__EVAL_18 = _EVAL_30;
  assign _EVAL_2 = bar__EVAL_34;
  assign error__EVAL_8 = bar__EVAL_30;
  assign _EVAL_3 = bar__EVAL_0;
  assign bar__EVAL = _EVAL_7;
  assign _EVAL_24 = bar__EVAL_21;
  assign bar__EVAL_3 = _EVAL_8;
  assign bar__EVAL_13 = error__EVAL;
  assign _EVAL_1 = bar__EVAL_23;
endmodule
