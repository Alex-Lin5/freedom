//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_101_assert(
  input  [3:0]  _EVAL,
  input  [3:0]  _EVAL_0,
  input         _EVAL_1,
  input  [1:0]  _EVAL_2,
  input  [3:0]  _EVAL_3,
  input  [2:0]  _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [2:0]  _EVAL_9,
  input  [31:0] _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input  [2:0]  _EVAL_17,
  input         _EVAL_18
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire [7:0] _EVAL_22;
  reg [3:0] _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire [31:0] _EVAL_27;
  wire [7:0] _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire [32:0] _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire [32:0] _EVAL_41;
  wire [6:0] _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  reg [2:0] _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_52;
  wire [32:0] _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire [32:0] _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire [32:0] _EVAL_62;
  wire [32:0] _EVAL_63;
  wire [31:0] _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire [31:0] _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire [32:0] _EVAL_72;
  wire [5:0] _EVAL_73;
  wire [31:0] _EVAL_74;
  wire  _EVAL_75;
  wire [6:0] _EVAL_77;
  wire  _EVAL_78;
  wire [32:0] _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  reg [2:0] _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire [5:0] _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  reg [5:0] _EVAL_100;
  wire [6:0] _EVAL_101;
  reg [6:0] _EVAL_102;
  wire  _EVAL_103;
  wire [6:0] _EVAL_104;
  wire [31:0] _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire [6:0] _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  reg  _EVAL_111;
  wire  _EVAL_112;
  wire [31:0] _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire [32:0] _EVAL_116;
  wire [32:0] _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire [32:0] _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire [32:0] _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  reg [5:0] _EVAL_129;
  wire  _EVAL_130;
  wire [31:0] _EVAL_131;
  wire [22:0] _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire [5:0] _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire [22:0] _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire [6:0] _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire [3:0] _EVAL_174;
  wire [6:0] _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire [1:0] _EVAL_181;
  wire [7:0] _EVAL_182;
  wire [32:0] _EVAL_183;
  wire  _EVAL_184;
  wire [32:0] _EVAL_185;
  wire [32:0] _EVAL_186;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire [6:0] _EVAL_191;
  wire [7:0] _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire [7:0] _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire [32:0] _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  reg [31:0] _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire [6:0] _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire [3:0] _EVAL_210;
  wire  _EVAL_211;
  reg [2:0] _EVAL_212;
  wire  _EVAL_213;
  wire [31:0] _EVAL_214;
  wire  _EVAL_215;
  wire [31:0] _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  reg [3:0] _EVAL_221;
  wire  _EVAL_222;
  wire [32:0] _EVAL_223;
  wire [3:0] _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire [6:0] _EVAL_228;
  wire [1:0] _EVAL_229;
  wire  _EVAL_230;
  wire [32:0] _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  reg [1:0] _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire [5:0] _EVAL_245;
  reg [31:0] _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire [6:0] _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire [5:0] _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire [7:0] _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_269;
  reg [5:0] _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire [32:0] _EVAL_277;
  reg  _EVAL_278;
  wire [32:0] _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire [5:0] _EVAL_287;
  wire  _EVAL_288;
  wire [32:0] _EVAL_290;
  reg [5:0] _EVAL_291;
  wire  _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_294;
  wire  _EVAL_295;
  wire  _EVAL_296;
  wire [31:0] _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_302;
  wire  _EVAL_303;
  wire [3:0] _EVAL_304;
  wire  _EVAL_305;
  wire [32:0] _EVAL_306;
  wire  _EVAL_307;
  wire  _EVAL_308;
  wire  _EVAL_309;
  wire [7:0] _EVAL_310;
  wire [32:0] _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire [32:0] _EVAL_317;
  wire  _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_320;
  wire [6:0] _EVAL_321;
  wire  _EVAL_322;
  wire  _EVAL_323;
  wire [32:0] _EVAL_324;
  wire  _EVAL_325;
  wire  _EVAL_326;
  wire  _EVAL_327;
  wire  _EVAL_328;
  wire  _EVAL_329;
  wire  _EVAL_330;
  reg [2:0] _EVAL_331;
  wire [7:0] _EVAL_332;
  wire  _EVAL_333;
  wire  _EVAL_334;
  wire  _EVAL_335;
  wire  _EVAL_336;
  wire  _EVAL_337;
  wire  _EVAL_338;
  wire  _EVAL_339;
  wire  _EVAL_340;
  reg [2:0] _EVAL_341;
  wire  _EVAL_342;
  wire  _EVAL_343;
  wire  _EVAL_344;
  wire  _EVAL_345;
  wire  _EVAL_346;
  wire  _EVAL_347;
  wire  _EVAL_348;
  wire  _EVAL_349;
  wire  _EVAL_350;
  wire  _EVAL_351;
  wire  _EVAL_352;
  wire  _EVAL_353;
  wire  _EVAL_354;
  wire  _EVAL_355;
  wire  _EVAL_357;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_149 = _EVAL_89 | _EVAL_1;
  assign _EVAL_173 = _EVAL_12 <= 3'h6;
  assign _EVAL_219 = _EVAL_316 & _EVAL_307;
  assign _EVAL_351 = _EVAL_330 | _EVAL_1;
  assign _EVAL_43 = _EVAL_240 & _EVAL_26;
  assign _EVAL_257 = _EVAL_35 & _EVAL_169;
  assign _EVAL_25 = ~_EVAL_288;
  assign _EVAL_287 = _EVAL_182[7:2];
  assign _EVAL_324 = _EVAL_120;
  assign _EVAL_64 = _EVAL_199[31:0];
  assign _EVAL_333 = _EVAL_16 & _EVAL_8;
  assign _EVAL_27 = _EVAL_10 ^ 32'h3000;
  assign _EVAL_298 = _EVAL_105 == 32'h0;
  assign _EVAL_36 = _EVAL_4 == 3'h1;
  assign _EVAL_231 = $signed(_EVAL_62) & -33'sh4000;
  assign _EVAL_154 = _EVAL_224 == 4'h0;
  assign _EVAL_284 = _EVAL_201 | _EVAL_1;
  assign _EVAL_147 = ~_EVAL_312;
  assign _EVAL_171 = _EVAL_344 | _EVAL_1;
  assign _EVAL_305 = _EVAL[0];
  assign _EVAL_245 = _EVAL_108[5:0];
  assign _EVAL_77 = _EVAL_100 - 6'h1;
  assign _EVAL_315 = _EVAL_9 == 3'h0;
  assign _EVAL_342 = _EVAL_333 & _EVAL_55;
  assign _EVAL_350 = _EVAL_9 == _EVAL_341;
  assign _EVAL_157 = _EVAL_180 & _EVAL_66;
  assign _EVAL_22 = _EVAL_152[7:0];
  assign _EVAL_185 = $signed(_EVAL_223) & -33'sh2000;
  assign _EVAL_52 = _EVAL_7 & _EVAL_34;
  assign _EVAL_327 = _EVAL_130 | _EVAL_1;
  assign _EVAL_259 = _EVAL_195[7:2];
  assign _EVAL_241 = _EVAL_9 <= 3'h1;
  assign _EVAL_229 = 2'h1 << _EVAL_305;
  assign _EVAL_292 = _EVAL_210 == 4'h0;
  assign _EVAL_142 = _EVAL_9 <= 3'h4;
  assign _EVAL_24 = $signed(_EVAL_306) == 33'sh0;
  assign _EVAL_302 = _EVAL_181[1];
  assign _EVAL_58 = $signed(_EVAL_324) == 33'sh0;
  assign _EVAL_45 = 4'h2 == _EVAL;
  assign _EVAL_198 = _EVAL_178 | _EVAL_1;
  assign _EVAL_172 = _EVAL_181[0];
  assign _EVAL_69 = _EVAL_0 == _EVAL_174;
  assign _EVAL_177 = _EVAL_234 | _EVAL_1;
  assign _EVAL_197 = _EVAL_112 | _EVAL_24;
  assign _EVAL_182 = ~_EVAL_22;
  assign _EVAL_155 = _EVAL_7 & _EVAL_49;
  assign _EVAL_258 = _EVAL_226 | _EVAL_188;
  assign _EVAL_248 = _EVAL_315 | _EVAL_1;
  assign _EVAL_299 = ~_EVAL_327;
  assign _EVAL_95 = _EVAL_165[5:0];
  assign _EVAL_332 = 8'h1 << _EVAL_12;
  assign _EVAL_81 = ~_EVAL_6;
  assign _EVAL_153 = _EVAL_344 | _EVAL_18;
  assign _EVAL_290 = {1'b0,$signed(_EVAL_214)};
  assign _EVAL_211 = _EVAL_333 | _EVAL_35;
  assign _EVAL_40 = _EVAL_222 | _EVAL_346;
  assign _EVAL_352 = _EVAL_4 == _EVAL_47;
  assign _EVAL_105 = _EVAL_10 & _EVAL_68;
  assign _EVAL_210 = ~_EVAL_0;
  assign _EVAL_101 = ~_EVAL_249;
  assign _EVAL_319 = _EVAL_241 | _EVAL_1;
  assign _EVAL_99 = ~_EVAL_248;
  assign _EVAL_232 = _EVAL_179 | _EVAL_1;
  assign _EVAL_215 = _EVAL_313 | _EVAL_148;
  assign _EVAL_116 = $signed(_EVAL_311) & -33'sh10000;
  assign _EVAL_63 = _EVAL_116;
  assign _EVAL_165 = _EVAL_291 - 6'h1;
  assign _EVAL_31 = _EVAL_104[0];
  assign _EVAL_328 = ~_EVAL_351;
  assign _EVAL_20 = _EVAL_157 | _EVAL_43;
  assign _EVAL_160 = ~_EVAL_261;
  assign _EVAL_338 = _EVAL_228[0];
  assign _EVAL_34 = _EVAL_4 == 3'h4;
  assign _EVAL_28 = 8'h1 << _EVAL_5;
  assign _EVAL_353 = _EVAL_115 | _EVAL_1;
  assign _EVAL_344 = ~_EVAL_11;
  assign _EVAL_119 = ~_EVAL_284;
  assign _EVAL_307 = ~_EVAL_159;
  assign _EVAL_242 = _EVAL_115 | _EVAL_60;
  assign _EVAL_326 = _EVAL_8 & _EVAL_33;
  assign _EVAL_106 = ~_EVAL_78;
  assign _EVAL_35 = _EVAL_14 & _EVAL_7;
  assign _EVAL_148 = $signed(_EVAL_317) == 33'sh0;
  assign _EVAL_254 = ~_EVAL_218;
  assign _EVAL_300 = _EVAL_65 | _EVAL_1;
  assign _EVAL_295 = ~_EVAL_18;
  assign _EVAL_201 = _EVAL_10 == _EVAL_246;
  assign _EVAL_260 = _EVAL_280 | _EVAL_1;
  assign _EVAL_26 = _EVAL_112 | _EVAL_148;
  assign _EVAL_48 = _EVAL_45 & _EVAL_173;
  assign _EVAL_123 = {1'b0,$signed(_EVAL_10)};
  assign _EVAL_235 = _EVAL_75 | _EVAL_1;
  assign _EVAL_170 = ~_EVAL_83;
  assign _EVAL_216 = _EVAL_10 ^ 32'h80000000;
  assign _EVAL_205 = ~_EVAL_300;
  assign _EVAL_251 = _EVAL_292 | _EVAL_1;
  assign _EVAL_97 = ~_EVAL_252;
  assign _EVAL_127 = _EVAL_17 == 3'h6;
  assign _EVAL_38 = _EVAL_17[2];
  assign _EVAL_223 = {1'b0,$signed(_EVAL_131)};
  assign _EVAL_107 = _EVAL_352 | _EVAL_1;
  assign _EVAL_222 = ~_EVAL_225;
  assign _EVAL_55 = _EVAL_100 == 6'h0;
  assign _EVAL_238 = ~_EVAL_39;
  assign _EVAL_318 = ~_EVAL_336;
  assign _EVAL_152 = 23'hff << _EVAL;
  assign _EVAL_121 = _EVAL_158 | _EVAL_281;
  assign _EVAL_128 = _EVAL_7 & _EVAL_44;
  assign _EVAL_166 = _EVAL_150 & _EVAL_307;
  assign _EVAL_227 = ~_EVAL_151;
  assign _EVAL_56 = _EVAL_17 == _EVAL_212;
  assign _EVAL_271 = ~_EVAL_303;
  assign _EVAL_33 = _EVAL_17 == 3'h1;
  assign _EVAL_311 = {1'b0,$signed(_EVAL_74)};
  assign _EVAL_140 = _EVAL_8 & _EVAL_135;
  assign _EVAL_277 = {1'b0,$signed(_EVAL_27)};
  assign _EVAL_175 = _EVAL_102 | _EVAL_42;
  assign _EVAL_357 = _EVAL_323 | _EVAL_1;
  assign _EVAL_138 = _EVAL_285 | _EVAL_1;
  assign _EVAL_354 = _EVAL_13 == _EVAL_278;
  assign _EVAL_159 = _EVAL_10[0];
  assign _EVAL_110 = ~_EVAL_1;
  assign _EVAL_280 = _EVAL == _EVAL_221;
  assign _EVAL_225 = |_EVAL_102;
  assign _EVAL_325 = ~_EVAL_260;
  assign _EVAL_120 = $signed(_EVAL_72) & -33'sh4000;
  assign _EVAL_334 = ~_EVAL_124;
  assign _EVAL_183 = $signed(_EVAL_123) & -33'sh5000;
  assign _EVAL_94 = _EVAL_196 | _EVAL_1;
  assign _EVAL_228 = _EVAL_102 >> _EVAL_12;
  assign _EVAL_339 = _EVAL_172 & _EVAL_166;
  assign _EVAL_253 = ~_EVAL_349;
  assign _EVAL_234 = _EVAL_2 == _EVAL_239;
  assign _EVAL_169 = _EVAL_291 == 6'h0;
  assign _EVAL_243 = _EVAL_7 & _EVAL_36;
  assign _EVAL_118 = ~_EVAL_177;
  assign _EVAL_158 = _EVAL_57 | _EVAL_293;
  assign _EVAL_194 = ~_EVAL_171;
  assign _EVAL_247 = ~_EVAL_94;
  assign _EVAL_323 = _EVAL_9 <= 3'h2;
  assign _EVAL_282 = _EVAL_17 == 3'h3;
  assign _EVAL_176 = ~_EVAL_90;
  assign _EVAL_237 = _EVAL_172 & _EVAL_217;
  assign _EVAL_60 = _EVAL_302 & _EVAL_150;
  assign _EVAL_276 = _EVAL_5 == _EVAL_331;
  assign _EVAL_320 = _EVAL_7 & _EVAL_122;
  assign _EVAL_230 = ~_EVAL_92;
  assign _EVAL_336 = _EVAL_4 == 3'h6;
  assign _EVAL_264 = _EVAL_24 | _EVAL_46;
  assign _EVAL_202 = _EVAL_3 == _EVAL_23;
  assign _EVAL_80 = _EVAL_172 & _EVAL_213;
  assign _EVAL_181 = _EVAL_229 | 2'h1;
  assign _EVAL_293 = $signed(_EVAL_63) == 33'sh0;
  assign _EVAL_286 = ~_EVAL_38;
  assign _EVAL_322 = _EVAL_333 & _EVAL_218;
  assign _EVAL_355 = _EVAL_5 <= 3'h6;
  assign _EVAL_316 = ~_EVAL_150;
  assign _EVAL_199 = _EVAL_204 + 32'h1;
  assign _EVAL_54 = _EVAL_197 | _EVAL_46;
  assign _EVAL_279 = _EVAL_37;
  assign _EVAL_186 = _EVAL_53;
  assign _EVAL_275 = _EVAL_35 & _EVAL_347;
  assign _EVAL_308 = ~_EVAL_107;
  assign _EVAL_297 = _EVAL_10 ^ 32'hc000000;
  assign _EVAL_348 = _EVAL_143 | _EVAL_293;
  assign _EVAL_163 = ~_EVAL_32;
  assign _EVAL_132 = 23'hff << _EVAL_3;
  assign _EVAL_59 = {1'b0,$signed(_EVAL_297)};
  assign _EVAL_192 = _EVAL_125 ? _EVAL_28 : 8'h0;
  assign _EVAL_68 = {{24'd0}, _EVAL_182};
  assign _EVAL_240 = _EVAL <= 4'h6;
  assign _EVAL_349 = _EVAL_276 | _EVAL_1;
  assign _EVAL_78 = _EVAL_355 | _EVAL_1;
  assign _EVAL_306 = _EVAL_79;
  assign _EVAL_312 = _EVAL_345 | _EVAL_1;
  assign _EVAL_265 = _EVAL_343 & _EVAL_173;
  assign _EVAL_112 = _EVAL_348 | _EVAL_281;
  assign _EVAL_98 = ~_EVAL_198;
  assign _EVAL_236 = ~_EVAL_232;
  assign _EVAL_86 = ~_EVAL_235;
  assign _EVAL_151 = _EVAL_81 | _EVAL_1;
  assign _EVAL_184 = ~_EVAL_294;
  assign _EVAL_53 = $signed(_EVAL_277) & -33'sh1000;
  assign _EVAL_126 = _EVAL_8 & _EVAL_254;
  assign _EVAL_303 = _EVAL_173 | _EVAL_1;
  assign _EVAL_288 = _EVAL_167 | _EVAL_1;
  assign _EVAL_71 = _EVAL_265 | _EVAL_1;
  assign _EVAL_72 = {1'b0,$signed(_EVAL_113)};
  assign _EVAL_65 = _EVAL_3 >= 4'h2;
  assign _EVAL_179 = _EVAL_48 & _EVAL_250;
  assign _EVAL_37 = $signed(_EVAL_59) & -33'sh400000;
  assign _EVAL_218 = _EVAL_129 == 6'h0;
  assign _EVAL_174 = {_EVAL_193,_EVAL_109,_EVAL_91,_EVAL_258};
  assign _EVAL_255 = |_EVAL_42;
  assign _EVAL_50 = _EVAL_17 == 3'h4;
  assign _EVAL_314 = ~_EVAL_272;
  assign _EVAL_217 = _EVAL_316 & _EVAL_159;
  assign _EVAL_161 = _EVAL_8 & _EVAL_282;
  assign _EVAL_83 = _EVAL_208 | _EVAL_1;
  assign _EVAL_301 = _EVAL_17 == 3'h5;
  assign _EVAL_252 = _EVAL_20 | _EVAL_1;
  assign _EVAL_84 = _EVAL_56 | _EVAL_1;
  assign _EVAL_109 = _EVAL_242 | _EVAL_339;
  assign _EVAL_267 = _EVAL_8 & _EVAL_301;
  assign _EVAL_133 = _EVAL_17 == 3'h2;
  assign _EVAL_87 = _EVAL_153 | _EVAL_1;
  assign _EVAL_113 = _EVAL_10 ^ 32'h1800000;
  assign _EVAL_262 = ~_EVAL_61;
  assign _EVAL_91 = _EVAL_226 | _EVAL_237;
  assign _EVAL_296 = _EVAL_8 & _EVAL_50;
  assign _EVAL_62 = {1'b0,$signed(_EVAL_216)};
  assign _EVAL_193 = _EVAL_242 | _EVAL_80;
  assign _EVAL_313 = _EVAL_121 | _EVAL_24;
  assign _EVAL_304 = ~_EVAL_174;
  assign _EVAL_135 = _EVAL_17 == 3'h7;
  assign _EVAL_343 = _EVAL <= 4'h2;
  assign _EVAL_131 = _EVAL_10 ^ 32'h40000000;
  assign _EVAL_213 = _EVAL_150 & _EVAL_159;
  assign _EVAL_309 = _EVAL_329 | _EVAL_1;
  assign _EVAL_330 = _EVAL_11 == _EVAL_111;
  assign _EVAL_283 = _EVAL_7 & _EVAL_336;
  assign _EVAL_114 = ~_EVAL_319;
  assign _EVAL_143 = _EVAL_335 | _EVAL_58;
  assign _EVAL_29 = _EVAL_4[0];
  assign _EVAL_191 = _EVAL_42 | _EVAL_102;
  assign _EVAL_340 = ~_EVAL_357;
  assign _EVAL_195 = ~_EVAL_310;
  assign _EVAL_189 = _EVAL_302 & _EVAL_316;
  assign _EVAL_108 = _EVAL_270 - 6'h1;
  assign _EVAL_226 = _EVAL_115 | _EVAL_189;
  assign _EVAL_200 = ~_EVAL_71;
  assign _EVAL_39 = _EVAL_295 | _EVAL_1;
  assign _EVAL_139 = ~_EVAL_164;
  assign _EVAL_79 = $signed(_EVAL_290) & -33'sh2000;
  assign _EVAL_49 = _EVAL_4 == 3'h0;
  assign _EVAL_32 = _EVAL_350 | _EVAL_1;
  assign _EVAL_104 = _EVAL_191 >> _EVAL_5;
  assign _EVAL_19 = _EVAL_154 | _EVAL_1;
  assign _EVAL_73 = _EVAL_77[5:0];
  assign _EVAL_141 = ~_EVAL_244;
  assign _EVAL_321 = _EVAL_129 - 6'h1;
  assign _EVAL_224 = _EVAL_0 & _EVAL_304;
  assign _EVAL_75 = _EVAL_30 | _EVAL_67;
  assign _EVAL_233 = ~_EVAL_138;
  assign _EVAL_30 = _EVAL_42 != _EVAL_249;
  assign _EVAL_125 = _EVAL_275 & _EVAL_318;
  assign _EVAL_70 = _EVAL_17 == 3'h0;
  assign _EVAL_124 = _EVAL_354 | _EVAL_1;
  assign _EVAL_317 = _EVAL_231;
  assign _EVAL_57 = _EVAL_206 | _EVAL_58;
  assign _EVAL_337 = ~_EVAL_84;
  assign _EVAL_41 = _EVAL_183;
  assign _EVAL_44 = _EVAL_4 == 3'h2;
  assign _EVAL_206 = _EVAL_335 | _EVAL_66;
  assign _EVAL_146 = _EVAL_321[5:0];
  assign _EVAL_220 = _EVAL_8 & _EVAL_70;
  assign _EVAL_250 = _EVAL_343 & _EVAL_215;
  assign _EVAL_214 = _EVAL_10 ^ 32'h20000000;
  assign _EVAL_117 = _EVAL_185;
  assign _EVAL_249 = _EVAL_192[6:0];
  assign _EVAL_207 = _EVAL_175 & _EVAL_101;
  assign _EVAL_188 = _EVAL_172 & _EVAL_219;
  assign _EVAL_335 = $signed(_EVAL_41) == 33'sh0;
  assign _EVAL_244 = _EVAL_137 | _EVAL_1;
  assign _EVAL_256 = _EVAL_2 <= 2'h2;
  assign _EVAL_115 = _EVAL >= 4'h2;
  assign _EVAL_281 = $signed(_EVAL_279) == 33'sh0;
  assign _EVAL_145 = ~_EVAL_19;
  assign _EVAL_310 = _EVAL_132[7:0];
  assign _EVAL_93 = _EVAL_240 & _EVAL_264;
  assign _EVAL_46 = $signed(_EVAL_117) == 33'sh0;
  assign _EVAL_103 = ~_EVAL_87;
  assign _EVAL_329 = _EVAL_2 == 2'h0;
  assign _EVAL_345 = _EVAL_9 <= 3'h3;
  assign _EVAL_66 = $signed(_EVAL_186) == 33'sh0;
  assign _EVAL_190 = _EVAL_4 == 3'h5;
  assign _EVAL_164 = _EVAL_162 | _EVAL_1;
  assign _EVAL_285 = _EVAL_157 | _EVAL_93;
  assign _EVAL_67 = ~_EVAL_255;
  assign _EVAL_272 = _EVAL_256 | _EVAL_1;
  assign _EVAL_96 = _EVAL_54 | _EVAL_148;
  assign _EVAL_346 = plusarg_reader_out == 32'h0;
  assign _EVAL_74 = _EVAL_10 ^ 32'h2000000;
  assign _EVAL_208 = _EVAL_40 | _EVAL_269;
  assign _EVAL_168 = ~_EVAL_149;
  assign _EVAL_90 = _EVAL_202 | _EVAL_1;
  assign _EVAL_261 = _EVAL_69 | _EVAL_1;
  assign _EVAL_294 = _EVAL_31 | _EVAL_1;
  assign _EVAL_89 = ~_EVAL_338;
  assign _EVAL_137 = _EVAL_9 != 3'h0;
  assign _EVAL_162 = _EVAL_2 != 2'h2;
  assign _EVAL_347 = _EVAL_270 == 6'h0;
  assign _EVAL_209 = _EVAL_8 & _EVAL_127;
  assign _EVAL_266 = ~_EVAL_353;
  assign _EVAL_144 = _EVAL_7 & _EVAL_190;
  assign _EVAL_263 = _EVAL_342 ? _EVAL_332 : 8'h0;
  assign _EVAL_130 = _EVAL_265 & _EVAL_178;
  assign _EVAL_42 = _EVAL_263[6:0];
  assign _EVAL_82 = ~_EVAL_251;
  assign _EVAL_180 = _EVAL <= 4'h8;
  assign _EVAL_61 = _EVAL_142 | _EVAL_1;
  assign _EVAL_167 = _EVAL_12 == _EVAL_85;
  assign _EVAL_21 = ~_EVAL_309;
  assign _EVAL_136 = _EVAL_240 & _EVAL_96;
  assign _EVAL_150 = _EVAL_10[1];
  assign _EVAL_203 = _EVAL_8 & _EVAL_133;
  assign _EVAL_122 = ~_EVAL_169;
  assign _EVAL_178 = _EVAL_157 | _EVAL_136;
  assign _EVAL_269 = _EVAL_204 < plusarg_reader_out;
  assign _EVAL_196 = _EVAL_4 <= 3'h6;
  assign _EVAL_92 = _EVAL_298 | _EVAL_1;
  always @(posedge _EVAL_15) begin
    if (_EVAL_257) begin
      _EVAL_23 <= _EVAL_3;
    end
    if (_EVAL_257) begin
      _EVAL_47 <= _EVAL_4;
    end
    if (_EVAL_322) begin
      _EVAL_85 <= _EVAL_12;
    end
    if (_EVAL_1) begin
      _EVAL_100 <= 6'h0;
    end else if (_EVAL_333) begin
      if (_EVAL_55) begin
        if (_EVAL_286) begin
          _EVAL_100 <= _EVAL_287;
        end else begin
          _EVAL_100 <= 6'h0;
        end
      end else begin
        _EVAL_100 <= _EVAL_73;
      end
    end
    if (_EVAL_1) begin
      _EVAL_102 <= 7'h0;
    end else begin
      _EVAL_102 <= _EVAL_207;
    end
    if (_EVAL_257) begin
      _EVAL_111 <= _EVAL_11;
    end
    if (_EVAL_1) begin
      _EVAL_129 <= 6'h0;
    end else if (_EVAL_333) begin
      if (_EVAL_218) begin
        if (_EVAL_286) begin
          _EVAL_129 <= _EVAL_287;
        end else begin
          _EVAL_129 <= 6'h0;
        end
      end else begin
        _EVAL_129 <= _EVAL_146;
      end
    end
    if (_EVAL_1) begin
      _EVAL_204 <= 32'h0;
    end else if (_EVAL_211) begin
      _EVAL_204 <= 32'h0;
    end else begin
      _EVAL_204 <= _EVAL_64;
    end
    if (_EVAL_322) begin
      _EVAL_212 <= _EVAL_17;
    end
    if (_EVAL_322) begin
      _EVAL_221 <= _EVAL;
    end
    if (_EVAL_257) begin
      _EVAL_239 <= _EVAL_2;
    end
    if (_EVAL_322) begin
      _EVAL_246 <= _EVAL_10;
    end
    if (_EVAL_1) begin
      _EVAL_270 <= 6'h0;
    end else if (_EVAL_35) begin
      if (_EVAL_347) begin
        if (_EVAL_29) begin
          _EVAL_270 <= _EVAL_259;
        end else begin
          _EVAL_270 <= 6'h0;
        end
      end else begin
        _EVAL_270 <= _EVAL_245;
      end
    end
    if (_EVAL_257) begin
      _EVAL_278 <= _EVAL_13;
    end
    if (_EVAL_1) begin
      _EVAL_291 <= 6'h0;
    end else if (_EVAL_35) begin
      if (_EVAL_169) begin
        if (_EVAL_29) begin
          _EVAL_291 <= _EVAL_259;
        end else begin
          _EVAL_291 <= 6'h0;
        end
      end else begin
        _EVAL_291 <= _EVAL_95;
      end
    end
    if (_EVAL_257) begin
      _EVAL_331 <= _EVAL_5;
    end
    if (_EVAL_322) begin
      _EVAL_341 <= _EVAL_9;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_99) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6bf469cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_328) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_253) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21001659)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_114) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_340) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(faf18ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_334) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1dafdc70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_7 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_145) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92a61064)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca4826f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e05e9a04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df634f7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_7 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b08e40b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5090a37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ebfc353)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(239bb4d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b65f128f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(136c683e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a301609f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7318577)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_314) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a4b1e77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b4ad127)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(101a5125)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_328) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5fc8c05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_243 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_325) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67a926fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_266) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1671bf40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1d3e2b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8cbdc90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_99) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb97ccfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_314) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4501eb95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ef5f2d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1bb2b4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(615bd548)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9953525e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_334) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f47095f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4bc71dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9b71052)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(930c0471)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a40905bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2aeaf440)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b23d9bd5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_99) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_299) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0b98acd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4e885a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2a93f20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_308) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f49aa13a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(909d2a15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_99) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66a33cf6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(600bf219)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_243 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ef4fe1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fcaaa82e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ddf07c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_337) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_176) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb068aa4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(509a0e0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf278f6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c257b2af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d73b32dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2242e9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95b41ef8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fcd5f5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2adc7244)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2fea48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_340) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9fa1c1c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3987bb92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56d7502c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_299) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5330fec1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_342 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9ff4426)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4185d32a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13d71a9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_253) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_308) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c205bac1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_243 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ce2cd1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_243 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d17f0c38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_340) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1fd20aa1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4915f2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40fb75f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdd6515d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_99) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_340) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32281688)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2360da43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c321ec83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18dfdd2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_230) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f10fcf2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48fbcc88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb6a0b86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_342 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e31bf012)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(172f2ee1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_114) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58de1a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_314) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bfdbe0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2ea0c0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dace447a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_176) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7efc77c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21507fd2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94d0f3e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_325) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c996892)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_326 & _EVAL_99) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efa2678c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_266) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_243 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4832ab6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_243 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9db9dd43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_230) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b40398f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_337) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1625ba1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a4b1e77)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_314) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_23 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_47 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_85 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_100 = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_102 = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_111 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_129 = _RAND_6[5:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_204 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_212 = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_221 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_239 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_246 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_270 = _RAND_12[5:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_278 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_291 = _RAND_14[5:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_331 = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_341 = _RAND_16[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
