//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_95_assert(
  input  [27:0] _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [9:0]  _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [2:0]  _EVAL_4,
  input         _EVAL_5,
  input  [1:0]  _EVAL_6,
  input  [2:0]  _EVAL_7,
  input  [1:0]  _EVAL_8,
  input  [9:0]  _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input  [3:0]  _EVAL_13,
  input         _EVAL_14
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [575:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_15;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire [1:0] _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire [1:0] _EVAL_24;
  reg  _EVAL_25;
  wire [27:0] _EVAL_26;
  wire  _EVAL_27;
  wire [31:0] _EVAL_29;
  wire [1:0] _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  reg [2:0] _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire [575:0] _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire [1023:0] _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire [3:0] _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  reg [1:0] _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire [1:0] _EVAL_69;
  wire [1:0] _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire [575:0] _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire [28:0] _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  reg  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire [27:0] _EVAL_96;
  wire [575:0] _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire [1023:0] _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_109;
  wire [575:0] _EVAL_110;
  wire  _EVAL_111;
  wire [1023:0] _EVAL_112;
  wire  _EVAL_113;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_114;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire [1:0] _EVAL_120;
  wire [575:0] _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  reg [9:0] _EVAL_125;
  reg [31:0] _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  reg [2:0] _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  reg  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  reg [9:0] _EVAL_149;
  wire [4:0] _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire [27:0] _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire [28:0] _EVAL_161;
  wire [3:0] _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  reg [1:0] _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire [575:0] _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire [28:0] _EVAL_177;
  wire  _EVAL_178;
  wire [575:0] _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire [3:0] _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire [1023:0] _EVAL_190;
  reg [575:0] _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire [3:0] _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  reg [2:0] _EVAL_206;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  reg  _EVAL_222;
  reg [27:0] _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire [1:0] _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire [1:0] _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire [575:0] _EVAL_241;
  wire [32:0] _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_47 = ~_EVAL_181;
  assign _EVAL_178 = _EVAL_30[0];
  assign _EVAL_228 = _EVAL_49 | _EVAL_50;
  assign _EVAL_209 = ~_EVAL_151;
  assign _EVAL_130 = _EVAL_44 & _EVAL_134;
  assign _EVAL_101 = _EVAL_224 ? _EVAL_190 : 1024'h0;
  assign _EVAL_91 = _EVAL_4 == 3'h6;
  assign _EVAL_162 = {_EVAL_212,_EVAL_139,_EVAL_228,_EVAL_235};
  assign _EVAL_66 = _EVAL == _EVAL_223;
  assign _EVAL_198 = ~_EVAL_1;
  assign _EVAL_180 = _EVAL_5 & _EVAL_183;
  assign _EVAL_210 = ~_EVAL_182;
  assign _EVAL_144 = _EVAL_215 | _EVAL_1;
  assign _EVAL_61 = ~_EVAL_80;
  assign _EVAL_173 = _EVAL_14 & _EVAL_63;
  assign _EVAL_172 = _EVAL_241[0];
  assign _EVAL_135 = _EVAL_134 & _EVAL_202;
  assign _EVAL_202 = _EVAL[0];
  assign _EVAL_161 = _EVAL_177;
  assign _EVAL_58 = _EVAL_205 | _EVAL_1;
  assign _EVAL_82 = _EVAL_44 & _EVAL_128;
  assign _EVAL_75 = _EVAL_121 | _EVAL_191;
  assign _EVAL_51 = ~_EVAL_98;
  assign _EVAL_165 = ~_EVAL_227;
  assign _EVAL_200 = ~_EVAL_13;
  assign _EVAL_118 = ~_EVAL_202;
  assign _EVAL_211 = _EVAL_7 <= 3'h3;
  assign _EVAL_127 = _EVAL_39[0];
  assign _EVAL_188 = _EVAL_126 < plusarg_reader_out;
  assign _EVAL_218 = ~_EVAL_20;
  assign _EVAL_93 = _EVAL_240 | _EVAL_1;
  assign _EVAL_53 = plusarg_reader_out == 32'h0;
  assign _EVAL_37 = _EVAL_229 | _EVAL_1;
  assign _EVAL_196 = _EVAL_68 | _EVAL_188;
  assign _EVAL_232 = ~_EVAL_222;
  assign _EVAL_65 = ~_EVAL_56;
  assign _EVAL_72 = ~_EVAL_85;
  assign _EVAL_56 = _EVAL_127 | _EVAL_1;
  assign _EVAL_174 = _EVAL_97 & _EVAL_110;
  assign _EVAL_102 = _EVAL_5 & _EVAL_201;
  assign _EVAL_81 = _EVAL_2 == _EVAL_125;
  assign _EVAL_94 = _EVAL_6 <= 2'h2;
  assign _EVAL_15 = _EVAL_4 == 3'h3;
  assign _EVAL_154 = _EVAL_109 & _EVAL_175;
  assign _EVAL_67 = _EVAL_107 | _EVAL_1;
  assign _EVAL_185 = _EVAL_103 | _EVAL_1;
  assign _EVAL_114 = _EVAL_10 & _EVAL_5;
  assign _EVAL_140 = _EVAL_5 & _EVAL_20;
  assign _EVAL_156 = _EVAL_116 | _EVAL_1;
  assign _EVAL_97 = _EVAL_191 | _EVAL_121;
  assign _EVAL_18 = _EVAL_5 & _EVAL_237;
  assign _EVAL_241 = _EVAL_191 >> _EVAL_9;
  assign _EVAL_219 = _EVAL_214 | _EVAL_1;
  assign _EVAL_163 = _EVAL_195 | _EVAL_114;
  assign _EVAL_183 = _EVAL_3 == 3'h4;
  assign _EVAL_234 = ~_EVAL_31;
  assign _EVAL_159 = ~_EVAL_12;
  assign _EVAL_233 = _EVAL_92 - 1'h1;
  assign _EVAL_45 = _EVAL_35 & _EVAL_218;
  assign _EVAL_212 = _EVAL_189 | _EVAL_113;
  assign _EVAL_168 = _EVAL_216 | _EVAL_1;
  assign _EVAL_117 = _EVAL_196 | _EVAL_1;
  assign _EVAL_99 = _EVAL_3 == _EVAL_206;
  assign _EVAL_134 = ~_EVAL_128;
  assign _EVAL_197 = _EVAL_4 == _EVAL_129;
  assign _EVAL_122 = ~_EVAL_171;
  assign _EVAL_78 = {1'b0,$signed(_EVAL_158)};
  assign _EVAL_46 = ~_EVAL_168;
  assign _EVAL_104 = _EVAL_226 & _EVAL_105;
  assign _EVAL_55 = ~_EVAL_138;
  assign _EVAL_128 = _EVAL[1];
  assign _EVAL_84 = _EVAL_99 | _EVAL_1;
  assign _EVAL_184 = _EVAL_13 & _EVAL_52;
  assign _EVAL_171 = _EVAL_159 | _EVAL_1;
  assign _EVAL_76 = _EVAL_195 & _EVAL_80;
  assign _EVAL_112 = 1024'h1 << _EVAL_2;
  assign _EVAL_36 = _EVAL_33 | _EVAL_1;
  assign _EVAL_22 = _EVAL_109 & _EVAL_43;
  assign _EVAL_148 = _EVAL_4 == 3'h1;
  assign _EVAL_31 = _EVAL_66 | _EVAL_1;
  assign _EVAL_194 = _EVAL_2 <= 10'h23f;
  assign _EVAL_24 = _EVAL_19 | 2'h1;
  assign _EVAL_103 = _EVAL_26 == 28'h0;
  assign _EVAL_220 = _EVAL_14 & _EVAL_61;
  assign _EVAL_153 = ~_EVAL_133;
  assign _EVAL_121 = _EVAL_101[575:0];
  assign _EVAL_113 = _EVAL_109 & _EVAL_74;
  assign _EVAL_43 = _EVAL_134 & _EVAL_118;
  assign _EVAL_214 = _EVAL_119 | _EVAL_77;
  assign _EVAL_44 = _EVAL_24[1];
  assign _EVAL_83 = _EVAL_14 & _EVAL_123;
  assign _EVAL_39 = _EVAL_75 >> _EVAL_2;
  assign _EVAL_145 = _EVAL_8 == _EVAL_167;
  assign _EVAL_169 = _EVAL_105 | _EVAL_1;
  assign _EVAL_143 = ~_EVAL_193;
  assign _EVAL_73 = _EVAL_146 | _EVAL_1;
  assign _EVAL_239 = _EVAL_9 == _EVAL_149;
  assign _EVAL_79 = _EVAL_226 | _EVAL_1;
  assign _EVAL_142 = _EVAL_13 == _EVAL_162;
  assign _EVAL_236 = _EVAL_114 & _EVAL_55;
  assign _EVAL_70 = _EVAL_25 - 1'h1;
  assign _EVAL_177 = $signed(_EVAL_78) & -29'sh400000;
  assign _EVAL_151 = _EVAL_211 | _EVAL_1;
  assign _EVAL_96 = {{26'd0}, _EVAL_69};
  assign _EVAL_95 = _EVAL_200 == 4'h0;
  assign _EVAL_227 = |_EVAL_191;
  assign _EVAL_30 = _EVAL_222 - 1'h1;
  assign _EVAL_111 = _EVAL_5 & _EVAL_186;
  assign _EVAL_204 = _EVAL_6[0];
  assign _EVAL_109 = _EVAL_24[0];
  assign _EVAL_195 = _EVAL_11 & _EVAL_14;
  assign _EVAL_199 = ~_EVAL_84;
  assign _EVAL_41 = _EVAL_5 & _EVAL_23;
  assign _EVAL_62 = _EVAL_197 | _EVAL_1;
  assign _EVAL_242 = _EVAL_126 + 32'h1;
  assign _EVAL_50 = _EVAL_109 & _EVAL_135;
  assign _EVAL_85 = _EVAL_239 | _EVAL_1;
  assign _EVAL_19 = 2'h1 << _EVAL_204;
  assign _EVAL_216 = ~_EVAL_172;
  assign _EVAL_217 = ~_EVAL_219;
  assign _EVAL_69 = ~_EVAL_120;
  assign _EVAL_100 = _EVAL_14 & _EVAL_91;
  assign _EVAL_139 = _EVAL_189 | _EVAL_154;
  assign _EVAL_90 = _EVAL_4 == 3'h2;
  assign _EVAL_175 = _EVAL_128 & _EVAL_118;
  assign _EVAL_68 = _EVAL_165 | _EVAL_53;
  assign _EVAL_23 = _EVAL_3 == 3'h0;
  assign _EVAL_54 = _EVAL_14 & _EVAL_15;
  assign _EVAL_244 = ~_EVAL_25;
  assign _EVAL_86 = ~_EVAL_67;
  assign _EVAL_215 = _EVAL_6 == _EVAL_64;
  assign _EVAL_160 = ~_EVAL_79;
  assign _EVAL_170 = _EVAL_233[0];
  assign _EVAL_192 = _EVAL_4 == 3'h7;
  assign _EVAL_40 = ~_EVAL_59;
  assign _EVAL_187 = ~_EVAL_176;
  assign _EVAL_116 = _EVAL_7 != 3'h0;
  assign _EVAL_21 = ~_EVAL_156;
  assign _EVAL_80 = ~_EVAL_92;
  assign _EVAL_164 = ~_EVAL_73;
  assign _EVAL_59 = _EVAL_95 | _EVAL_1;
  assign _EVAL_230 = _EVAL_138 - 1'h1;
  assign _EVAL_181 = _EVAL_145 | _EVAL_1;
  assign _EVAL_88 = _EVAL_14 & _EVAL_148;
  assign _EVAL_33 = _EVAL_8 >= 2'h2;
  assign _EVAL_133 = _EVAL_104 | _EVAL_1;
  assign _EVAL_176 = _EVAL_81 | _EVAL_1;
  assign _EVAL_71 = _EVAL_230[0];
  assign _EVAL_226 = _EVAL_9 <= 10'h23f;
  assign _EVAL_29 = _EVAL_242[31:0];
  assign _EVAL_150 = 5'h3 << _EVAL_6;
  assign _EVAL_120 = _EVAL_150[1:0];
  assign _EVAL_166 = ~_EVAL_37;
  assign _EVAL_231 = _EVAL_221 | _EVAL_1;
  assign _EVAL_235 = _EVAL_49 | _EVAL_22;
  assign _EVAL_146 = _EVAL_3 <= 3'h6;
  assign _EVAL_229 = _EVAL_6 >= 2'h2;
  assign _EVAL_155 = |_EVAL_121;
  assign _EVAL_193 = _EVAL_142 | _EVAL_1;
  assign _EVAL_203 = $signed(_EVAL_161) == 29'sh0;
  assign _EVAL_205 = _EVAL_7 == _EVAL_34;
  assign _EVAL_119 = _EVAL_121 != _EVAL_179;
  assign _EVAL_32 = ~_EVAL_36;
  assign _EVAL_182 = _EVAL_194 | _EVAL_1;
  assign _EVAL_186 = _EVAL_3 == 3'h2;
  assign _EVAL_63 = _EVAL_4 == 3'h5;
  assign _EVAL_38 = _EVAL_137 | _EVAL_1;
  assign _EVAL_208 = _EVAL_70[0];
  assign _EVAL_27 = ~_EVAL_169;
  assign _EVAL_201 = _EVAL_3 == 3'h1;
  assign _EVAL_240 = _EVAL_7 <= 3'h1;
  assign _EVAL_190 = 1024'h1 << _EVAL_9;
  assign _EVAL_110 = ~_EVAL_179;
  assign _EVAL_49 = _EVAL_229 | _EVAL_130;
  assign _EVAL_124 = ~_EVAL_117;
  assign _EVAL_60 = _EVAL_7 <= 3'h4;
  assign _EVAL_137 = _EVAL_184 == 4'h0;
  assign _EVAL_106 = _EVAL_14 & _EVAL_192;
  assign _EVAL_26 = _EVAL & _EVAL_96;
  assign _EVAL_189 = _EVAL_229 | _EVAL_82;
  assign _EVAL_52 = ~_EVAL_162;
  assign _EVAL_147 = _EVAL_14 & _EVAL_136;
  assign _EVAL_98 = _EVAL_60 | _EVAL_1;
  assign _EVAL_238 = _EVAL_5 & _EVAL_57;
  assign _EVAL_20 = _EVAL_3 == 3'h6;
  assign _EVAL_157 = ~_EVAL_93;
  assign _EVAL_57 = _EVAL_3 == 3'h5;
  assign _EVAL_179 = _EVAL_48[575:0];
  assign _EVAL_224 = _EVAL_195 & _EVAL_244;
  assign _EVAL_105 = _EVAL_94 & _EVAL_203;
  assign _EVAL_77 = ~_EVAL_155;
  assign _EVAL_221 = _EVAL_7 == 3'h0;
  assign _EVAL_17 = ~_EVAL_185;
  assign _EVAL_16 = _EVAL_14 & _EVAL_90;
  assign _EVAL_123 = _EVAL_4 == 3'h4;
  assign _EVAL_48 = _EVAL_45 ? _EVAL_112 : 1024'h0;
  assign _EVAL_141 = ~_EVAL_62;
  assign _EVAL_225 = ~_EVAL_38;
  assign _EVAL_158 = _EVAL ^ 28'hc000000;
  assign _EVAL_237 = ~_EVAL_55;
  assign _EVAL_35 = _EVAL_114 & _EVAL_232;
  assign _EVAL_89 = ~_EVAL_231;
  assign _EVAL_107 = _EVAL_7 <= 3'h2;
  assign _EVAL_136 = _EVAL_4 == 3'h0;
  assign _EVAL_213 = ~_EVAL_144;
  assign _EVAL_243 = ~_EVAL_58;
  assign _EVAL_74 = _EVAL_128 & _EVAL_202;
  always @(posedge _EVAL_0) begin
    if (_EVAL_1) begin
      _EVAL_25 <= 1'h0;
    end else if (_EVAL_195) begin
      if (_EVAL_244) begin
        _EVAL_25 <= 1'h0;
      end else begin
        _EVAL_25 <= _EVAL_208;
      end
    end
    if (_EVAL_76) begin
      _EVAL_34 <= _EVAL_7;
    end
    if (_EVAL_76) begin
      _EVAL_64 <= _EVAL_6;
    end
    if (_EVAL_1) begin
      _EVAL_92 <= 1'h0;
    end else if (_EVAL_195) begin
      if (_EVAL_80) begin
        _EVAL_92 <= 1'h0;
      end else begin
        _EVAL_92 <= _EVAL_170;
      end
    end
    if (_EVAL_236) begin
      _EVAL_125 <= _EVAL_2;
    end
    if (_EVAL_1) begin
      _EVAL_126 <= 32'h0;
    end else if (_EVAL_163) begin
      _EVAL_126 <= 32'h0;
    end else begin
      _EVAL_126 <= _EVAL_29;
    end
    if (_EVAL_76) begin
      _EVAL_129 <= _EVAL_4;
    end
    if (_EVAL_1) begin
      _EVAL_138 <= 1'h0;
    end else if (_EVAL_114) begin
      if (_EVAL_55) begin
        _EVAL_138 <= 1'h0;
      end else begin
        _EVAL_138 <= _EVAL_71;
      end
    end
    if (_EVAL_76) begin
      _EVAL_149 <= _EVAL_9;
    end
    if (_EVAL_236) begin
      _EVAL_167 <= _EVAL_8;
    end
    if (_EVAL_1) begin
      _EVAL_191 <= 576'h0;
    end else begin
      _EVAL_191 <= _EVAL_174;
    end
    if (_EVAL_236) begin
      _EVAL_206 <= _EVAL_3;
    end
    if (_EVAL_1) begin
      _EVAL_222 <= 1'h0;
    end else if (_EVAL_114) begin
      if (_EVAL_232) begin
        _EVAL_222 <= 1'h0;
      end else begin
        _EVAL_222 <= _EVAL_178;
      end
    end
    if (_EVAL_76) begin
      _EVAL_223 <= _EVAL;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fba1d34a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f5d0292)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a269a788)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(333cf7c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(298b0a80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dba2cfb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a93fa8d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(83b13d00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55a2ed4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59416da7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(443136d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bf87dd0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3fa24e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f9afd3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6c17ac2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17c7a34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9382678)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff119467)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62985c96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8c8230c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0671c02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5154001e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75458866)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9d11f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34becfc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(adfc3ac2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(478464ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb4bc42a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd25e753)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d403b413)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33bfedc7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30becf39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c588958)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd10db74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2505badf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35214b80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35a72927)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb6ac07a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(142f6ca6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(208679dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d403b413)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8e1798c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae068599)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54849923)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da9d1cdd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4a48f18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e32fc76c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a823a5ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23f521a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3544ad4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ae784e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2521483)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5a4f347)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a33f57e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7aa1724)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90e5af7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9437933a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(662b4a53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0e24ec5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9806a97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_199) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d49b5bb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c42a47bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f1fe8bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_199) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a955a9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(727db7d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_198) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f5e234e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_198) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acc21b26)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b30a19bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_147 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff4effb6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1960e4f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(468b873d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_54 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17ebeb30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f6e7447)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c393cf7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_88 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d8bb28b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_100 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(479a8644)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_25 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_34 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_64 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_92 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_125 = _RAND_4[9:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_126 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_129 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_138 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_149 = _RAND_8[9:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_167 = _RAND_9[1:0];
  _RAND_10 = {18{`RANDOM}};
  _EVAL_191 = _RAND_10[575:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_206 = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_222 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_223 = _RAND_13[27:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
