//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_113(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  output [31:0] _EVAL_2,
  input  [1:0]  _EVAL_3,
  input  [29:0] _EVAL_4,
  input         _EVAL_5,
  input  [31:0] _EVAL_6,
  input         _EVAL_7,
  input  [31:0] _EVAL_8,
  input         _EVAL_9,
  input  [31:0] _EVAL_10,
  input         _EVAL_11,
  output        _EVAL_12,
  input         _EVAL_13,
  input  [31:0] _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18,
  input         _EVAL_19,
  input  [1:0]  _EVAL_20,
  input         _EVAL_21,
  input  [29:0] _EVAL_22,
  input  [1:0]  _EVAL_23,
  input         _EVAL_24,
  input         _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  input  [29:0] _EVAL_30,
  input  [29:0] _EVAL_31,
  input  [1:0]  _EVAL_32,
  input         _EVAL_33,
  input         _EVAL_34,
  input  [31:0] _EVAL_35,
  input  [1:0]  _EVAL_36,
  input  [29:0] _EVAL_37,
  input  [1:0]  _EVAL_38,
  input  [31:0] _EVAL_39,
  input         _EVAL_40,
  input         _EVAL_41,
  input         _EVAL_42,
  input         _EVAL_43,
  input         _EVAL_44,
  input  [31:0] _EVAL_45,
  input         _EVAL_46,
  input  [31:0] _EVAL_47,
  input         _EVAL_48,
  input  [1:0]  _EVAL_49,
  input         _EVAL_50,
  input         _EVAL_51,
  input         _EVAL_52,
  input  [1:0]  _EVAL_53,
  input         _EVAL_54,
  input  [31:0] _EVAL_55,
  input         _EVAL_56,
  input  [1:0]  _EVAL_57,
  input  [29:0] _EVAL_58,
  input         _EVAL_59,
  input  [29:0] _EVAL_60,
  input  [29:0] _EVAL_61
);
  wire  _EVAL_62;
  wire [32:0] _EVAL_63;
  wire [32:0] _EVAL_64;
  wire [32:0] _EVAL_65;
  wire  _EVAL_66;
  wire [32:0] _EVAL_67;
  wire [32:0] _EVAL_68;
  wire  _EVAL_69;
  wire [31:0] _EVAL_70;
  wire [2:0] _EVAL_71;
  wire [32:0] _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire [32:0] _EVAL_76;
  wire  pmp__EVAL;
  wire [31:0] pmp__EVAL_0;
  wire [29:0] pmp__EVAL_1;
  wire  pmp__EVAL_2;
  wire  pmp__EVAL_3;
  wire  pmp__EVAL_4;
  wire [29:0] pmp__EVAL_5;
  wire  pmp__EVAL_6;
  wire [1:0] pmp__EVAL_7;
  wire  pmp__EVAL_8;
  wire  pmp__EVAL_9;
  wire [1:0] pmp__EVAL_10;
  wire [1:0] pmp__EVAL_11;
  wire [1:0] pmp__EVAL_12;
  wire  pmp__EVAL_13;
  wire  pmp__EVAL_14;
  wire  pmp__EVAL_15;
  wire [1:0] pmp__EVAL_16;
  wire  pmp__EVAL_17;
  wire  pmp__EVAL_18;
  wire  pmp__EVAL_19;
  wire [29:0] pmp__EVAL_20;
  wire  pmp__EVAL_21;
  wire  pmp__EVAL_22;
  wire  pmp__EVAL_23;
  wire [31:0] pmp__EVAL_24;
  wire  pmp__EVAL_25;
  wire  pmp__EVAL_26;
  wire [31:0] pmp__EVAL_27;
  wire [31:0] pmp__EVAL_28;
  wire [31:0] pmp__EVAL_29;
  wire  pmp__EVAL_30;
  wire [1:0] pmp__EVAL_31;
  wire [1:0] pmp__EVAL_32;
  wire [29:0] pmp__EVAL_33;
  wire [31:0] pmp__EVAL_34;
  wire  pmp__EVAL_35;
  wire  pmp__EVAL_36;
  wire  pmp__EVAL_37;
  wire [31:0] pmp__EVAL_38;
  wire [31:0] pmp__EVAL_39;
  wire [1:0] pmp__EVAL_40;
  wire [29:0] pmp__EVAL_41;
  wire [29:0] pmp__EVAL_42;
  wire  pmp__EVAL_43;
  wire  pmp__EVAL_44;
  wire [29:0] pmp__EVAL_45;
  wire [31:0] pmp__EVAL_46;
  wire [1:0] pmp__EVAL_47;
  wire  pmp__EVAL_48;
  wire  pmp__EVAL_49;
  wire  pmp__EVAL_50;
  wire  pmp__EVAL_51;
  wire  pmp__EVAL_52;
  wire [29:0] pmp__EVAL_53;
  wire  pmp__EVAL_54;
  wire  pmp__EVAL_55;
  wire  pmp__EVAL_56;
  wire  pmp__EVAL_57;
  wire  pmp__EVAL_58;
  wire  pmp__EVAL_59;
  wire  pmp__EVAL_60;
  wire  pmp__EVAL_61;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire [31:0] _EVAL_79;
  wire [31:0] _EVAL_80;
  wire [13:0] _EVAL_81;
  wire [32:0] _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire [32:0] _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire [31:0] _EVAL_88;
  wire [31:0] _EVAL_89;
  wire [32:0] _EVAL_90;
  wire [32:0] _EVAL_91;
  wire [13:0] _EVAL_92;
  wire [13:0] _EVAL_93;
  wire [32:0] _EVAL_94;
  wire [1:0] _EVAL_95;
  wire [32:0] _EVAL_96;
  wire [32:0] _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire [32:0] _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire [31:0] _EVAL_105;
  wire [32:0] _EVAL_106;
  wire [32:0] _EVAL_107;
  wire  _EVAL_108;
  wire [31:0] _EVAL_109;
  wire [32:0] _EVAL_110;
  wire [32:0] _EVAL_111;
  wire [32:0] _EVAL_112;
  wire [32:0] _EVAL_113;
  wire [19:0] _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire [11:0] _EVAL_117;
  wire [32:0] _EVAL_118;
  wire [31:0] _EVAL_119;
  wire [32:0] _EVAL_120;
  wire [32:0] _EVAL_121;
  wire [32:0] _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire [32:0] _EVAL_127;
  wire [19:0] _EVAL_128;
  wire [32:0] _EVAL_129;
  wire [32:0] _EVAL_130;
  wire  _EVAL_131;
  wire [32:0] _EVAL_132;
  wire [32:0] _EVAL_133;
  wire  _EVAL_134;
  wire [32:0] _EVAL_135;
  wire  _EVAL_136;
  wire [32:0] _EVAL_137;
  wire [32:0] _EVAL_138;
  wire  _EVAL_139;
  wire [31:0] _EVAL_140;
  wire [32:0] _EVAL_141;
  wire  _EVAL_142;
  wire [32:0] _EVAL_143;
  _EVAL_105 pmp (
    ._EVAL(pmp__EVAL),
    ._EVAL_0(pmp__EVAL_0),
    ._EVAL_1(pmp__EVAL_1),
    ._EVAL_2(pmp__EVAL_2),
    ._EVAL_3(pmp__EVAL_3),
    ._EVAL_4(pmp__EVAL_4),
    ._EVAL_5(pmp__EVAL_5),
    ._EVAL_6(pmp__EVAL_6),
    ._EVAL_7(pmp__EVAL_7),
    ._EVAL_8(pmp__EVAL_8),
    ._EVAL_9(pmp__EVAL_9),
    ._EVAL_10(pmp__EVAL_10),
    ._EVAL_11(pmp__EVAL_11),
    ._EVAL_12(pmp__EVAL_12),
    ._EVAL_13(pmp__EVAL_13),
    ._EVAL_14(pmp__EVAL_14),
    ._EVAL_15(pmp__EVAL_15),
    ._EVAL_16(pmp__EVAL_16),
    ._EVAL_17(pmp__EVAL_17),
    ._EVAL_18(pmp__EVAL_18),
    ._EVAL_19(pmp__EVAL_19),
    ._EVAL_20(pmp__EVAL_20),
    ._EVAL_21(pmp__EVAL_21),
    ._EVAL_22(pmp__EVAL_22),
    ._EVAL_23(pmp__EVAL_23),
    ._EVAL_24(pmp__EVAL_24),
    ._EVAL_25(pmp__EVAL_25),
    ._EVAL_26(pmp__EVAL_26),
    ._EVAL_27(pmp__EVAL_27),
    ._EVAL_28(pmp__EVAL_28),
    ._EVAL_29(pmp__EVAL_29),
    ._EVAL_30(pmp__EVAL_30),
    ._EVAL_31(pmp__EVAL_31),
    ._EVAL_32(pmp__EVAL_32),
    ._EVAL_33(pmp__EVAL_33),
    ._EVAL_34(pmp__EVAL_34),
    ._EVAL_35(pmp__EVAL_35),
    ._EVAL_36(pmp__EVAL_36),
    ._EVAL_37(pmp__EVAL_37),
    ._EVAL_38(pmp__EVAL_38),
    ._EVAL_39(pmp__EVAL_39),
    ._EVAL_40(pmp__EVAL_40),
    ._EVAL_41(pmp__EVAL_41),
    ._EVAL_42(pmp__EVAL_42),
    ._EVAL_43(pmp__EVAL_43),
    ._EVAL_44(pmp__EVAL_44),
    ._EVAL_45(pmp__EVAL_45),
    ._EVAL_46(pmp__EVAL_46),
    ._EVAL_47(pmp__EVAL_47),
    ._EVAL_48(pmp__EVAL_48),
    ._EVAL_49(pmp__EVAL_49),
    ._EVAL_50(pmp__EVAL_50),
    ._EVAL_51(pmp__EVAL_51),
    ._EVAL_52(pmp__EVAL_52),
    ._EVAL_53(pmp__EVAL_53),
    ._EVAL_54(pmp__EVAL_54),
    ._EVAL_55(pmp__EVAL_55),
    ._EVAL_56(pmp__EVAL_56),
    ._EVAL_57(pmp__EVAL_57),
    ._EVAL_58(pmp__EVAL_58),
    ._EVAL_59(pmp__EVAL_59),
    ._EVAL_60(pmp__EVAL_60),
    ._EVAL_61(pmp__EVAL_61)
  );
  assign _EVAL_128 = _EVAL_39[31:12];
  assign _EVAL_129 = {1'b0,$signed(_EVAL_89)};
  assign pmp__EVAL_53 = _EVAL_61;
  assign _EVAL_132 = $signed(_EVAL_118) & -33'sh1000;
  assign pmp__EVAL_25 = _EVAL_52;
  assign _EVAL_82 = {1'b0,$signed(_EVAL_119)};
  assign _EVAL_136 = _EVAL_87 | _EVAL_73;
  assign pmp__EVAL_17 = _EVAL_27;
  assign _EVAL_124 = $signed(_EVAL_67) == 33'sh0;
  assign _EVAL_76 = _EVAL_135;
  assign pmp__EVAL_7 = _EVAL_53;
  assign _EVAL_116 = $signed(_EVAL_64) == 33'sh0;
  assign pmp__EVAL_39 = _EVAL_45;
  assign pmp__EVAL_26 = _EVAL_43;
  assign pmp__EVAL_42 = _EVAL_60;
  assign pmp__EVAL_10 = _EVAL_23;
  assign _EVAL_64 = _EVAL_102;
  assign _EVAL_137 = {1'b0,$signed(_EVAL_140)};
  assign _EVAL_118 = {1'b0,$signed(_EVAL_79)};
  assign pmp__EVAL_11 = _EVAL_32;
  assign _EVAL_94 = $signed(_EVAL_82) & -33'sh1000;
  assign _EVAL_88 = _EVAL_80 ^ 32'h80000000;
  assign _EVAL_135 = $signed(_EVAL_129) & -33'sh2000;
  assign pmp__EVAL_20 = _EVAL_37;
  assign _EVAL_84 = _EVAL_142 | _EVAL_116;
  assign _EVAL_122 = _EVAL_132;
  assign pmp__EVAL_19 = _EVAL_21;
  assign pmp__EVAL_43 = _EVAL_51;
  assign _EVAL_123 = $signed(_EVAL_122) == 33'sh0;
  assign _EVAL_107 = _EVAL_94;
  assign _EVAL_79 = _EVAL_80 ^ 32'h3000;
  assign _EVAL_98 = $signed(_EVAL_91) == 33'sh0;
  assign pmp__EVAL_40 = _EVAL_49;
  assign _EVAL_2 = {_EVAL_114,_EVAL_117};
  assign _EVAL_103 = _EVAL_84 | _EVAL_125;
  assign _EVAL_106 = {1'b0,$signed(_EVAL_80)};
  assign pmp__EVAL_29 = _EVAL_55;
  assign _EVAL_142 = _EVAL_62 | _EVAL_98;
  assign _EVAL_117 = _EVAL_39[11:0];
  assign pmp__EVAL_3 = _EVAL_44;
  assign _EVAL_141 = _EVAL_121;
  assign pmp__EVAL_21 = _EVAL_48;
  assign pmp__EVAL_12 = _EVAL_20;
  assign _EVAL_78 = ~_EVAL_69;
  assign _EVAL_131 = _EVAL_71 <= 3'h3;
  assign _EVAL_87 = _EVAL_134 | _EVAL_126;
  assign pmp__EVAL_27 = _EVAL_35;
  assign _EVAL_67 = _EVAL_138;
  assign pmp__EVAL_0 = _EVAL_14;
  assign _EVAL_73 = $signed(_EVAL_141) == 33'sh0;
  assign _EVAL_139 = _EVAL_136 | _EVAL_101;
  assign pmp__EVAL_28 = _EVAL_10;
  assign _EVAL_68 = _EVAL_112;
  assign pmp__EVAL_22 = _EVAL_28;
  assign pmp__EVAL_14 = _EVAL_29;
  assign _EVAL_114 = _EVAL_39[31:12];
  assign _EVAL_108 = $signed(_EVAL_76) == 33'sh0;
  assign _EVAL_85 = $signed(_EVAL_137) & 33'sheb004000;
  assign _EVAL_115 = _EVAL_103 | _EVAL_108;
  assign _EVAL_75 = _EVAL_123 | _EVAL_66;
  assign _EVAL_113 = {1'b0,$signed(_EVAL_105)};
  assign pmp__EVAL_57 = _EVAL_25;
  assign _EVAL_111 = _EVAL_143;
  assign _EVAL_91 = _EVAL_97;
  assign pmp__EVAL_60 = _EVAL_50;
  assign pmp__EVAL_13 = _EVAL_13;
  assign pmp__EVAL_33 = _EVAL_4;
  assign _EVAL_86 = $signed(_EVAL_63) == 33'sh0;
  assign _EVAL_100 = _EVAL_115 & _EVAL_139;
  assign _EVAL_138 = $signed(_EVAL_113) & -33'sh4000;
  assign pmp__EVAL_16 = _EVAL_38;
  assign _EVAL_63 = _EVAL_96;
  assign _EVAL_119 = _EVAL_80 ^ 32'h4000;
  assign pmp__EVAL_59 = _EVAL_18;
  assign pmp__EVAL_32 = _EVAL_57;
  assign pmp__EVAL_6 = _EVAL_33;
  assign _EVAL_80 = {_EVAL_128,_EVAL_117};
  assign _EVAL_90 = {1'b0,$signed(_EVAL_88)};
  assign pmp__EVAL_15 = _EVAL_1;
  assign _EVAL_97 = $signed(_EVAL_90) & -33'sh4000;
  assign pmp__EVAL_45 = _EVAL_30;
  assign pmp__EVAL_23 = _EVAL_46;
  assign _EVAL_104 = _EVAL_77 & pmp__EVAL;
  assign pmp__EVAL_38 = {_EVAL_128,_EVAL_117};
  assign _EVAL_77 = _EVAL_100 & _EVAL_78;
  assign _EVAL_126 = $signed(_EVAL_130) == 33'sh0;
  assign _EVAL_134 = $signed(_EVAL_65) == 33'sh0;
  assign pmp__EVAL_44 = _EVAL;
  assign pmp__EVAL_58 = _EVAL_9;
  assign pmp__EVAL_8 = _EVAL_26;
  assign _EVAL_127 = {1'b0,$signed(_EVAL_70)};
  assign pmp__EVAL_49 = _EVAL_54;
  assign _EVAL_125 = $signed(_EVAL_107) == 33'sh0;
  assign _EVAL_101 = $signed(_EVAL_72) == 33'sh0;
  assign _EVAL_121 = $signed(_EVAL_129) & 33'sheb004000;
  assign pmp__EVAL_18 = _EVAL_15;
  assign _EVAL_96 = $signed(_EVAL_127) & -33'sh10000;
  assign _EVAL_81 = _EVAL_92 & 14'h2000;
  assign _EVAL_62 = _EVAL_83 | _EVAL_124;
  assign pmp__EVAL_50 = _EVAL_59;
  assign _EVAL_130 = _EVAL_85;
  assign _EVAL_133 = $signed(_EVAL_106) & 33'shea004000;
  assign pmp__EVAL_47 = _EVAL_71[1:0];
  assign _EVAL_12 = |_EVAL_81;
  assign _EVAL_71 = {_EVAL_40,_EVAL_3};
  assign pmp__EVAL_48 = _EVAL_0;
  assign _EVAL_65 = _EVAL_133;
  assign _EVAL_93 = {_EVAL_95,12'h0};
  assign _EVAL_83 = _EVAL_74 | _EVAL_99;
  assign pmp__EVAL_51 = _EVAL_5;
  assign pmp__EVAL_61 = _EVAL_56;
  assign pmp__EVAL_1 = _EVAL_58;
  assign _EVAL_74 = _EVAL_75 | _EVAL_86;
  assign _EVAL_72 = _EVAL_110;
  assign pmp__EVAL_41 = _EVAL_31;
  assign _EVAL_112 = $signed(_EVAL_106) & -33'sh1000;
  assign _EVAL_120 = {1'b0,$signed(_EVAL_109)};
  assign pmp__EVAL_5 = _EVAL_22;
  assign pmp__EVAL_55 = _EVAL_34;
  assign pmp__EVAL_2 = _EVAL_41;
  assign pmp__EVAL_24 = _EVAL_47;
  assign pmp__EVAL_52 = _EVAL_16;
  assign pmp__EVAL_31 = _EVAL_36;
  assign pmp__EVAL_35 = _EVAL_19;
  assign _EVAL_92 = ~_EVAL_93;
  assign pmp__EVAL_37 = _EVAL_42;
  assign pmp__EVAL_36 = _EVAL_24;
  assign _EVAL_105 = _EVAL_80 ^ 32'h1800000;
  assign _EVAL_99 = $signed(_EVAL_68) == 33'sh0;
  assign _EVAL_109 = _EVAL_80 ^ 32'hc000000;
  assign pmp__EVAL_56 = _EVAL_7;
  assign pmp__EVAL_4 = _EVAL_11;
  assign _EVAL_70 = _EVAL_80 ^ 32'h2000000;
  assign _EVAL_102 = $signed(_EVAL_137) & -33'sh2000;
  assign _EVAL_95 = _EVAL_104 ? 2'h3 : 2'h0;
  assign _EVAL_89 = _EVAL_80 ^ 32'h40000000;
  assign pmp__EVAL_30 = _EVAL_17;
  assign pmp__EVAL_46 = _EVAL_8;
  assign _EVAL_66 = $signed(_EVAL_111) == 33'sh0;
  assign _EVAL_110 = $signed(_EVAL_90) & 33'sheb004000;
  assign _EVAL_69 = _EVAL_131 & _EVAL_99;
  assign _EVAL_143 = $signed(_EVAL_120) & -33'sh400000;
  assign pmp__EVAL_34 = _EVAL_6;
  assign _EVAL_140 = _EVAL_80 ^ 32'h20000000;
endmodule
