//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_17(
  input  [30:0] _EVAL,
  input         _EVAL_0,
  input  [2:0]  _EVAL_1,
  output        _EVAL_2,
  input         _EVAL_3,
  output        _EVAL_4,
  input         _EVAL_5,
  output [31:0] _EVAL_6,
  input         _EVAL_7,
  output [2:0]  _EVAL_8,
  output        _EVAL_9,
  input  [4:0]  _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  output [3:0]  _EVAL_13,
  output [30:0] _EVAL_14,
  output        _EVAL_15,
  output [2:0]  _EVAL_16,
  input  [31:0] _EVAL_17,
  input  [3:0]  _EVAL_18,
  input         _EVAL_19,
  input  [2:0]  _EVAL_20,
  output        _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23,
  output [2:0]  _EVAL_24,
  output [4:0]  _EVAL_25,
  output        _EVAL_26,
  output        _EVAL_27,
  input  [2:0]  _EVAL_28
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  _EVAL_29 [0:0];
  wire  _EVAL_29__EVAL_30_data;
  wire  _EVAL_29__EVAL_30_addr;
  wire  _EVAL_29__EVAL_31_data;
  wire  _EVAL_29__EVAL_31_addr;
  wire  _EVAL_29__EVAL_31_mask;
  wire  _EVAL_29__EVAL_31_en;
  wire  _EVAL_32;
  wire  _EVAL_33;
  reg [4:0] _EVAL_34 [0:0];
  wire [4:0] _EVAL_34__EVAL_35_data;
  wire  _EVAL_34__EVAL_35_addr;
  wire [4:0] _EVAL_34__EVAL_36_data;
  wire  _EVAL_34__EVAL_36_addr;
  wire  _EVAL_34__EVAL_36_mask;
  wire  _EVAL_34__EVAL_36_en;
  reg  _EVAL_37 [0:0];
  wire  _EVAL_37__EVAL_38_data;
  wire  _EVAL_37__EVAL_38_addr;
  wire  _EVAL_37__EVAL_39_data;
  wire  _EVAL_37__EVAL_39_addr;
  wire  _EVAL_37__EVAL_39_mask;
  wire  _EVAL_37__EVAL_39_en;
  wire  _EVAL_40;
  reg  _EVAL_41;
  reg [2:0] _EVAL_42 [0:0];
  wire [2:0] _EVAL_42__EVAL_43_data;
  wire  _EVAL_42__EVAL_43_addr;
  wire [2:0] _EVAL_42__EVAL_44_data;
  wire  _EVAL_42__EVAL_44_addr;
  wire  _EVAL_42__EVAL_44_mask;
  wire  _EVAL_42__EVAL_44_en;
  wire  _EVAL_45;
  wire  _EVAL_46;
  reg [31:0] _EVAL_47 [0:0];
  wire [31:0] _EVAL_47__EVAL_48_data;
  wire  _EVAL_47__EVAL_48_addr;
  wire [31:0] _EVAL_47__EVAL_49_data;
  wire  _EVAL_47__EVAL_49_addr;
  wire  _EVAL_47__EVAL_49_mask;
  wire  _EVAL_47__EVAL_49_en;
  reg [3:0] _EVAL_50 [0:0];
  wire [3:0] _EVAL_50__EVAL_51_data;
  wire  _EVAL_50__EVAL_51_addr;
  wire [3:0] _EVAL_50__EVAL_52_data;
  wire  _EVAL_50__EVAL_52_addr;
  wire  _EVAL_50__EVAL_52_mask;
  wire  _EVAL_50__EVAL_52_en;
  wire  _EVAL_53;
  reg  _EVAL_54 [0:0];
  wire  _EVAL_54__EVAL_55_data;
  wire  _EVAL_54__EVAL_55_addr;
  wire  _EVAL_54__EVAL_56_data;
  wire  _EVAL_54__EVAL_56_addr;
  wire  _EVAL_54__EVAL_56_mask;
  wire  _EVAL_54__EVAL_56_en;
  reg [2:0] _EVAL_57 [0:0];
  wire [2:0] _EVAL_57__EVAL_58_data;
  wire  _EVAL_57__EVAL_58_addr;
  wire [2:0] _EVAL_57__EVAL_59_data;
  wire  _EVAL_57__EVAL_59_addr;
  wire  _EVAL_57__EVAL_59_mask;
  wire  _EVAL_57__EVAL_59_en;
  reg  _EVAL_60 [0:0];
  wire  _EVAL_60__EVAL_61_data;
  wire  _EVAL_60__EVAL_61_addr;
  wire  _EVAL_60__EVAL_62_data;
  wire  _EVAL_60__EVAL_62_addr;
  wire  _EVAL_60__EVAL_62_mask;
  wire  _EVAL_60__EVAL_62_en;
  reg [2:0] _EVAL_63 [0:0];
  wire [2:0] _EVAL_63__EVAL_64_data;
  wire  _EVAL_63__EVAL_64_addr;
  wire [2:0] _EVAL_63__EVAL_65_data;
  wire  _EVAL_63__EVAL_65_addr;
  wire  _EVAL_63__EVAL_65_mask;
  wire  _EVAL_63__EVAL_65_en;
  reg [30:0] _EVAL_66 [0:0];
  wire [30:0] _EVAL_66__EVAL_67_data;
  wire  _EVAL_66__EVAL_67_addr;
  wire [30:0] _EVAL_66__EVAL_68_data;
  wire  _EVAL_66__EVAL_68_addr;
  wire  _EVAL_66__EVAL_68_mask;
  wire  _EVAL_66__EVAL_68_en;
  wire  _EVAL_69;
  reg  _EVAL_71 [0:0];
  wire  _EVAL_71__EVAL_72_data;
  wire  _EVAL_71__EVAL_72_addr;
  wire  _EVAL_71__EVAL_73_data;
  wire  _EVAL_71__EVAL_73_addr;
  wire  _EVAL_71__EVAL_73_mask;
  wire  _EVAL_71__EVAL_73_en;
  wire  _EVAL_74;
  assign _EVAL_29__EVAL_30_addr = 1'h0;
  assign _EVAL_29__EVAL_30_data = _EVAL_29[_EVAL_29__EVAL_30_addr];
  assign _EVAL_29__EVAL_31_data = _EVAL_5;
  assign _EVAL_29__EVAL_31_addr = 1'h0;
  assign _EVAL_29__EVAL_31_mask = 1'h1;
  assign _EVAL_29__EVAL_31_en = _EVAL_69 ? _EVAL_40 : _EVAL_32;
  assign _EVAL_34__EVAL_35_addr = 1'h0;
  assign _EVAL_34__EVAL_35_data = _EVAL_34[_EVAL_34__EVAL_35_addr];
  assign _EVAL_34__EVAL_36_data = _EVAL_10;
  assign _EVAL_34__EVAL_36_addr = 1'h0;
  assign _EVAL_34__EVAL_36_mask = 1'h1;
  assign _EVAL_34__EVAL_36_en = _EVAL_69 ? _EVAL_40 : _EVAL_32;
  assign _EVAL_37__EVAL_38_addr = 1'h0;
  assign _EVAL_37__EVAL_38_data = _EVAL_37[_EVAL_37__EVAL_38_addr];
  assign _EVAL_37__EVAL_39_data = _EVAL_0;
  assign _EVAL_37__EVAL_39_addr = 1'h0;
  assign _EVAL_37__EVAL_39_mask = 1'h1;
  assign _EVAL_37__EVAL_39_en = _EVAL_69 ? _EVAL_40 : _EVAL_32;
  assign _EVAL_42__EVAL_43_addr = 1'h0;
  assign _EVAL_42__EVAL_43_data = _EVAL_42[_EVAL_42__EVAL_43_addr];
  assign _EVAL_42__EVAL_44_data = _EVAL_20;
  assign _EVAL_42__EVAL_44_addr = 1'h0;
  assign _EVAL_42__EVAL_44_mask = 1'h1;
  assign _EVAL_42__EVAL_44_en = _EVAL_69 ? _EVAL_40 : _EVAL_32;
  assign _EVAL_47__EVAL_48_addr = 1'h0;
  assign _EVAL_47__EVAL_48_data = _EVAL_47[_EVAL_47__EVAL_48_addr];
  assign _EVAL_47__EVAL_49_data = _EVAL_17;
  assign _EVAL_47__EVAL_49_addr = 1'h0;
  assign _EVAL_47__EVAL_49_mask = 1'h1;
  assign _EVAL_47__EVAL_49_en = _EVAL_69 ? _EVAL_40 : _EVAL_32;
  assign _EVAL_50__EVAL_51_addr = 1'h0;
  assign _EVAL_50__EVAL_51_data = _EVAL_50[_EVAL_50__EVAL_51_addr];
  assign _EVAL_50__EVAL_52_data = _EVAL_18;
  assign _EVAL_50__EVAL_52_addr = 1'h0;
  assign _EVAL_50__EVAL_52_mask = 1'h1;
  assign _EVAL_50__EVAL_52_en = _EVAL_69 ? _EVAL_40 : _EVAL_32;
  assign _EVAL_54__EVAL_55_addr = 1'h0;
  assign _EVAL_54__EVAL_55_data = _EVAL_54[_EVAL_54__EVAL_55_addr];
  assign _EVAL_54__EVAL_56_data = _EVAL_19;
  assign _EVAL_54__EVAL_56_addr = 1'h0;
  assign _EVAL_54__EVAL_56_mask = 1'h1;
  assign _EVAL_54__EVAL_56_en = _EVAL_69 ? _EVAL_40 : _EVAL_32;
  assign _EVAL_57__EVAL_58_addr = 1'h0;
  assign _EVAL_57__EVAL_58_data = _EVAL_57[_EVAL_57__EVAL_58_addr];
  assign _EVAL_57__EVAL_59_data = _EVAL_1;
  assign _EVAL_57__EVAL_59_addr = 1'h0;
  assign _EVAL_57__EVAL_59_mask = 1'h1;
  assign _EVAL_57__EVAL_59_en = _EVAL_69 ? _EVAL_40 : _EVAL_32;
  assign _EVAL_60__EVAL_61_addr = 1'h0;
  assign _EVAL_60__EVAL_61_data = _EVAL_60[_EVAL_60__EVAL_61_addr];
  assign _EVAL_60__EVAL_62_data = _EVAL_7;
  assign _EVAL_60__EVAL_62_addr = 1'h0;
  assign _EVAL_60__EVAL_62_mask = 1'h1;
  assign _EVAL_60__EVAL_62_en = _EVAL_69 ? _EVAL_40 : _EVAL_32;
  assign _EVAL_63__EVAL_64_addr = 1'h0;
  assign _EVAL_63__EVAL_64_data = _EVAL_63[_EVAL_63__EVAL_64_addr];
  assign _EVAL_63__EVAL_65_data = _EVAL_28;
  assign _EVAL_63__EVAL_65_addr = 1'h0;
  assign _EVAL_63__EVAL_65_mask = 1'h1;
  assign _EVAL_63__EVAL_65_en = _EVAL_69 ? _EVAL_40 : _EVAL_32;
  assign _EVAL_66__EVAL_67_addr = 1'h0;
  assign _EVAL_66__EVAL_67_data = _EVAL_66[_EVAL_66__EVAL_67_addr];
  assign _EVAL_66__EVAL_68_data = _EVAL;
  assign _EVAL_66__EVAL_68_addr = 1'h0;
  assign _EVAL_66__EVAL_68_mask = 1'h1;
  assign _EVAL_66__EVAL_68_en = _EVAL_69 ? _EVAL_40 : _EVAL_32;
  assign _EVAL_71__EVAL_72_addr = 1'h0;
  assign _EVAL_71__EVAL_72_data = _EVAL_71[_EVAL_71__EVAL_72_addr];
  assign _EVAL_71__EVAL_73_data = _EVAL_22;
  assign _EVAL_71__EVAL_73_addr = 1'h0;
  assign _EVAL_71__EVAL_73_mask = 1'h1;
  assign _EVAL_71__EVAL_73_en = _EVAL_69 ? _EVAL_40 : _EVAL_32;
  assign _EVAL_2 = ~_EVAL_41;
  assign _EVAL_33 = _EVAL_74 != _EVAL_53;
  assign _EVAL_16 = _EVAL_69 ? _EVAL_1 : _EVAL_57__EVAL_58_data;
  assign _EVAL_46 = ~_EVAL_69;
  assign _EVAL_53 = _EVAL_69 ? 1'h0 : _EVAL_45;
  assign _EVAL_24 = _EVAL_69 ? _EVAL_20 : _EVAL_42__EVAL_43_data;
  assign _EVAL_74 = _EVAL_69 ? _EVAL_40 : _EVAL_32;
  assign _EVAL_6 = _EVAL_69 ? _EVAL_17 : _EVAL_47__EVAL_48_data;
  assign _EVAL_45 = _EVAL_12 & _EVAL_21;
  assign _EVAL_26 = _EVAL_69 ? _EVAL_22 : _EVAL_71__EVAL_72_data;
  assign _EVAL_8 = _EVAL_69 ? _EVAL_28 : _EVAL_63__EVAL_64_data;
  assign _EVAL_32 = _EVAL_2 & _EVAL_3;
  assign _EVAL_27 = _EVAL_69 ? _EVAL_5 : _EVAL_29__EVAL_30_data;
  assign _EVAL_4 = _EVAL_69 ? _EVAL_7 : _EVAL_60__EVAL_61_data;
  assign _EVAL_69 = ~_EVAL_41;
  assign _EVAL_9 = _EVAL_69 ? _EVAL_0 : _EVAL_37__EVAL_38_data;
  assign _EVAL_21 = _EVAL_3 | _EVAL_46;
  assign _EVAL_15 = _EVAL_69 ? _EVAL_19 : _EVAL_54__EVAL_55_data;
  assign _EVAL_25 = _EVAL_69 ? _EVAL_10 : _EVAL_34__EVAL_35_data;
  assign _EVAL_14 = _EVAL_69 ? _EVAL : _EVAL_66__EVAL_67_data;
  assign _EVAL_13 = _EVAL_69 ? _EVAL_18 : _EVAL_50__EVAL_51_data;
  assign _EVAL_40 = _EVAL_12 ? 1'h0 : _EVAL_32;
  always @(posedge _EVAL_11) begin
    if(_EVAL_29__EVAL_31_en & _EVAL_29__EVAL_31_mask) begin
      _EVAL_29[_EVAL_29__EVAL_31_addr] <= _EVAL_29__EVAL_31_data;
    end
    if(_EVAL_34__EVAL_36_en & _EVAL_34__EVAL_36_mask) begin
      _EVAL_34[_EVAL_34__EVAL_36_addr] <= _EVAL_34__EVAL_36_data;
    end
    if(_EVAL_37__EVAL_39_en & _EVAL_37__EVAL_39_mask) begin
      _EVAL_37[_EVAL_37__EVAL_39_addr] <= _EVAL_37__EVAL_39_data;
    end
    if (_EVAL_23) begin
      _EVAL_41 <= 1'h0;
    end else if (_EVAL_33) begin
      if (_EVAL_69) begin
        if (_EVAL_12) begin
          _EVAL_41 <= 1'h0;
        end else begin
          _EVAL_41 <= _EVAL_32;
        end
      end else begin
        _EVAL_41 <= _EVAL_32;
      end
    end
    if(_EVAL_42__EVAL_44_en & _EVAL_42__EVAL_44_mask) begin
      _EVAL_42[_EVAL_42__EVAL_44_addr] <= _EVAL_42__EVAL_44_data;
    end
    if(_EVAL_47__EVAL_49_en & _EVAL_47__EVAL_49_mask) begin
      _EVAL_47[_EVAL_47__EVAL_49_addr] <= _EVAL_47__EVAL_49_data;
    end
    if(_EVAL_50__EVAL_52_en & _EVAL_50__EVAL_52_mask) begin
      _EVAL_50[_EVAL_50__EVAL_52_addr] <= _EVAL_50__EVAL_52_data;
    end
    if(_EVAL_54__EVAL_56_en & _EVAL_54__EVAL_56_mask) begin
      _EVAL_54[_EVAL_54__EVAL_56_addr] <= _EVAL_54__EVAL_56_data;
    end
    if(_EVAL_57__EVAL_59_en & _EVAL_57__EVAL_59_mask) begin
      _EVAL_57[_EVAL_57__EVAL_59_addr] <= _EVAL_57__EVAL_59_data;
    end
    if(_EVAL_60__EVAL_62_en & _EVAL_60__EVAL_62_mask) begin
      _EVAL_60[_EVAL_60__EVAL_62_addr] <= _EVAL_60__EVAL_62_data;
    end
    if(_EVAL_63__EVAL_65_en & _EVAL_63__EVAL_65_mask) begin
      _EVAL_63[_EVAL_63__EVAL_65_addr] <= _EVAL_63__EVAL_65_data;
    end
    if(_EVAL_66__EVAL_68_en & _EVAL_66__EVAL_68_mask) begin
      _EVAL_66[_EVAL_66__EVAL_68_addr] <= _EVAL_66__EVAL_68_data;
    end
    if(_EVAL_71__EVAL_73_en & _EVAL_71__EVAL_73_mask) begin
      _EVAL_71[_EVAL_71__EVAL_73_addr] <= _EVAL_71__EVAL_73_data;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_29[initvar] = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_34[initvar] = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_37[initvar] = _RAND_2[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_42[initvar] = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_47[initvar] = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_50[initvar] = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_54[initvar] = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_57[initvar] = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_60[initvar] = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_63[initvar] = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_66[initvar] = _RAND_11[30:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    _EVAL_71[initvar] = _RAND_12[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _EVAL_41 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
