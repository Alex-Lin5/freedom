//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_133(
  output        _EVAL,
  input         _EVAL_0,
  input  [31:0] _EVAL_1,
  input  [6:0]  _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  output        _EVAL_5,
  output        _EVAL_6,
  output        _EVAL_7,
  input         _EVAL_8,
  output [4:0]  _EVAL_9,
  output        _EVAL_10,
  output [1:0]  _EVAL_11,
  input         _EVAL_12,
  output        _EVAL_13,
  output        _EVAL_14,
  output [31:0] _EVAL_15,
  output [3:0]  _EVAL_16,
  output        _EVAL_17,
  input         _EVAL_18,
  output        _EVAL_19,
  output [31:0] _EVAL_20,
  output        _EVAL_21,
  input  [1:0]  _EVAL_22,
  input         _EVAL_23,
  output        _EVAL_24,
  output [29:0] _EVAL_25,
  output [1:0]  _EVAL_26,
  output [31:0] _EVAL_27,
  output        _EVAL_28,
  output [31:0] _EVAL_29,
  output [29:0] _EVAL_30,
  input         _EVAL_31,
  input         _EVAL_32,
  output [1:0]  _EVAL_33,
  output [1:0]  _EVAL_34,
  output [1:0]  _EVAL_35,
  output [31:0] _EVAL_36,
  output        _EVAL_37,
  output [29:0] _EVAL_38,
  input         _EVAL_39,
  output        _EVAL_40,
  output        _EVAL_41,
  input         _EVAL_42,
  input  [4:0]  _EVAL_43,
  input  [31:0] _EVAL_44,
  input  [4:0]  _EVAL_45,
  input  [1:0]  _EVAL_46,
  input         _EVAL_47,
  input  [31:0] _EVAL_48,
  output [1:0]  _EVAL_49,
  output        _EVAL_50,
  output [31:0] _EVAL_51,
  output        _EVAL_52,
  input         _EVAL_53,
  output [1:0]  _EVAL_54,
  output        _EVAL_55,
  output        _EVAL_56,
  input         _EVAL_57,
  output        _EVAL_58,
  input         _EVAL_59,
  output [4:0]  _EVAL_60,
  output        _EVAL_61,
  output [31:0] _EVAL_62,
  input         _EVAL_63,
  output [1:0]  _EVAL_64,
  output        _EVAL_65,
  output [31:0] _EVAL_66,
  output        _EVAL_67,
  output [1:0]  _EVAL_68,
  input  [31:0] _EVAL_69,
  output [1:0]  _EVAL_70,
  input  [7:0]  _EVAL_71,
  input  [31:0] _EVAL_72,
  output        _EVAL_73,
  input         _EVAL_74,
  output [31:0] _EVAL_75,
  output [6:0]  _EVAL_76,
  output        _EVAL_77,
  output        _EVAL_78,
  output        _EVAL_79,
  input         _EVAL_80,
  input         _EVAL_81,
  input         _EVAL_82,
  input         _EVAL_83,
  input         _EVAL_84,
  input         _EVAL_85,
  output        _EVAL_86,
  output        _EVAL_87,
  output        _EVAL_88,
  output [1:0]  _EVAL_89,
  input         _EVAL_90,
  output [31:0] _EVAL_91,
  input         _EVAL_92,
  output        _EVAL_93,
  output        _EVAL_94,
  output [31:0] _EVAL_95,
  output        _EVAL_96,
  output        _EVAL_97,
  output        _EVAL_98,
  output        _EVAL_99,
  input         _EVAL_100,
  output        _EVAL_101,
  output        _EVAL_102,
  input         _EVAL_103,
  output [31:0] _EVAL_104,
  input         _EVAL_105,
  input         _EVAL_106,
  input         _EVAL_107,
  output [31:0] _EVAL_108,
  input         _EVAL_109,
  output [1:0]  _EVAL_110,
  input         _EVAL_111,
  output [31:0] _EVAL_112,
  input  [31:0] _EVAL_113,
  output        _EVAL_114,
  input         _EVAL_115,
  input         _EVAL_116,
  input         _EVAL_117,
  input         _EVAL_118,
  input         _EVAL_119,
  output        _EVAL_120,
  output        _EVAL_121,
  input         _EVAL_122,
  output        _EVAL_123,
  output        _EVAL_124,
  output [31:0] _EVAL_125,
  input         _EVAL_126,
  output        _EVAL_127,
  output [7:0]  _EVAL_128,
  output        _EVAL_129,
  output        _EVAL_130,
  input         _EVAL_131,
  output        _EVAL_132,
  output [29:0] _EVAL_133,
  output        _EVAL_134,
  input         _EVAL_135,
  output [29:0] _EVAL_136,
  output        _EVAL_137,
  output [29:0] _EVAL_138,
  output        _EVAL_139,
  input         _EVAL_140,
  input         _EVAL_141,
  output [1:0]  _EVAL_142,
  output        _EVAL_143,
  output        _EVAL_144,
  output        _EVAL_145,
  output [31:0] _EVAL_146,
  input         _EVAL_147,
  output [31:0] _EVAL_148,
  input         _EVAL_149,
  input         _EVAL_150,
  input         _EVAL_151,
  input  [31:0] _EVAL_152,
  output [3:0]  _EVAL_153,
  input         _EVAL_154,
  output [29:0] _EVAL_155,
  output [29:0] _EVAL_156,
  input         _EVAL_157,
  input         _EVAL_158,
  output        _EVAL_159,
  input         _EVAL_160,
  output        _EVAL_161
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_162;
  wire [31:0] _EVAL_163;
  wire [31:0] _EVAL_164;
  wire  _EVAL_165;
  wire [31:0] _EVAL_166;
  wire [31:0] _EVAL_167;
  wire [4:0] _EVAL_168;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire [31:0] _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire [31:0] _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_180;
  wire [4:0] _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_184;
  wire [1:0] _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire [31:0] _EVAL_191;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire [31:0] _EVAL_195;
  wire  _EVAL_196;
  wire [31:0] bpu__EVAL;
  wire  bpu__EVAL_0;
  wire  bpu__EVAL_1;
  wire  bpu__EVAL_2;
  wire  bpu__EVAL_3;
  wire  bpu__EVAL_4;
  wire  bpu__EVAL_5;
  wire  bpu__EVAL_6;
  wire [1:0] bpu__EVAL_7;
  wire [31:0] bpu__EVAL_8;
  wire  bpu__EVAL_9;
  wire  bpu__EVAL_10;
  wire  bpu__EVAL_11;
  wire  bpu__EVAL_12;
  wire  bpu__EVAL_13;
  wire  bpu__EVAL_14;
  wire  bpu__EVAL_15;
  wire  bpu__EVAL_16;
  wire  bpu__EVAL_17;
  wire [1:0] bpu__EVAL_18;
  wire [1:0] bpu__EVAL_19;
  wire  bpu__EVAL_20;
  wire [31:0] bpu__EVAL_21;
  wire  bpu__EVAL_22;
  wire [31:0] bpu__EVAL_23;
  wire  bpu__EVAL_24;
  wire  bpu__EVAL_25;
  wire  bpu__EVAL_26;
  wire  bpu__EVAL_27;
  wire  bpu__EVAL_28;
  wire [31:0] bpu__EVAL_29;
  wire  bpu__EVAL_30;
  wire [31:0] bpu__EVAL_31;
  wire  bpu__EVAL_32;
  wire  bpu__EVAL_33;
  wire [1:0] bpu__EVAL_34;
  wire  bpu__EVAL_35;
  wire  bpu__EVAL_36;
  wire  bpu__EVAL_37;
  wire  bpu__EVAL_38;
  wire  bpu__EVAL_39;
  wire  bpu__EVAL_40;
  wire  bpu__EVAL_41;
  wire [1:0] bpu__EVAL_42;
  wire  bpu__EVAL_43;
  wire  _EVAL_197;
  wire [31:0] _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire [31:0] _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire [31:0] _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire [3:0] _EVAL_223;
  wire [31:0] _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire [31:0] _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire [23:0] _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire [32:0] _EVAL_240;
  wire [5:0] _EVAL_241;
  wire  _EVAL_242;
  wire [3:0] _EVAL_243;
  wire [31:0] _EVAL_244;
  wire [31:0] _EVAL_245;
  wire  csr__EVAL;
  wire [1:0] csr__EVAL_0;
  wire [31:0] csr__EVAL_1;
  wire  csr__EVAL_2;
  wire  csr__EVAL_3;
  wire [31:0] csr__EVAL_4;
  wire  csr__EVAL_5;
  wire  csr__EVAL_6;
  wire  csr__EVAL_7;
  wire  csr__EVAL_8;
  wire  csr__EVAL_9;
  wire  csr__EVAL_10;
  wire  csr__EVAL_11;
  wire  csr__EVAL_12;
  wire [1:0] csr__EVAL_13;
  wire [1:0] csr__EVAL_14;
  wire [31:0] csr__EVAL_15;
  wire  csr__EVAL_16;
  wire  csr__EVAL_17;
  wire  csr__EVAL_18;
  wire  csr__EVAL_19;
  wire  csr__EVAL_20;
  wire  csr__EVAL_21;
  wire  csr__EVAL_22;
  wire  csr__EVAL_23;
  wire [1:0] csr__EVAL_24;
  wire  csr__EVAL_25;
  wire [1:0] csr__EVAL_26;
  wire [31:0] csr__EVAL_27;
  wire [31:0] csr__EVAL_28;
  wire  csr__EVAL_29;
  wire  csr__EVAL_30;
  wire [1:0] csr__EVAL_31;
  wire  csr__EVAL_32;
  wire  csr__EVAL_33;
  wire [31:0] csr__EVAL_34;
  wire  csr__EVAL_35;
  wire  csr__EVAL_36;
  wire  csr__EVAL_37;
  wire  csr__EVAL_38;
  wire  csr__EVAL_39;
  wire [29:0] csr__EVAL_40;
  wire  csr__EVAL_41;
  wire [29:0] csr__EVAL_42;
  wire [1:0] csr__EVAL_43;
  wire [31:0] csr__EVAL_44;
  wire  csr__EVAL_45;
  wire [31:0] csr__EVAL_46;
  wire  csr__EVAL_47;
  wire  csr__EVAL_48;
  wire  csr__EVAL_49;
  wire [31:0] csr__EVAL_50;
  wire  csr__EVAL_51;
  wire [31:0] csr__EVAL_52;
  wire  csr__EVAL_53;
  wire  csr__EVAL_54;
  wire  csr__EVAL_55;
  wire [31:0] csr__EVAL_56;
  wire  csr__EVAL_57;
  wire  csr__EVAL_58;
  wire  csr__EVAL_59;
  wire [1:0] csr__EVAL_60;
  wire  csr__EVAL_61;
  wire  csr__EVAL_62;
  wire  csr__EVAL_63;
  wire [31:0] csr__EVAL_64;
  wire  csr__EVAL_65;
  wire  csr__EVAL_66;
  wire [1:0] csr__EVAL_67;
  wire  csr__EVAL_68;
  wire  csr__EVAL_69;
  wire [31:0] csr__EVAL_70;
  wire [31:0] csr__EVAL_71;
  wire  csr__EVAL_72;
  wire [31:0] csr__EVAL_73;
  wire  csr__EVAL_74;
  wire  csr__EVAL_75;
  wire  csr__EVAL_76;
  wire  csr__EVAL_77;
  wire  csr__EVAL_78;
  wire  csr__EVAL_79;
  wire  csr__EVAL_80;
  wire  csr__EVAL_81;
  wire [7:0] csr__EVAL_82;
  wire  csr__EVAL_83;
  wire  csr__EVAL_84;
  wire  csr__EVAL_85;
  wire  csr__EVAL_86;
  wire [29:0] csr__EVAL_87;
  wire  csr__EVAL_88;
  wire [1:0] csr__EVAL_89;
  wire  csr__EVAL_90;
  wire  csr__EVAL_91;
  wire [1:0] csr__EVAL_92;
  wire  csr__EVAL_93;
  wire [31:0] csr__EVAL_94;
  wire  csr__EVAL_95;
  wire  csr__EVAL_96;
  wire [31:0] csr__EVAL_97;
  wire  csr__EVAL_98;
  wire  csr__EVAL_99;
  wire [1:0] csr__EVAL_100;
  wire [31:0] csr__EVAL_101;
  wire  csr__EVAL_102;
  wire [31:0] csr__EVAL_103;
  wire [31:0] csr__EVAL_104;
  wire [29:0] csr__EVAL_105;
  wire  csr__EVAL_106;
  wire  csr__EVAL_107;
  wire [2:0] csr__EVAL_108;
  wire  csr__EVAL_109;
  wire  csr__EVAL_110;
  wire  csr__EVAL_111;
  wire  csr__EVAL_112;
  wire [11:0] csr__EVAL_113;
  wire  csr__EVAL_114;
  wire  csr__EVAL_115;
  wire [31:0] csr__EVAL_116;
  wire  csr__EVAL_117;
  wire [31:0] csr__EVAL_118;
  wire  csr__EVAL_119;
  wire  csr__EVAL_120;
  wire  csr__EVAL_121;
  wire [26:0] csr__EVAL_122;
  wire [1:0] csr__EVAL_123;
  wire [31:0] csr__EVAL_124;
  wire [1:0] csr__EVAL_125;
  wire  csr__EVAL_126;
  wire  csr__EVAL_127;
  wire  csr__EVAL_128;
  wire  csr__EVAL_129;
  wire [31:0] csr__EVAL_130;
  wire  csr__EVAL_131;
  wire  csr__EVAL_132;
  wire [31:0] csr__EVAL_133;
  wire [2:0] csr__EVAL_134;
  wire  csr__EVAL_135;
  wire  csr__EVAL_136;
  wire  csr__EVAL_137;
  wire  csr__EVAL_138;
  wire [1:0] csr__EVAL_139;
  wire [31:0] csr__EVAL_140;
  wire  csr__EVAL_141;
  wire  csr__EVAL_142;
  wire [1:0] csr__EVAL_143;
  wire [29:0] csr__EVAL_144;
  wire [31:0] csr__EVAL_145;
  wire  csr__EVAL_146;
  wire  csr__EVAL_147;
  wire [29:0] csr__EVAL_148;
  wire  csr__EVAL_149;
  wire  csr__EVAL_150;
  wire [11:0] csr__EVAL_151;
  wire  csr__EVAL_152;
  wire  csr__EVAL_153;
  wire  csr__EVAL_154;
  wire  csr__EVAL_155;
  wire  csr__EVAL_156;
  wire  csr__EVAL_157;
  wire [31:0] csr__EVAL_158;
  wire  csr__EVAL_159;
  wire [29:0] csr__EVAL_160;
  wire [31:0] csr__EVAL_161;
  wire [1:0] csr__EVAL_162;
  wire [29:0] csr__EVAL_163;
  wire  csr__EVAL_164;
  wire [31:0] csr__EVAL_165;
  wire  csr__EVAL_166;
  wire  csr__EVAL_167;
  wire  csr__EVAL_168;
  wire [31:0] csr__EVAL_169;
  wire  csr__EVAL_170;
  wire [1:0] csr__EVAL_171;
  wire  csr__EVAL_172;
  wire  csr__EVAL_173;
  wire  csr__EVAL_174;
  wire  csr__EVAL_175;
  wire [1:0] csr__EVAL_176;
  wire [1:0] csr__EVAL_177;
  wire  csr__EVAL_178;
  wire  csr__EVAL_179;
  wire  csr__EVAL_180;
  wire  csr__EVAL_181;
  wire  csr__EVAL_182;
  wire  csr__EVAL_183;
  wire  csr__EVAL_184;
  wire  csr__EVAL_185;
  wire  csr__EVAL_186;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire [3:0] _EVAL_262;
  wire  _EVAL_263;
  wire [7:0] _EVAL_264;
  wire  _EVAL_265;
  wire [31:0] _EVAL_266;
  wire  _EVAL_268;
  wire [31:0] _EVAL_269;
  wire  _EVAL_270;
  wire [1:0] _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire [31:0] _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire [3:0] _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire [31:0] _EVAL_285;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire  _EVAL_294;
  wire  _EVAL_295;
  wire  _EVAL_296;
  wire  _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_308;
  wire  _EVAL_309;
  wire [31:0] _EVAL_310;
  wire  _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_317;
  wire  _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_320;
  wire [31:0] _EVAL_322;
  wire  _EVAL_323;
  wire [2:0] _EVAL_324;
  wire  _EVAL_325;
  wire  _EVAL_326;
  wire  _EVAL_327;
  wire  _EVAL_328;
  wire  _EVAL_329;
  wire  _EVAL_330;
  wire [15:0] _EVAL_331;
  wire  _EVAL_332;
  wire  _EVAL_333;
  wire [31:0] _EVAL_334;
  wire  _EVAL_335;
  wire  _EVAL_336;
  reg  _EVAL_337;
  wire  _EVAL_338;
  wire [15:0] _EVAL_339;
  wire  _EVAL_340;
  wire  _EVAL_341;
  wire  _EVAL_342;
  wire  _EVAL_343;
  wire  _EVAL_344;
  wire [4:0] _EVAL_345;
  wire  _EVAL_346;
  wire  _EVAL_347;
  wire [4:0] _EVAL_348;
  wire [31:0] _EVAL_349;
  wire [31:0] _EVAL_350;
  wire  _EVAL_352;
  wire  _EVAL_353;
  wire  _EVAL_354;
  wire [31:0] _EVAL_355;
  wire  _EVAL_356;
  wire  _EVAL_357;
  wire  _EVAL_359;
  wire [31:0] _EVAL_361;
  wire  _EVAL_362;
  wire  _EVAL_363;
  wire [31:0] _EVAL_364;
  wire  _EVAL_365;
  wire  _EVAL_366;
  wire  _EVAL_367;
  wire  _EVAL_368;
  wire  _EVAL_369;
  wire  _EVAL_370;
  wire  _EVAL_371;
  wire [3:0] _EVAL_372;
  wire [31:0] _EVAL_373;
  wire  _EVAL_374;
  wire  _EVAL_375;
  wire  _EVAL_376;
  wire  _EVAL_377;
  wire  _EVAL_378;
  wire  _EVAL_379;
  wire  _EVAL_380;
  wire  _EVAL_381;
  wire  _EVAL_382;
  wire  _EVAL_384;
  wire  _EVAL_385;
  wire [1:0] _EVAL_386;
  wire  _EVAL_387;
  wire  _EVAL_389;
  wire  _EVAL_390;
  wire  _EVAL_391;
  wire  _EVAL_392;
  wire  _EVAL_393;
  wire  _EVAL_394;
  wire  _EVAL_395;
  wire  _EVAL_396;
  wire  _EVAL_397;
  wire  _EVAL_398;
  wire  _EVAL_400;
  wire  _EVAL_401;
  wire  _EVAL_402;
  wire  _EVAL_403;
  wire  _EVAL_404;
  wire  _EVAL_405;
  wire [23:0] _EVAL_406;
  wire [31:0] _EVAL_407;
  wire  _EVAL_408;
  wire  _EVAL_409;
  wire  _EVAL_410;
  wire  _EVAL_411;
  wire  _EVAL_412;
  wire  _EVAL_413;
  wire [1:0] _EVAL_414;
  wire  _EVAL_415;
  wire  _EVAL_417;
  wire  _EVAL_418;
  wire  _EVAL_419;
  wire  _EVAL_420;
  wire  _EVAL_421;
  wire  _EVAL_422;
  wire  _EVAL_423;
  wire  _EVAL_424;
  wire  _EVAL_425;
  wire [2:0] _EVAL_426;
  wire [10:0] _EVAL_427;
  wire  _EVAL_428;
  wire [10:0] _EVAL_429;
  wire  _EVAL_430;
  wire  _EVAL_431;
  wire  _EVAL_432;
  wire  _EVAL_433;
  wire  _EVAL_434;
  wire [31:0] _EVAL_435;
  wire  _EVAL_436;
  wire  _EVAL_437;
  wire  _EVAL_438;
  wire  _EVAL_439;
  wire  _EVAL_440;
  wire [31:0] _EVAL_441;
  wire  _EVAL_442;
  wire  _EVAL_443;
  wire [1:0] _EVAL_444;
  wire  _EVAL_445;
  wire [31:0] _EVAL_447;
  wire  _EVAL_448;
  wire  _EVAL_449;
  wire [1:0] _EVAL_450;
  wire [31:0] _EVAL_451;
  wire  _EVAL_452;
  wire  _EVAL_453;
  wire  _EVAL_454;
  wire  _EVAL_455;
  wire  _EVAL_457;
  wire  _EVAL_458;
  wire  _EVAL_459;
  wire  _EVAL_460;
  wire  _EVAL_461;
  wire  _EVAL_462;
  wire  _EVAL_463;
  wire  _EVAL_464;
  wire  _EVAL_465;
  wire [31:0] _EVAL_466;
  wire  _EVAL_467;
  wire [23:0] _EVAL_469;
  wire  _EVAL_470;
  wire  _EVAL_471;
  wire  _EVAL_472;
  reg  _EVAL_473;
  wire  _EVAL_475;
  wire [31:0] _EVAL_477;
  wire [31:0] _EVAL_478;
  wire  _EVAL_479;
  wire  _EVAL_480;
  wire [31:0] _EVAL_481;
  wire  _EVAL_482;
  wire  _EVAL_483;
  wire  _EVAL_484;
  wire [31:0] _EVAL_485;
  wire  _EVAL_486;
  wire  _EVAL_487;
  wire  _EVAL_488;
  wire  _EVAL_489;
  wire  _EVAL_490;
  wire  _EVAL_491;
  wire  _EVAL_494;
  wire  _EVAL_495;
  wire  _EVAL_496;
  wire  _EVAL_497;
  wire  _EVAL_498;
  wire [1:0] _EVAL_499;
  wire [31:0] _EVAL_500;
  wire  _EVAL_501;
  wire  _EVAL_502;
  wire  _EVAL_503;
  wire [2:0] _EVAL_504;
  wire  _EVAL_505;
  wire  _EVAL_506;
  wire  _EVAL_507;
  wire  _EVAL_508;
  wire  _EVAL_509;
  wire [31:0] _EVAL_510;
  wire  _EVAL_511;
  wire  _EVAL_512;
  wire  _EVAL_513;
  wire  _EVAL_514;
  wire  _EVAL_515;
  wire  _EVAL_516;
  wire  _EVAL_517;
  wire  _EVAL_518;
  wire  _EVAL_519;
  wire [31:0] _EVAL_520;
  wire  _EVAL_521;
  wire [31:0] _EVAL_522;
  wire  _EVAL_523;
  wire [4:0] _EVAL_525;
  wire [30:0] _EVAL_526;
  wire  _EVAL_527;
  wire  _EVAL_528;
  wire  _EVAL_529;
  wire  _EVAL_530;
  wire  _EVAL_531;
  wire  _EVAL_532;
  wire [31:0] _EVAL_533;
  wire  _EVAL_534;
  wire [31:0] _EVAL_535;
  wire  _EVAL_536;
  wire [31:0] _EVAL_537;
  wire  _EVAL_538;
  wire  _EVAL_539;
  wire  _EVAL_540;
  wire [31:0] _EVAL_541;
  wire  _EVAL_542;
  wire  _EVAL_543;
  wire  _EVAL_544;
  wire  _EVAL_545;
  wire [31:0] _EVAL_546;
  wire [31:0] _EVAL_547;
  wire  _EVAL_548;
  wire  _EVAL_549;
  wire  _EVAL_550;
  wire  _EVAL_551;
  wire  _EVAL_552;
  wire  _EVAL_553;
  wire [29:0] _EVAL_554;
  wire [31:0] _EVAL_555;
  wire  _EVAL_556;
  wire  _EVAL_557;
  wire  _EVAL_558;
  wire  _EVAL_559;
  wire [7:0] _EVAL_560;
  wire [3:0] _EVAL_561;
  wire  _EVAL_562;
  wire  _EVAL_563;
  wire  _EVAL_564;
  wire  _EVAL_566;
  wire  _EVAL_567;
  wire  _EVAL_568;
  wire  _EVAL_570;
  wire  _EVAL_572;
  wire [23:0] _EVAL_573;
  wire  _EVAL_574;
  wire  _EVAL_575;
  wire  _EVAL_576;
  wire  _EVAL_577;
  wire  _EVAL_578;
  wire  _EVAL_579;
  wire  _EVAL_580;
  wire  _EVAL_581;
  wire  _EVAL_582;
  wire [3:0] _EVAL_583;
  wire  _EVAL_584;
  wire  _EVAL_585;
  wire [15:0] _EVAL_586;
  wire  _EVAL_587;
  wire  _EVAL_588;
  wire  _EVAL_589;
  wire  _EVAL_590;
  wire [3:0] _EVAL_591;
  wire  _EVAL_593;
  wire  _EVAL_594;
  wire  _EVAL_595;
  wire  _EVAL_596;
  wire [31:0] _EVAL_597;
  wire  _EVAL_598;
  wire  _EVAL_599;
  wire  _EVAL_600;
  wire  _EVAL_601;
  wire [4:0] _EVAL_602;
  wire  _EVAL_603;
  wire  _EVAL_604;
  wire  _EVAL_605;
  wire  _EVAL_606;
  wire  _EVAL_607;
  wire  _EVAL_608;
  wire  _EVAL_609;
  wire [15:0] _EVAL_610;
  wire [1:0] _EVAL_611;
  wire [31:0] _EVAL_612;
  wire  _EVAL_613;
  wire  _EVAL_614;
  wire [31:0] _EVAL_615;
  wire [3:0] _EVAL_616;
  wire  _EVAL_617;
  wire [4:0] _EVAL_618;
  wire [3:0] _EVAL_619;
  wire  _EVAL_620;
  wire  _EVAL_621;
  wire [4:0] _EVAL_622;
  wire  _EVAL_623;
  wire  _EVAL_624;
  wire  _EVAL_625;
  wire [31:0] _EVAL_626;
  wire  _EVAL_627;
  wire  _EVAL_628;
  wire  _EVAL_629;
  wire  _EVAL_630;
  wire [3:0] _EVAL_631;
  wire  _EVAL_632;
  wire [31:0] _EVAL_633;
  reg  _EVAL_634;
  wire  _EVAL_635;
  wire [4:0] _EVAL_637;
  wire  _EVAL_638;
  wire [7:0] _EVAL_639;
  wire  _EVAL_640;
  wire [31:0] _EVAL_641;
  wire  _EVAL_642;
  wire  _EVAL_643;
  wire [1:0] _EVAL_644;
  wire  _EVAL_645;
  wire  _EVAL_646;
  wire  _EVAL_647;
  wire  _EVAL_648;
  wire [31:0] _EVAL_649;
  wire  _EVAL_650;
  wire  _EVAL_651;
  wire  _EVAL_652;
  wire  _EVAL_653;
  wire  _EVAL_655;
  wire [31:0] _EVAL_656;
  wire [23:0] _EVAL_657;
  wire  _EVAL_658;
  wire  _EVAL_660;
  wire  _EVAL_661;
  wire  _EVAL_662;
  wire [1:0] _EVAL_663;
  wire  _EVAL_664;
  wire  _EVAL_665;
  wire  _EVAL_666;
  wire  _EVAL_667;
  wire  _EVAL_668;
  wire  _EVAL_669;
  wire  _EVAL_670;
  wire  _EVAL_671;
  wire  _EVAL_672;
  wire  _EVAL_674;
  wire  _EVAL_675;
  wire  _EVAL_676;
  wire  _EVAL_677;
  wire  _EVAL_679;
  wire  _EVAL_680;
  wire  _EVAL_681;
  wire  _EVAL_682;
  wire  _EVAL_683;
  wire  _EVAL_684;
  wire  _EVAL_685;
  wire  _EVAL_686;
  wire [31:0] _EVAL_687;
  wire  _EVAL_688;
  wire  _EVAL_689;
  wire [3:0] _EVAL_690;
  wire  _EVAL_692;
  wire  _EVAL_693;
  wire  div__EVAL;
  wire  div__EVAL_0;
  wire [31:0] div__EVAL_1;
  wire  div__EVAL_2;
  wire  div__EVAL_3;
  wire [3:0] div__EVAL_4;
  wire  div__EVAL_5;
  wire [31:0] div__EVAL_6;
  wire [4:0] div__EVAL_7;
  wire [4:0] div__EVAL_8;
  wire [31:0] div__EVAL_9;
  wire  div__EVAL_10;
  wire  div__EVAL_11;
  wire [31:0] _EVAL_694;
  wire  _EVAL_695;
  wire  _EVAL_696;
  wire  _EVAL_697;
  wire [31:0] _EVAL_698;
  reg  _EVAL_699;
  wire [31:0] _EVAL_700;
  wire  _EVAL_701;
  wire [31:0] _EVAL_702;
  wire [4:0] _EVAL_703;
  wire  _EVAL_704;
  wire  _EVAL_705;
  wire  _EVAL_706;
  wire  _EVAL_707;
  wire [31:0] _EVAL_708;
  wire  _EVAL_709;
  wire  _EVAL_710;
  wire [31:0] _EVAL_711;
  wire  _EVAL_712;
  wire [31:0] _EVAL_713;
  wire  _EVAL_714;
  wire [15:0] _EVAL_716;
  wire  _EVAL_717;
  wire  _EVAL_718;
  wire  _EVAL_720;
  wire  _EVAL_721;
  wire  _EVAL_722;
  wire [9:0] _EVAL_723;
  wire  _EVAL_724;
  wire  _EVAL_725;
  wire  _EVAL_726;
  wire  _EVAL_727;
  wire [4:0] _EVAL_729;
  wire  _EVAL_730;
  wire  _EVAL_732;
  wire  _EVAL_733;
  wire [23:0] _EVAL_734;
  wire  _EVAL_735;
  wire [31:0] _EVAL_736;
  wire [31:0] _EVAL_737;
  wire [31:0] m__EVAL;
  wire [31:0] m__EVAL_0;
  wire [3:0] m__EVAL_1;
  wire  m__EVAL_2;
  wire  m__EVAL_3;
  wire  m__EVAL_4;
  wire [31:0] m__EVAL_5;
  wire  _EVAL_738;
  wire [31:0] _EVAL_740;
  wire  _EVAL_741;
  wire [31:0] _EVAL_743;
  wire  _EVAL_745;
  wire  _EVAL_746;
  wire  _EVAL_747;
  wire  _EVAL_748;
  wire  _EVAL_749;
  wire  _EVAL_750;
  wire  _EVAL_751;
  wire  _EVAL_752;
  wire  _EVAL_753;
  wire  _EVAL_754;
  wire [2:0] _EVAL_755;
  wire  _EVAL_756;
  wire  _EVAL_757;
  wire [4:0] _EVAL_758;
  wire  _EVAL_759;
  wire  _EVAL_760;
  wire  _EVAL_761;
  wire  _EVAL_762;
  wire  _EVAL_763;
  wire  _EVAL_764;
  wire [31:0] _EVAL_765;
  wire [32:0] _EVAL_766;
  wire [31:0] _EVAL_767;
  wire  _EVAL_768;
  wire  _EVAL_769;
  wire  _EVAL_770;
  wire  _EVAL_771;
  wire [1:0] _EVAL_772;
  wire  _EVAL_773;
  wire  _EVAL_774;
  wire  _EVAL_775;
  wire [31:0] _EVAL_776;
  wire  _EVAL_777;
  wire  _EVAL_778;
  wire  _EVAL_780;
  wire  _EVAL_781;
  wire  _EVAL_782;
  wire [7:0] _EVAL_783;
  wire  _EVAL_784;
  wire  _EVAL_785;
  wire [31:0] _EVAL_786;
  wire  _EVAL_787;
  wire  _EVAL_788;
  wire  _EVAL_789;
  wire [1:0] _EVAL_790;
  wire  _EVAL_791;
  wire  _EVAL_792;
  wire [29:0] _EVAL_793;
  wire  _EVAL_794;
  wire  _EVAL_795;
  wire  _EVAL_796;
  wire [4:0] _EVAL_797;
  wire  _EVAL_798;
  wire  _EVAL_800;
  wire  _EVAL_801;
  wire  _EVAL_803;
  wire  _EVAL_804;
  wire  _EVAL_805;
  wire  _EVAL_806;
  wire  _EVAL_807;
  wire  _EVAL_808;
  wire  _EVAL_810;
  wire  _EVAL_811;
  wire  _EVAL_812;
  wire [31:0] _EVAL_813;
  wire  _EVAL_814;
  wire  _EVAL_816;
  wire [31:0] _EVAL_817;
  wire  _EVAL_818;
  wire  _EVAL_819;
  wire [31:0] _EVAL_820;
  wire  _EVAL_821;
  wire  _EVAL_822;
  wire [1:0] _EVAL_824;
  wire  _EVAL_825;
  wire [31:0] _EVAL_826;
  wire  _EVAL_827;
  wire [31:0] _EVAL_828;
  wire  _EVAL_829;
  wire  _EVAL_830;
  wire [23:0] _EVAL_831;
  wire  _EVAL_833;
  wire  _EVAL_834;
  wire  _EVAL_835;
  wire  _EVAL_836;
  wire  _EVAL_837;
  wire  _EVAL_838;
  wire  _EVAL_840;
  wire [31:0] _EVAL_841;
  wire [3:0] _EVAL_842;
  wire  _EVAL_843;
  wire [31:0] _EVAL_844;
  wire  _EVAL_845;
  wire  _EVAL_846;
  wire  _EVAL_847;
  wire  _EVAL_848;
  wire  _EVAL_849;
  wire  _EVAL_850;
  wire [31:0] _EVAL_851;
  wire  _EVAL_852;
  wire  _EVAL_853;
  wire [31:0] _EVAL_854;
  wire  _EVAL_855;
  wire  _EVAL_856;
  wire  _EVAL_857;
  wire  _EVAL_858;
  wire [4:0] _EVAL_859;
  wire  _EVAL_860;
  wire  _EVAL_861;
  wire  _EVAL_862;
  wire  _EVAL_863;
  wire [31:0] _EVAL_864;
  wire  _EVAL_865;
  wire  _EVAL_866;
  wire  _EVAL_867;
  wire  _EVAL_868;
  wire  _EVAL_869;
  wire  _EVAL_870;
  wire  _EVAL_872;
  wire [5:0] _EVAL_873;
  wire  _EVAL_874;
  wire  _EVAL_875;
  wire  _EVAL_876;
  wire  _EVAL_877;
  wire  _EVAL_878;
  wire [31:0] _EVAL_879;
  wire  _EVAL_880;
  wire  _EVAL_881;
  wire  _EVAL_882;
  wire  _EVAL_883;
  wire  _EVAL_884;
  wire [31:0] _EVAL_885;
  wire [7:0] _EVAL_886;
  wire  _EVAL_887;
  wire  _EVAL_888;
  wire  _EVAL_889;
  wire  _EVAL_890;
  wire  _EVAL_891;
  wire  _EVAL_892;
  wire  _EVAL_893;
  wire [3:0] _EVAL_894;
  wire [31:0] _EVAL_895;
  wire  _EVAL_896;
  wire  _EVAL_897;
  wire [3:0] _EVAL_898;
  wire [31:0] _EVAL_899;
  wire  _EVAL_900;
  wire [3:0] _EVAL_901;
  wire [31:0] _EVAL_902;
  wire  _EVAL_903;
  wire  _EVAL_904;
  wire [31:0] _EVAL_906;
  wire [10:0] _EVAL_907;
  wire [31:0] _EVAL_908;
  wire [31:0] _EVAL_909;
  wire [10:0] _EVAL_910;
  wire  _EVAL_911;
  wire  _EVAL_912;
  wire [31:0] _EVAL_913;
  wire  _EVAL_914;
  wire  _EVAL_915;
  wire  _EVAL_916;
  wire  _EVAL_917;
  wire  _EVAL_918;
  wire  _EVAL_919;
  wire [5:0] _EVAL_920;
  wire  _EVAL_922;
  wire [31:0] _EVAL_923;
  wire  _EVAL_924;
  wire  _EVAL_925;
  wire  _EVAL_926;
  wire  _EVAL_927;
  wire [31:0] _EVAL_928;
  wire  _EVAL_929;
  wire  _EVAL_930;
  wire  _EVAL_931;
  wire  _EVAL_933;
  wire [31:0] _EVAL_934;
  wire [31:0] _EVAL_935;
  wire  _EVAL_936;
  wire  _EVAL_937;
  wire  _EVAL_940;
  wire  _EVAL_941;
  wire  _EVAL_942;
  wire  _EVAL_943;
  wire [31:0] _EVAL_944;
  wire  _EVAL_945;
  wire [31:0] _EVAL_946;
  wire  _EVAL_947;
  wire  _EVAL_948;
  wire [31:0] _EVAL_949;
  wire [1:0] _EVAL_950;
  wire  _EVAL_951;
  wire [31:0] _EVAL_952;
  wire  _EVAL_953;
  wire  _EVAL_954;
  wire  _EVAL_955;
  wire  _EVAL_956;
  wire [5:0] _EVAL_957;
  wire [31:0] _EVAL_958;
  wire [31:0] _EVAL_959;
  wire  _EVAL_961;
  wire  _EVAL_962;
  wire [31:0] _EVAL_963;
  wire  _EVAL_964;
  wire [5:0] _EVAL_965;
  wire [10:0] _EVAL_966;
  wire  _EVAL_967;
  wire [23:0] _EVAL_968;
  wire [31:0] _EVAL_969;
  wire  _EVAL_970;
  wire  _EVAL_971;
  wire  _EVAL_972;
  wire  _EVAL_973;
  wire  _EVAL_974;
  wire  _EVAL_975;
  wire  _EVAL_976;
  wire  _EVAL_978;
  wire [7:0] _EVAL_979;
  wire  _EVAL_980;
  wire  _EVAL_981;
  wire  _EVAL_982;
  wire  _EVAL_983;
  wire  _EVAL_984;
  wire  _EVAL_985;
  wire  _EVAL_986;
  wire  _EVAL_987;
  wire  _EVAL_989;
  wire  _EVAL_992;
  wire [31:0] _EVAL_993;
  wire  _EVAL_994;
  wire  _EVAL_995;
  wire  _EVAL_997;
  wire [31:0] _EVAL_998;
  wire [31:0] _EVAL_999;
  wire [31:0] _EVAL_1000;
  wire  _EVAL_1001;
  wire  _EVAL_1002;
  wire  _EVAL_1004;
  wire [31:0] _EVAL_1005;
  wire [31:0] _EVAL_1006;
  wire  _EVAL_1007;
  wire  _EVAL_1008;
  wire  _EVAL_1009;
  wire  _EVAL_1010;
  wire  _EVAL_1011;
  wire  _EVAL_1012;
  wire  _EVAL_1014;
  wire  _EVAL_1015;
  wire [3:0] _EVAL_1016;
  wire [31:0] _EVAL_1017;
  wire [3:0] _EVAL_1018;
  wire  _EVAL_1020;
  wire  _EVAL_1021;
  wire  _EVAL_1022;
  wire  _EVAL_1023;
  wire  _EVAL_1024;
  wire [31:0] _EVAL_1025;
  wire  _EVAL_1026;
  wire  _EVAL_1027;
  wire [29:0] _EVAL_1028;
  wire [3:0] _EVAL_1029;
  wire  _EVAL_1030;
  wire  _EVAL_1031;
  wire [10:0] _EVAL_1032;
  wire  _EVAL_1033;
  wire [31:0] _EVAL_1034;
  wire  _EVAL_1035;
  wire  _EVAL_1036;
  wire  _EVAL_1037;
  wire  _EVAL_1038;
  wire  _EVAL_1040;
  wire  _EVAL_1042;
  wire [31:0] _EVAL_1043;
  wire  _EVAL_1044;
  wire  _EVAL_1045;
  wire  _EVAL_1046;
  wire  _EVAL_1047;
  wire [23:0] _EVAL_1048;
  wire  _EVAL_1051;
  wire [1:0] _EVAL_1052;
  wire  _EVAL_1053;
  wire  _EVAL_1054;
  wire  _EVAL_1055;
  wire  _EVAL_1056;
  wire  _EVAL_1057;
  wire  _EVAL_1058;
  wire  _EVAL_1059;
  wire  _EVAL_1060;
  wire  _EVAL_1061;
  wire  _EVAL_1062;
  wire  _EVAL_1063;
  wire [31:0] _EVAL_1064;
  wire  _EVAL_1065;
  wire [31:0] _EVAL_1066;
  wire  _EVAL_1067;
  wire  _EVAL_1069;
  wire  _EVAL_1070;
  wire [31:0] _EVAL_1071;
  wire  _EVAL_1072;
  wire  _EVAL_1073;
  wire  _EVAL_1074;
  wire [23:0] _EVAL_1075;
  wire  _EVAL_1076;
  wire  _EVAL_1077;
  wire [31:0] _EVAL_1078;
  wire  _EVAL_1079;
  wire  _EVAL_1081;
  wire [3:0] _EVAL_1082;
  wire  _EVAL_1083;
  wire [2:0] _EVAL_1084;
  wire  _EVAL_1085;
  wire [7:0] _EVAL_1086;
  wire  _EVAL_1087;
  wire [31:0] alu__EVAL;
  wire [31:0] alu__EVAL_0;
  wire  alu__EVAL_1;
  wire [31:0] alu__EVAL_2;
  wire [3:0] alu__EVAL_3;
  wire [31:0] alu__EVAL_4;
  wire  _EVAL_1088;
  wire [31:0] _EVAL_1089;
  wire [31:0] _EVAL_1090;
  wire [7:0] _EVAL_1091;
  wire  _EVAL_1092;
  wire [31:0] _EVAL_1093;
  wire  _EVAL_1094;
  wire  _EVAL_1095;
  wire  _EVAL_1096;
  wire  _EVAL_1097;
  wire  _EVAL_1098;
  wire  _EVAL_1099;
  wire [7:0] _EVAL_1100;
  wire [31:0] _EVAL_1101;
  wire  _EVAL_1102;
  wire  _EVAL_1103;
  wire  _EVAL_1104;
  wire  _EVAL_1105;
  wire  _EVAL_1106;
  wire  _EVAL_1108;
  wire  _EVAL_1109;
  wire [31:0] _EVAL_1110;
  wire  _EVAL_1111;
  wire  _EVAL_1112;
  wire  _EVAL_1113;
  wire  _EVAL_1114;
  wire  _EVAL_1115;
  wire  _EVAL_1116;
  wire  _EVAL_1117;
  wire  _EVAL_1118;
  wire  _EVAL_1119;
  wire [31:0] _EVAL_1121;
  wire  _EVAL_1122;
  wire  _EVAL_1123;
  wire  _EVAL_1125;
  wire [31:0] _EVAL_1126;
  wire [1:0] _EVAL_1127;
  wire  ibuf__EVAL;
  wire  ibuf__EVAL_0;
  wire  ibuf__EVAL_1;
  wire  ibuf__EVAL_2;
  wire  ibuf__EVAL_3;
  wire  ibuf__EVAL_4;
  wire  ibuf__EVAL_5;
  wire  ibuf__EVAL_6;
  wire  ibuf__EVAL_7;
  wire  ibuf__EVAL_8;
  wire [4:0] ibuf__EVAL_9;
  wire  ibuf__EVAL_10;
  wire [4:0] ibuf__EVAL_11;
  wire [7:0] ibuf__EVAL_12;
  wire  ibuf__EVAL_13;
  wire [4:0] ibuf__EVAL_14;
  wire [31:0] ibuf__EVAL_15;
  wire [31:0] ibuf__EVAL_16;
  wire  ibuf__EVAL_17;
  wire [4:0] ibuf__EVAL_18;
  wire [31:0] ibuf__EVAL_19;
  wire  ibuf__EVAL_20;
  wire  ibuf__EVAL_21;
  wire  ibuf__EVAL_22;
  wire  ibuf__EVAL_23;
  wire [31:0] ibuf__EVAL_24;
  wire [4:0] ibuf__EVAL_25;
  wire  ibuf__EVAL_26;
  wire  ibuf__EVAL_27;
  wire [7:0] ibuf__EVAL_28;
  wire [31:0] ibuf__EVAL_29;
  wire  _EVAL_1128;
  wire  _EVAL_1129;
  wire  _EVAL_1130;
  wire  _EVAL_1131;
  wire  _EVAL_1132;
  wire  _EVAL_1133;
  wire  _EVAL_1134;
  wire  _EVAL_1135;
  wire  _EVAL_1136;
  wire  _EVAL_1137;
  wire  _EVAL_1138;
  wire  _EVAL_1139;
  wire [31:0] _EVAL_1140;
  wire [31:0] _EVAL_1141;
  wire  _EVAL_1142;
  wire  _EVAL_1143;
  wire  _EVAL_1144;
  wire  _EVAL_1145;
  wire  _EVAL_1146;
  wire  _EVAL_1147;
  wire  _EVAL_1148;
  wire [31:0] _EVAL_1149;
  wire [3:0] _EVAL_1150;
  wire [31:0] _EVAL_1151;
  wire  _EVAL_1152;
  wire  _EVAL_1153;
  wire  _EVAL_1154;
  wire  _EVAL_1155;
  wire  _EVAL_1156;
  wire  _EVAL_1159;
  wire  _EVAL_1160;
  wire  _EVAL_1161;
  wire  _EVAL_1162;
  wire [31:0] _EVAL_1163;
  wire [4:0] _EVAL_1164;
  wire  _EVAL_1165;
  wire  _EVAL_1166;
  wire  _EVAL_1167;
  wire  _EVAL_1168;
  wire  _EVAL_1170;
  wire  _EVAL_1171;
  wire  _EVAL_1172;
  wire [31:0] _EVAL_1174;
  wire  _EVAL_1175;
  wire  _EVAL_1176;
  wire  _EVAL_1177;
  wire  _EVAL_1178;
  wire  _EVAL_1180;
  wire  _EVAL_1181;
  wire [4:0] _EVAL_1182;
  wire  _EVAL_1184;
  wire  _EVAL_1185;
  wire  _EVAL_1186;
  wire  _EVAL_1187;
  wire  _EVAL_1188;
  wire  _EVAL_1189;
  wire  _EVAL_1190;
  wire  _EVAL_1191;
  wire [31:0] _EVAL_1192;
  wire  _EVAL_1193;
  wire  _EVAL_1195;
  wire [4:0] _EVAL_1196;
  wire  _EVAL_1197;
  wire [31:0] _EVAL_1198;
  wire  _EVAL_1199;
  wire [31:0] _EVAL_1200;
  wire  _EVAL_1201;
  wire  _EVAL_1202;
  wire  _EVAL_1203;
  wire  _EVAL_1204;
  wire  _EVAL_1205;
  wire  _EVAL_1207;
  wire  _EVAL_1208;
  wire  _EVAL_1209;
  wire  _EVAL_1211;
  wire  _EVAL_1212;
  wire  _EVAL_1213;
  wire [31:0] _EVAL_1214;
  wire  _EVAL_1215;
  wire  _EVAL_1216;
  wire  _EVAL_1217;
  wire [31:0] _EVAL_1218;
  wire  _EVAL_1219;
  wire  _EVAL_1220;
  wire  _EVAL_1221;
  wire  _EVAL_1222;
  wire [2:0] _EVAL_1223;
  wire  _EVAL_1224;
  wire  _EVAL_1225;
  wire  _EVAL_1226;
  wire [23:0] _EVAL_1227;
  wire  _EVAL_1228;
  wire  _EVAL_1229;
  wire [31:0] _EVAL_1230;
  reg [31:0] _EVAL_1231 [0:30];
  wire [31:0] _EVAL_1231__EVAL_1232_data;
  wire [4:0] _EVAL_1231__EVAL_1232_addr;
  wire [31:0] _EVAL_1231__EVAL_1233_data;
  wire [4:0] _EVAL_1231__EVAL_1233_addr;
  wire [31:0] _EVAL_1231__EVAL_1234_data;
  wire [4:0] _EVAL_1231__EVAL_1234_addr;
  wire  _EVAL_1231__EVAL_1234_mask;
  wire  _EVAL_1231__EVAL_1234_en;
  wire  _EVAL_1236;
  wire  _EVAL_1237;
  wire  _EVAL_1238;
  wire  _EVAL_1239;
  wire [1:0] _EVAL_1240;
  wire  _EVAL_1241;
  wire  _EVAL_1242;
  wire  _EVAL_1243;
  wire  _EVAL_1244;
  wire  _EVAL_1245;
  wire  _EVAL_1246;
  wire [31:0] _EVAL_1247;
  wire  _EVAL_1248;
  wire  _EVAL_1249;
  wire  _EVAL_1251;
  wire  _EVAL_1252;
  wire  _EVAL_1253;
  wire  _EVAL_1254;
  wire  _EVAL_1255;
  wire  _EVAL_1256;
  wire  _EVAL_1257;
  wire  _EVAL_1258;
  wire  _EVAL_1260;
  wire [4:0] _EVAL_1261;
  wire  _EVAL_1262;
  wire  _EVAL_1263;
  wire [3:0] _EVAL_1264;
  wire  _EVAL_1265;
  wire  _EVAL_1266;
  wire  _EVAL_1267;
  wire  _EVAL_1268;
  wire  _EVAL_1269;
  wire [31:0] _EVAL_1270;
  wire  _EVAL_1271;
  wire  _EVAL_1272;
  wire  _EVAL_1273;
  wire  _EVAL_1274;
  wire  _EVAL_1275;
  wire  _EVAL_1276;
  wire [31:0] _EVAL_1278;
  wire  _EVAL_1279;
  wire [7:0] _EVAL_1280;
  wire  _EVAL_1281;
  wire  _EVAL_1282;
  wire  _EVAL_1284;
  wire  _EVAL_1285;
  wire  _EVAL_1286;
  wire [3:0] _EVAL_1287;
  wire [10:0] _EVAL_1288;
  wire  _EVAL_1289;
  wire  _EVAL_1290;
  wire  _EVAL_1292;
  wire [4:0] _EVAL_1294;
  wire  _EVAL_1295;
  wire  _EVAL_1296;
  wire  _EVAL_1297;
  wire  _EVAL_1298;
  wire  _EVAL_1300;
  wire  _EVAL_1301;
  wire  _EVAL_1302;
  wire  _EVAL_1303;
  wire  _EVAL_1304;
  wire  _EVAL_1305;
  wire  _EVAL_1306;
  wire  _EVAL_1307;
  wire  _EVAL_1308;
  wire [31:0] _EVAL_1309;
  wire  _EVAL_1310;
  wire  _EVAL_1311;
  wire  _EVAL_1312;
  wire  _EVAL_1313;
  wire  _EVAL_1314;
  wire  _EVAL_1315;
  wire  _EVAL_1316;
  wire  _EVAL_1317;
  wire  _EVAL_1319;
  wire [1:0] _EVAL_1320;
  wire  _EVAL_1321;
  wire  _EVAL_1322;
  wire  _EVAL_1323;
  wire  _EVAL_1324;
  wire  gated_clock_rocket_clock_gate_in;
  wire  gated_clock_rocket_clock_gate_test_en;
  wire  gated_clock_rocket_clock_gate_en;
  wire  gated_clock_rocket_clock_gate_out;
  reg [31:0] _EVAL_1325;
  reg  _EVAL_1326;
  reg [2:0] _EVAL_1327;
  reg [7:0] _EVAL_1328;
  reg [31:0] _EVAL_1329;
  reg  _EVAL_1330;
  reg [31:0] _EVAL_1331;
  reg [31:0] _EVAL_1332;
  reg  _EVAL_1333;
  reg  _EVAL_1334;
  reg [2:0] _EVAL_1335;
  reg [29:0] _EVAL_1336;
  reg [4:0] _EVAL_1337;
  reg  _EVAL_1338;
  reg  _EVAL_1339;
  reg [2:0] _EVAL_1340;
  reg  _EVAL_1341;
  reg  _EVAL_1342;
  reg  _EVAL_1343;
  reg  _EVAL_1344;
  reg [31:0] _EVAL_1345;
  reg  _EVAL_1346;
  reg [31:0] _EVAL_1347;
  reg  _EVAL_1348;
  reg  _EVAL_1349;
  reg [31:0] _EVAL_1350;
  reg  _EVAL_1351;
  reg  _EVAL_1352;
  reg  _EVAL_1353;
  reg  _EVAL_1354;
  reg  _EVAL_1355;
  reg [31:0] _EVAL_1356;
  reg  _EVAL_1357;
  reg [1:0] _EVAL_1358;
  reg  _EVAL_1359;
  reg [31:0] _EVAL_1360;
  reg  _EVAL_1361;
  reg  _EVAL_1362;
  reg  _EVAL_1363;
  reg [31:0] _EVAL_1364;
  reg [4:0] _EVAL_1365;
  reg  _EVAL_1366;
  reg  _EVAL_1367;
  reg  _EVAL_1368;
  reg  _EVAL_1369;
  reg [1:0] _EVAL_1370;
  reg  _EVAL_1371;
  reg  _EVAL_1372;
  reg  _EVAL_1373;
  reg  _EVAL_1374;
  reg  _EVAL_1375;
  reg [3:0] _EVAL_1376;
  reg [31:0] _EVAL_1377;
  reg  _EVAL_1378;
  reg  _EVAL_1379;
  reg  _EVAL_1380;
  reg  _EVAL_1381;
  reg  _EVAL_1383;
  reg [4:0] _EVAL_1384;
  reg [1:0] _EVAL_1386;
  reg  _EVAL_1387;
  reg  _EVAL_1388;
  reg  _EVAL_1390;
  reg  _EVAL_1391;
  reg  _EVAL_1392;
  reg  _EVAL_1393;
  reg  _EVAL_1394;
  reg  _EVAL_1395;
  reg  _EVAL_1397;
  reg [31:0] _EVAL_1398;
  reg [1:0] _EVAL_1399;
  reg [29:0] _EVAL_1400;
  reg [31:0] _EVAL_1401;
  reg [31:0] _EVAL_1402;
  reg [2:0] _EVAL_1403;
  reg [31:0] _EVAL_1404;
  reg  _EVAL_1405;
  reg  _EVAL_1406;
  reg  _EVAL_1407;
  reg  _EVAL_1409;
  reg  _EVAL_1410;
  reg  _EVAL_1411;
  reg  _EVAL_1412;
  reg [1:0] _EVAL_1413;
  reg [31:0] _EVAL_1414;
  reg  _EVAL_1415;
  reg  _EVAL_1416;
  reg [31:0] _EVAL_1417;
  reg [31:0] _EVAL_1418;
  reg [31:0] _EVAL_1419;
  reg  _EVAL_1420;
  reg  _EVAL_1421;
  reg  _EVAL_1422;
  reg [7:0] _EVAL_1423;
  reg [31:0] _EVAL_1424;
  reg  _EVAL_1425;
  wire  _EVAL_1426;
  _EVAL_128 bpu (
    ._EVAL(bpu__EVAL),
    ._EVAL_0(bpu__EVAL_0),
    ._EVAL_1(bpu__EVAL_1),
    ._EVAL_2(bpu__EVAL_2),
    ._EVAL_3(bpu__EVAL_3),
    ._EVAL_4(bpu__EVAL_4),
    ._EVAL_5(bpu__EVAL_5),
    ._EVAL_6(bpu__EVAL_6),
    ._EVAL_7(bpu__EVAL_7),
    ._EVAL_8(bpu__EVAL_8),
    ._EVAL_9(bpu__EVAL_9),
    ._EVAL_10(bpu__EVAL_10),
    ._EVAL_11(bpu__EVAL_11),
    ._EVAL_12(bpu__EVAL_12),
    ._EVAL_13(bpu__EVAL_13),
    ._EVAL_14(bpu__EVAL_14),
    ._EVAL_15(bpu__EVAL_15),
    ._EVAL_16(bpu__EVAL_16),
    ._EVAL_17(bpu__EVAL_17),
    ._EVAL_18(bpu__EVAL_18),
    ._EVAL_19(bpu__EVAL_19),
    ._EVAL_20(bpu__EVAL_20),
    ._EVAL_21(bpu__EVAL_21),
    ._EVAL_22(bpu__EVAL_22),
    ._EVAL_23(bpu__EVAL_23),
    ._EVAL_24(bpu__EVAL_24),
    ._EVAL_25(bpu__EVAL_25),
    ._EVAL_26(bpu__EVAL_26),
    ._EVAL_27(bpu__EVAL_27),
    ._EVAL_28(bpu__EVAL_28),
    ._EVAL_29(bpu__EVAL_29),
    ._EVAL_30(bpu__EVAL_30),
    ._EVAL_31(bpu__EVAL_31),
    ._EVAL_32(bpu__EVAL_32),
    ._EVAL_33(bpu__EVAL_33),
    ._EVAL_34(bpu__EVAL_34),
    ._EVAL_35(bpu__EVAL_35),
    ._EVAL_36(bpu__EVAL_36),
    ._EVAL_37(bpu__EVAL_37),
    ._EVAL_38(bpu__EVAL_38),
    ._EVAL_39(bpu__EVAL_39),
    ._EVAL_40(bpu__EVAL_40),
    ._EVAL_41(bpu__EVAL_41),
    ._EVAL_42(bpu__EVAL_42),
    ._EVAL_43(bpu__EVAL_43)
  );
  _EVAL_127 csr (
    ._EVAL(csr__EVAL),
    ._EVAL_0(csr__EVAL_0),
    ._EVAL_1(csr__EVAL_1),
    ._EVAL_2(csr__EVAL_2),
    ._EVAL_3(csr__EVAL_3),
    ._EVAL_4(csr__EVAL_4),
    ._EVAL_5(csr__EVAL_5),
    ._EVAL_6(csr__EVAL_6),
    ._EVAL_7(csr__EVAL_7),
    ._EVAL_8(csr__EVAL_8),
    ._EVAL_9(csr__EVAL_9),
    ._EVAL_10(csr__EVAL_10),
    ._EVAL_11(csr__EVAL_11),
    ._EVAL_12(csr__EVAL_12),
    ._EVAL_13(csr__EVAL_13),
    ._EVAL_14(csr__EVAL_14),
    ._EVAL_15(csr__EVAL_15),
    ._EVAL_16(csr__EVAL_16),
    ._EVAL_17(csr__EVAL_17),
    ._EVAL_18(csr__EVAL_18),
    ._EVAL_19(csr__EVAL_19),
    ._EVAL_20(csr__EVAL_20),
    ._EVAL_21(csr__EVAL_21),
    ._EVAL_22(csr__EVAL_22),
    ._EVAL_23(csr__EVAL_23),
    ._EVAL_24(csr__EVAL_24),
    ._EVAL_25(csr__EVAL_25),
    ._EVAL_26(csr__EVAL_26),
    ._EVAL_27(csr__EVAL_27),
    ._EVAL_28(csr__EVAL_28),
    ._EVAL_29(csr__EVAL_29),
    ._EVAL_30(csr__EVAL_30),
    ._EVAL_31(csr__EVAL_31),
    ._EVAL_32(csr__EVAL_32),
    ._EVAL_33(csr__EVAL_33),
    ._EVAL_34(csr__EVAL_34),
    ._EVAL_35(csr__EVAL_35),
    ._EVAL_36(csr__EVAL_36),
    ._EVAL_37(csr__EVAL_37),
    ._EVAL_38(csr__EVAL_38),
    ._EVAL_39(csr__EVAL_39),
    ._EVAL_40(csr__EVAL_40),
    ._EVAL_41(csr__EVAL_41),
    ._EVAL_42(csr__EVAL_42),
    ._EVAL_43(csr__EVAL_43),
    ._EVAL_44(csr__EVAL_44),
    ._EVAL_45(csr__EVAL_45),
    ._EVAL_46(csr__EVAL_46),
    ._EVAL_47(csr__EVAL_47),
    ._EVAL_48(csr__EVAL_48),
    ._EVAL_49(csr__EVAL_49),
    ._EVAL_50(csr__EVAL_50),
    ._EVAL_51(csr__EVAL_51),
    ._EVAL_52(csr__EVAL_52),
    ._EVAL_53(csr__EVAL_53),
    ._EVAL_54(csr__EVAL_54),
    ._EVAL_55(csr__EVAL_55),
    ._EVAL_56(csr__EVAL_56),
    ._EVAL_57(csr__EVAL_57),
    ._EVAL_58(csr__EVAL_58),
    ._EVAL_59(csr__EVAL_59),
    ._EVAL_60(csr__EVAL_60),
    ._EVAL_61(csr__EVAL_61),
    ._EVAL_62(csr__EVAL_62),
    ._EVAL_63(csr__EVAL_63),
    ._EVAL_64(csr__EVAL_64),
    ._EVAL_65(csr__EVAL_65),
    ._EVAL_66(csr__EVAL_66),
    ._EVAL_67(csr__EVAL_67),
    ._EVAL_68(csr__EVAL_68),
    ._EVAL_69(csr__EVAL_69),
    ._EVAL_70(csr__EVAL_70),
    ._EVAL_71(csr__EVAL_71),
    ._EVAL_72(csr__EVAL_72),
    ._EVAL_73(csr__EVAL_73),
    ._EVAL_74(csr__EVAL_74),
    ._EVAL_75(csr__EVAL_75),
    ._EVAL_76(csr__EVAL_76),
    ._EVAL_77(csr__EVAL_77),
    ._EVAL_78(csr__EVAL_78),
    ._EVAL_79(csr__EVAL_79),
    ._EVAL_80(csr__EVAL_80),
    ._EVAL_81(csr__EVAL_81),
    ._EVAL_82(csr__EVAL_82),
    ._EVAL_83(csr__EVAL_83),
    ._EVAL_84(csr__EVAL_84),
    ._EVAL_85(csr__EVAL_85),
    ._EVAL_86(csr__EVAL_86),
    ._EVAL_87(csr__EVAL_87),
    ._EVAL_88(csr__EVAL_88),
    ._EVAL_89(csr__EVAL_89),
    ._EVAL_90(csr__EVAL_90),
    ._EVAL_91(csr__EVAL_91),
    ._EVAL_92(csr__EVAL_92),
    ._EVAL_93(csr__EVAL_93),
    ._EVAL_94(csr__EVAL_94),
    ._EVAL_95(csr__EVAL_95),
    ._EVAL_96(csr__EVAL_96),
    ._EVAL_97(csr__EVAL_97),
    ._EVAL_98(csr__EVAL_98),
    ._EVAL_99(csr__EVAL_99),
    ._EVAL_100(csr__EVAL_100),
    ._EVAL_101(csr__EVAL_101),
    ._EVAL_102(csr__EVAL_102),
    ._EVAL_103(csr__EVAL_103),
    ._EVAL_104(csr__EVAL_104),
    ._EVAL_105(csr__EVAL_105),
    ._EVAL_106(csr__EVAL_106),
    ._EVAL_107(csr__EVAL_107),
    ._EVAL_108(csr__EVAL_108),
    ._EVAL_109(csr__EVAL_109),
    ._EVAL_110(csr__EVAL_110),
    ._EVAL_111(csr__EVAL_111),
    ._EVAL_112(csr__EVAL_112),
    ._EVAL_113(csr__EVAL_113),
    ._EVAL_114(csr__EVAL_114),
    ._EVAL_115(csr__EVAL_115),
    ._EVAL_116(csr__EVAL_116),
    ._EVAL_117(csr__EVAL_117),
    ._EVAL_118(csr__EVAL_118),
    ._EVAL_119(csr__EVAL_119),
    ._EVAL_120(csr__EVAL_120),
    ._EVAL_121(csr__EVAL_121),
    ._EVAL_122(csr__EVAL_122),
    ._EVAL_123(csr__EVAL_123),
    ._EVAL_124(csr__EVAL_124),
    ._EVAL_125(csr__EVAL_125),
    ._EVAL_126(csr__EVAL_126),
    ._EVAL_127(csr__EVAL_127),
    ._EVAL_128(csr__EVAL_128),
    ._EVAL_129(csr__EVAL_129),
    ._EVAL_130(csr__EVAL_130),
    ._EVAL_131(csr__EVAL_131),
    ._EVAL_132(csr__EVAL_132),
    ._EVAL_133(csr__EVAL_133),
    ._EVAL_134(csr__EVAL_134),
    ._EVAL_135(csr__EVAL_135),
    ._EVAL_136(csr__EVAL_136),
    ._EVAL_137(csr__EVAL_137),
    ._EVAL_138(csr__EVAL_138),
    ._EVAL_139(csr__EVAL_139),
    ._EVAL_140(csr__EVAL_140),
    ._EVAL_141(csr__EVAL_141),
    ._EVAL_142(csr__EVAL_142),
    ._EVAL_143(csr__EVAL_143),
    ._EVAL_144(csr__EVAL_144),
    ._EVAL_145(csr__EVAL_145),
    ._EVAL_146(csr__EVAL_146),
    ._EVAL_147(csr__EVAL_147),
    ._EVAL_148(csr__EVAL_148),
    ._EVAL_149(csr__EVAL_149),
    ._EVAL_150(csr__EVAL_150),
    ._EVAL_151(csr__EVAL_151),
    ._EVAL_152(csr__EVAL_152),
    ._EVAL_153(csr__EVAL_153),
    ._EVAL_154(csr__EVAL_154),
    ._EVAL_155(csr__EVAL_155),
    ._EVAL_156(csr__EVAL_156),
    ._EVAL_157(csr__EVAL_157),
    ._EVAL_158(csr__EVAL_158),
    ._EVAL_159(csr__EVAL_159),
    ._EVAL_160(csr__EVAL_160),
    ._EVAL_161(csr__EVAL_161),
    ._EVAL_162(csr__EVAL_162),
    ._EVAL_163(csr__EVAL_163),
    ._EVAL_164(csr__EVAL_164),
    ._EVAL_165(csr__EVAL_165),
    ._EVAL_166(csr__EVAL_166),
    ._EVAL_167(csr__EVAL_167),
    ._EVAL_168(csr__EVAL_168),
    ._EVAL_169(csr__EVAL_169),
    ._EVAL_170(csr__EVAL_170),
    ._EVAL_171(csr__EVAL_171),
    ._EVAL_172(csr__EVAL_172),
    ._EVAL_173(csr__EVAL_173),
    ._EVAL_174(csr__EVAL_174),
    ._EVAL_175(csr__EVAL_175),
    ._EVAL_176(csr__EVAL_176),
    ._EVAL_177(csr__EVAL_177),
    ._EVAL_178(csr__EVAL_178),
    ._EVAL_179(csr__EVAL_179),
    ._EVAL_180(csr__EVAL_180),
    ._EVAL_181(csr__EVAL_181),
    ._EVAL_182(csr__EVAL_182),
    ._EVAL_183(csr__EVAL_183),
    ._EVAL_184(csr__EVAL_184),
    ._EVAL_185(csr__EVAL_185),
    ._EVAL_186(csr__EVAL_186)
  );
  _EVAL_130 div (
    ._EVAL(div__EVAL),
    ._EVAL_0(div__EVAL_0),
    ._EVAL_1(div__EVAL_1),
    ._EVAL_2(div__EVAL_2),
    ._EVAL_3(div__EVAL_3),
    ._EVAL_4(div__EVAL_4),
    ._EVAL_5(div__EVAL_5),
    ._EVAL_6(div__EVAL_6),
    ._EVAL_7(div__EVAL_7),
    ._EVAL_8(div__EVAL_8),
    ._EVAL_9(div__EVAL_9),
    ._EVAL_10(div__EVAL_10),
    ._EVAL_11(div__EVAL_11)
  );
  _EVAL_131 m (
    ._EVAL(m__EVAL),
    ._EVAL_0(m__EVAL_0),
    ._EVAL_1(m__EVAL_1),
    ._EVAL_2(m__EVAL_2),
    ._EVAL_3(m__EVAL_3),
    ._EVAL_4(m__EVAL_4),
    ._EVAL_5(m__EVAL_5)
  );
  _EVAL_129 alu (
    ._EVAL(alu__EVAL),
    ._EVAL_0(alu__EVAL_0),
    ._EVAL_1(alu__EVAL_1),
    ._EVAL_2(alu__EVAL_2),
    ._EVAL_3(alu__EVAL_3),
    ._EVAL_4(alu__EVAL_4)
  );
  _EVAL_126 ibuf (
    ._EVAL(ibuf__EVAL),
    ._EVAL_0(ibuf__EVAL_0),
    ._EVAL_1(ibuf__EVAL_1),
    ._EVAL_2(ibuf__EVAL_2),
    ._EVAL_3(ibuf__EVAL_3),
    ._EVAL_4(ibuf__EVAL_4),
    ._EVAL_5(ibuf__EVAL_5),
    ._EVAL_6(ibuf__EVAL_6),
    ._EVAL_7(ibuf__EVAL_7),
    ._EVAL_8(ibuf__EVAL_8),
    ._EVAL_9(ibuf__EVAL_9),
    ._EVAL_10(ibuf__EVAL_10),
    ._EVAL_11(ibuf__EVAL_11),
    ._EVAL_12(ibuf__EVAL_12),
    ._EVAL_13(ibuf__EVAL_13),
    ._EVAL_14(ibuf__EVAL_14),
    ._EVAL_15(ibuf__EVAL_15),
    ._EVAL_16(ibuf__EVAL_16),
    ._EVAL_17(ibuf__EVAL_17),
    ._EVAL_18(ibuf__EVAL_18),
    ._EVAL_19(ibuf__EVAL_19),
    ._EVAL_20(ibuf__EVAL_20),
    ._EVAL_21(ibuf__EVAL_21),
    ._EVAL_22(ibuf__EVAL_22),
    ._EVAL_23(ibuf__EVAL_23),
    ._EVAL_24(ibuf__EVAL_24),
    ._EVAL_25(ibuf__EVAL_25),
    ._EVAL_26(ibuf__EVAL_26),
    ._EVAL_27(ibuf__EVAL_27),
    ._EVAL_28(ibuf__EVAL_28),
    ._EVAL_29(ibuf__EVAL_29)
  );
  EICG_wrapper gated_clock_rocket_clock_gate (
    .in(gated_clock_rocket_clock_gate_in),
    .test_en(gated_clock_rocket_clock_gate_test_en),
    .en(gated_clock_rocket_clock_gate_en),
    .out(gated_clock_rocket_clock_gate_out)
  );
  assign _EVAL_1231__EVAL_1232_addr = ~_EVAL_1261;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _EVAL_1231__EVAL_1232_data = _EVAL_1231[_EVAL_1231__EVAL_1232_addr];
  `else
  assign _EVAL_1231__EVAL_1232_data = _EVAL_1231__EVAL_1232_addr >= 5'h1f ? _RAND_5[31:0] :
    _EVAL_1231[_EVAL_1231__EVAL_1232_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _EVAL_1231__EVAL_1233_addr = ~_EVAL_859;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _EVAL_1231__EVAL_1233_data = _EVAL_1231[_EVAL_1231__EVAL_1233_addr];
  `else
  assign _EVAL_1231__EVAL_1233_data = _EVAL_1231__EVAL_1233_addr >= 5'h1f ? _RAND_6[31:0] :
    _EVAL_1231[_EVAL_1231__EVAL_1233_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _EVAL_1231__EVAL_1234_data = _EVAL_1130 ? _EVAL_1 : _EVAL_1090;
  assign _EVAL_1231__EVAL_1234_addr = ~_EVAL_1182;
  assign _EVAL_1231__EVAL_1234_mask = 1'h1;
  assign _EVAL_1231__EVAL_1234_en = _EVAL_668 & _EVAL_428;
  assign _EVAL = csr__EVAL_150;
  assign _EVAL_983 = _EVAL_374 | _EVAL_890;
  assign _EVAL_193 = _EVAL_954 | _EVAL_961;
  assign _EVAL_259 = ~_EVAL_712;
  assign _EVAL_668 = _EVAL_1067 | _EVAL_627;
  assign _EVAL_1062 = _EVAL_927 & _EVAL_83;
  assign _EVAL_622 = _EVAL_2[5:1];
  assign _EVAL_1252 = _EVAL_1417[31];
  assign _EVAL_29 = _EVAL_975 ? csr__EVAL_161 : _EVAL_407;
  assign _EVAL_1279 = _EVAL_322 == 32'h2013;
  assign bpu__EVAL_21 = csr__EVAL_169;
  assign _EVAL_1323 = _EVAL_308 | _EVAL_1021;
  assign _EVAL_1083 = _EVAL_1391 & _EVAL_1246;
  assign _EVAL_959 = _EVAL_1356;
  assign ibuf__EVAL_2 = _EVAL_158;
  assign div__EVAL_9 = _EVAL_1415 ? _EVAL_1066 : _EVAL_998;
  assign _EVAL_751 = _EVAL_1327 == 3'h2;
  assign _EVAL_767 = ibuf__EVAL_19 & 32'h1058;
  assign _EVAL_371 = _EVAL_1070 | csr__EVAL_168;
  assign _EVAL_1162 = _EVAL_1261 == _EVAL_181;
  assign _EVAL_1214 = ~_EVAL_1192;
  assign csr__EVAL_135 = _EVAL_135;
  assign _EVAL_1007 = _EVAL_1111 | _EVAL_1104;
  assign _EVAL_1016 = ibuf__EVAL_6 ? 4'h1 : _EVAL_901;
  assign _EVAL_685 = _EVAL_311 | _EVAL_442;
  assign _EVAL_911 = _EVAL_1375 & _EVAL_1330;
  assign _EVAL_575 = _EVAL_643 | _EVAL_1191;
  assign _EVAL_947 = _EVAL_946 == 32'h6033;
  assign _EVAL_816 = _EVAL_510 == 32'h0;
  assign _EVAL_961 = _EVAL_1337 == 5'hb;
  assign _EVAL_514 = _EVAL_1374 & _EVAL_326;
  assign _EVAL_93 = csr__EVAL_170;
  assign _EVAL_1199 = _EVAL_1030 | _EVAL_1292;
  assign _EVAL_445 = _EVAL_632 | _EVAL_1133;
  assign bpu__EVAL_23 = ibuf__EVAL_15;
  assign _EVAL_1076 = _EVAL_1395 & _EVAL_819;
  assign _EVAL_922 = _EVAL_494 | _EVAL_178;
  assign csr__EVAL_18 = _EVAL_3;
  assign bpu__EVAL_41 = csr__EVAL_61;
  assign _EVAL_423 = _EVAL_1125 | _EVAL_858;
  assign _EVAL_104 = csr__EVAL_116;
  assign _EVAL_252 = ~_EVAL_1195;
  assign _EVAL_850 = _EVAL_1422 & _EVAL_777;
  assign _EVAL_191 = ibuf__EVAL_19 & 32'h2004074;
  assign _EVAL_1027 = _EVAL_1403 != 3'h0;
  assign _EVAL_1125 = _EVAL_755 == 3'h6;
  assign _EVAL_805 = _EVAL_847;
  assign _EVAL_831 = _EVAL_968 & _EVAL_657;
  assign _EVAL_710 = _EVAL_767 == 32'h1040;
  assign _EVAL_1217 = _EVAL_626[0];
  assign _EVAL_1245 = _EVAL_1009 | ibuf__EVAL_27;
  assign _EVAL_1056 = _EVAL_181 == _EVAL_1261;
  assign _EVAL_417 = _EVAL_1129 | _EVAL_1316;
  assign _EVAL_313 = _EVAL_652;
  assign _EVAL_196 = _EVAL_233 | _EVAL_1113;
  assign _EVAL_1221 = _EVAL_797 != 5'h0;
  assign _EVAL_943 = _EVAL_1141 == 32'h0;
  assign _EVAL_1303 = _EVAL_256 | _EVAL_257;
  assign _EVAL_886 = _EVAL_783;
  assign _EVAL_749 = _EVAL_797 == _EVAL_525;
  assign _EVAL_1059 = |_EVAL_1075;
  assign _EVAL_187 = _EVAL_1395 & _EVAL_1148;
  assign _EVAL_223 = _EVAL_1062 ? 4'h4 : _EVAL_619;
  assign _EVAL_33 = _EVAL_1370;
  assign _EVAL_1225 = _EVAL_285 == 32'h20;
  assign _EVAL_475 = _EVAL_1311 | _EVAL_1161;
  assign _EVAL_7 = csr__EVAL_68;
  assign _EVAL_1065 = _EVAL_946 == 32'h33;
  assign _EVAL_1085 = ~_EVAL_483;
  assign _EVAL_632 = _EVAL_830 | _EVAL_289;
  assign _EVAL_714 = _EVAL_390 | ibuf__EVAL_6;
  assign _EVAL_629 = _EVAL_1020 & _EVAL_1085;
  assign _EVAL_486 = _EVAL_556 & _EVAL_605;
  assign _EVAL_590 = _EVAL_322 == 32'h3073;
  assign _EVAL_861 = _EVAL_548 | _EVAL_852;
  assign m__EVAL_3 = _EVAL_74;
  assign _EVAL_495 = _EVAL_879 == 32'ha000202f;
  assign _EVAL_528 = _EVAL_757 | _EVAL_507;
  assign _EVAL_317 = _EVAL_841 == 32'h4;
  assign _EVAL_847 = _EVAL_1207 ? $signed(1'sh0) : $signed(_EVAL_1226);
  assign _EVAL_409 = _EVAL_1199 | csr__EVAL_115;
  assign _EVAL_1140 = {_EVAL_526, 1'h0};
  assign _EVAL_681 = _EVAL_628 | _EVAL_753;
  assign _EVAL_1426 = _EVAL_801 | _EVAL_943;
  assign _EVAL_355 = ibuf__EVAL_19 & 32'h6018;
  assign _EVAL_679 = _EVAL_984 | _EVAL_1301;
  assign _EVAL_662 = _EVAL_841 == 32'h3;
  assign _EVAL_757 = _EVAL_384 | _EVAL_424;
  assign ibuf__EVAL_14 = _EVAL_45;
  assign _EVAL_1316 = _EVAL_934 == 32'h10;
  assign _EVAL_362 = _EVAL_191 == 32'h2000030;
  assign _EVAL_957 = {_EVAL_168,1'h0};
  assign bpu__EVAL_29 = _EVAL_1347;
  assign _EVAL_247 = _EVAL_322 == 32'h4013;
  assign _EVAL_774 = _EVAL_797 == _EVAL_168;
  assign _EVAL_120 = csr__EVAL_6;
  assign _EVAL_791 = _EVAL_361 == 32'h4040;
  assign _EVAL_389 = _EVAL_380 | _EVAL_995;
  assign _EVAL_849 = _EVAL_322 == 32'h3013;
  assign _EVAL_460 = _EVAL_1187 | _EVAL_1406;
  assign csr__EVAL_102 = _EVAL_843 | _EVAL_877;
  assign _EVAL_378 = _EVAL_529 | _EVAL_671;
  assign _EVAL_137 = csr__EVAL_99;
  assign _EVAL_810 = _EVAL_927 & _EVAL_116;
  assign _EVAL_535 = _EVAL_1130 ? _EVAL_1 : _EVAL_1090;
  assign _EVAL_987 = _EVAL_1379 & _EVAL_1037;
  assign _EVAL_203 = _EVAL_1181 | _EVAL_718;
  assign _EVAL_934 = ibuf__EVAL_19 & 32'h14;
  assign _EVAL_344 = _EVAL_1017 == 32'h4050;
  assign _EVAL_392 = _EVAL_413 | _EVAL_206;
  assign _EVAL_333 = _EVAL_1154 | _EVAL_989;
  assign _EVAL_1001 = _EVAL_1102 & _EVAL_720;
  assign _EVAL_576 = _EVAL_746 | _EVAL_434;
  assign _EVAL_305 = _EVAL_505 | _EVAL_590;
  assign _EVAL_1241 = _EVAL_392 | _EVAL_359;
  assign _EVAL_27 = csr__EVAL_97;
  assign _EVAL_496 = ibuf__EVAL_23 & _EVAL_186;
  assign _EVAL_1097 = ~_EVAL_1105;
  assign _EVAL_225 = _EVAL_656;
  assign _EVAL_240 = $signed(_EVAL_743) + $signed(_EVAL_913);
  assign _EVAL_730 = _EVAL_431 & _EVAL_1209;
  assign _EVAL_470 = _EVAL_1055 & _EVAL_1391;
  assign _EVAL_700 = ibuf__EVAL_19 & 32'h50;
  assign csr__EVAL_62 = _EVAL_117;
  assign _EVAL_1201 = _EVAL_279 | csr__EVAL_111;
  assign _EVAL_298 = _EVAL_813 == 32'h2008;
  assign _EVAL_1175 = _EVAL_196 | _EVAL_275;
  assign _EVAL_487 = _EVAL_298 & _EVAL_1045;
  assign _EVAL_75 = csr__EVAL_124;
  assign _EVAL_277 = _EVAL_946 == 32'h2006033;
  assign _EVAL_979 = _EVAL_1278[7:0];
  assign _EVAL_666 = _EVAL_928 == 32'h40;
  assign _EVAL_727 = _EVAL_463 | _EVAL_1367;
  assign _EVAL_1106 = _EVAL_1008 & _EVAL_607;
  assign csr__EVAL_121 = _EVAL_431 & _EVAL_1209;
  assign _EVAL_435 = _EVAL_633;
  assign _EVAL_1275 = _EVAL_1103 | _EVAL_943;
  assign _EVAL_1314 = _EVAL_870 | _EVAL_1326;
  assign _EVAL_775 = _EVAL_1261 != 5'h0;
  assign _EVAL_347 = _EVAL_738 | _EVAL_289;
  assign _EVAL_755 = {_EVAL_491,_EVAL_1176,_EVAL_642};
  assign bpu__EVAL_15 = csr__EVAL_39;
  assign _EVAL_303 = csr__EVAL_114 | bpu__EVAL_9;
  assign _EVAL_1224 = bpu__EVAL_2 | _EVAL_1092;
  assign _EVAL_1239 = _EVAL_1201 | _EVAL_665;
  assign _EVAL_621 = _EVAL_1426 | _EVAL_593;
  assign bpu__EVAL_27 = csr__EVAL_107;
  assign _EVAL_452 = _EVAL_703 == 5'h5;
  assign csr__EVAL_28 = {_EVAL_610,_EVAL_716};
  assign _EVAL_572 = _EVAL_782 | _EVAL_1238;
  assign div__EVAL_8 = _EVAL_1417[11:7];
  assign _EVAL_1053 = _EVAL_1337 == 5'ha;
  assign bpu__EVAL_37 = csr__EVAL_159;
  assign _EVAL_1088 = _EVAL_294 | _EVAL_251;
  assign _EVAL_613 = _EVAL_1305 | _EVAL_473;
  assign _EVAL_67 = csr__EVAL_110;
  assign _EVAL_541 = ibuf__EVAL_19 & 32'h6034;
  assign _EVAL_1144 = _EVAL_677;
  assign bpu__EVAL_4 = csr__EVAL_142;
  assign _EVAL_1004 = _EVAL_322 == 32'h13;
  assign _EVAL_320 = _EVAL_946 == 32'h5033;
  assign _EVAL_674 = _EVAL_969 == 32'h7000;
  assign _EVAL_161 = csr__EVAL_76;
  assign _EVAL_985 = _EVAL_703 == 5'h0;
  assign _EVAL_257 = _EVAL_946 == 32'h7033;
  assign _EVAL_212 = ~_EVAL_704;
  assign _EVAL_227 = _EVAL_841 == 32'hc;
  assign _EVAL_112 = ~_EVAL_164;
  assign gated_clock_rocket_clock_gate_test_en = _EVAL_154;
  assign _EVAL_1082 = _EVAL_436 ? 4'he : 4'h3;
  assign _EVAL_226 = _EVAL_1258 | _EVAL_542;
  assign _EVAL_950 = _EVAL_1407 ? 2'h0 : 2'h2;
  assign _EVAL_718 = _EVAL_238 ? 1'h0 : _EVAL_1378;
  assign _EVAL_560 = _EVAL_1086;
  assign _EVAL_605 = _EVAL_1412 | _EVAL_1083;
  assign _EVAL_649 = ibuf__EVAL_19 & 32'h18000008;
  assign _EVAL_534 = _EVAL_931 | _EVAL_304;
  assign csr__EVAL_153 = _EVAL_111;
  assign _EVAL_845 = _EVAL_530 | _EVAL_412;
  assign _EVAL_1126 = {_EVAL_805,_EVAL_1032,_EVAL_886,_EVAL_1142,_EVAL_920,_EVAL_243,_EVAL_312};
  assign _EVAL_98 = csr__EVAL_75;
  assign _EVAL_945 = _EVAL_423 & _EVAL_237;
  assign _EVAL_500 = ibuf__EVAL_19 & 32'h4004;
  assign _EVAL_624 = _EVAL_423 | _EVAL_856;
  assign bpu__EVAL_0 = csr__EVAL_128;
  assign _EVAL_1196 = _EVAL_1364[19:15];
  assign _EVAL_881 = _EVAL_997 | _EVAL_725;
  assign _EVAL_601 = _EVAL_681 | _EVAL_255;
  assign _EVAL_955 = _EVAL_686 | _EVAL_682;
  assign _EVAL_544 = _EVAL_518 & _EVAL_1097;
  assign _EVAL_814 = _EVAL_879 == 32'h800202f;
  assign _EVAL_973 = _EVAL_663 == 2'h3;
  assign _EVAL_783 = _EVAL_660 ? $signed({8{_EVAL_847}}) : $signed(_EVAL_1280);
  assign _EVAL_1031 = _EVAL_194 & _EVAL_1317;
  assign _EVAL_1073 = _EVAL_897 | _EVAL_925;
  assign _EVAL_87 = csr__EVAL_53;
  assign _EVAL_51 = alu__EVAL_4;
  assign _EVAL_319 = _EVAL_1353 | _EVAL_1422;
  assign _EVAL_763 = _EVAL_1043 == 32'h0;
  assign _EVAL_1220 = _EVAL_1121 == 32'h40000008;
  assign _EVAL_91 = 32'h0;
  assign _EVAL_769 = csr__EVAL_56[12];
  assign div__EVAL_4 = _EVAL_1376;
  assign _EVAL_310 = ibuf__EVAL_19 & 32'h7f;
  assign _EVAL_114 = csr__EVAL_3;
  assign _EVAL_1112 = _EVAL_213 | _EVAL_495;
  assign _EVAL_520 = _EVAL_1231__EVAL_1232_data;
  assign _EVAL_698 = ibuf__EVAL_19 & 32'h64;
  assign _EVAL_236 = _EVAL_469 & _EVAL_657;
  assign _EVAL_965 = {1'h0,_EVAL_42,_EVAL_18,1'h0,_EVAL_106,_EVAL_59};
  assign _EVAL_1272 = _EVAL_386 == 2'h1;
  assign _EVAL_1101 = _EVAL_914 ? _EVAL_1347 : 32'h0;
  assign _EVAL_891 = _EVAL_980 & _EVAL_1253;
  assign ibuf__EVAL_10 = _EVAL_119;
  assign _EVAL_697 = _EVAL_1255 | _EVAL_791;
  assign _EVAL_206 = _EVAL_879 == 32'he000202f;
  assign _EVAL_271 = {ibuf__EVAL_7,ibuf__EVAL_27};
  assign _EVAL_1045 = ~_EVAL_781;
  assign _EVAL_1190 = _EVAL_1413 == 2'h1;
  assign ibuf__EVAL = _EVAL_821 | _EVAL_987;
  assign _EVAL_1135 = _EVAL_242 | _EVAL_227;
  assign _EVAL_740 = ibuf__EVAL_19 & 32'h1050;
  assign _EVAL_129 = ibuf__EVAL_17;
  assign _EVAL_295 = _EVAL_612 == 32'h0;
  assign bpu__EVAL_30 = csr__EVAL_178;
  assign _EVAL_658 = ~_EVAL_821;
  assign _EVAL_548 = _EVAL_458 | _EVAL_376;
  assign _EVAL_906 = _EVAL_240[31:0];
  assign _EVAL_437 = |_EVAL_734;
  assign _EVAL_199 = |_EVAL_236;
  assign _EVAL_511 = _EVAL_927 & _EVAL_39;
  assign _EVAL_594 = _EVAL_1422 ^ _EVAL_1172;
  assign _EVAL_1165 = _EVAL_881 | _EVAL_422;
  assign _EVAL_434 = ibuf__EVAL_19 == 32'h7b200073;
  assign _EVAL_89 = csr__EVAL_123;
  assign alu__EVAL_2 = _EVAL_1163;
  assign _EVAL_1160 = _EVAL_430 | _EVAL_263;
  assign _EVAL_982 = _EVAL_369 & _EVAL_1167;
  assign _EVAL_1058 = _EVAL_322 == 32'h1023;
  assign _EVAL_610 = _EVAL_346 ? _EVAL_331 : 16'h0;
  assign _EVAL_1174 = _EVAL_246 ? _EVAL_535 : _EVAL_520;
  assign _EVAL_1168 = ibuf__EVAL_19 == 32'h30200073;
  assign _EVAL_6 = csr__EVAL_79;
  assign _EVAL_198 = _EVAL_1025;
  assign _EVAL_694 = _EVAL_1140 >> _EVAL_1261;
  assign _EVAL_771 = _EVAL_451 == 32'h2001030;
  assign _EVAL_902 = ibuf__EVAL_19 & 32'h24;
  assign _EVAL_1048 = {{14'd0}, _EVAL_723};
  assign _EVAL_633 = _EVAL_1153 ? $signed(_EVAL_1110) : $signed(_EVAL_817);
  assign _EVAL_1218 = _EVAL_1367 ? $signed(_EVAL_944) : $signed({{28{_EVAL_591[3]}},_EVAL_591});
  assign _EVAL_290 = csr__EVAL_56[2];
  assign _EVAL_1268 = _EVAL_490 | _EVAL_81;
  assign _EVAL_1294 = _EVAL_1424[19:15];
  assign _EVAL_1267 = _EVAL_1197 & _EVAL_544;
  assign _EVAL_687 = ibuf__EVAL_19 & 32'hf9f0707f;
  assign _EVAL_300 = _EVAL_1322 | _EVAL_670;
  assign _EVAL_882 = _EVAL_1337 == 5'h6;
  assign _EVAL_1285 = _EVAL_679 | _EVAL_506;
  assign _EVAL_1141 = ibuf__EVAL_19 & 32'h18;
  assign _EVAL_1266 = _EVAL_322 == 32'h7013;
  assign _EVAL_598 = csr__EVAL | _EVAL_484;
  assign _EVAL_948 = _EVAL_168 == _EVAL_1261;
  assign _EVAL_764 = _EVAL_1348 & _EVAL_1042;
  assign _EVAL_587 = _EVAL_896 | _EVAL_1095;
  assign _EVAL_123 = 1'h0;
  assign _EVAL_424 = _EVAL_522 == 32'h2004020;
  assign _EVAL_384 = _EVAL_189 | _EVAL_362;
  assign _EVAL_1099 = _EVAL_982 & _EVAL_1152;
  assign _EVAL_1024 = _EVAL_150 & _EVAL_4;
  assign _EVAL_1313 = _EVAL_1148 & _EVAL_160;
  assign _EVAL_171 = _EVAL_761 | _EVAL_888;
  assign csr__EVAL_101 = _EVAL_614 ? _EVAL_1377 : 32'h0;
  assign _EVAL_485 = _EVAL_918 ? _EVAL_535 : _EVAL_1071;
  assign _EVAL_1046 = _EVAL_513 | _EVAL_1065;
  assign _EVAL_1180 = _EVAL_1339 != _EVAL_1334;
  assign _EVAL_1044 = _EVAL_322 == 32'h1073;
  assign _EVAL_1254 = _EVAL_765 == 32'h40;
  assign _EVAL_125 = csr__EVAL_165;
  assign _EVAL_608 = _EVAL_403 | _EVAL_395;
  assign _EVAL_712 = _EVAL_627 & _EVAL_773;
  assign _EVAL_35 = csr__EVAL_177;
  assign _EVAL_37 = csr__EVAL_54;
  assign _EVAL_136 = csr__EVAL_105;
  assign _EVAL_615 = ibuf__EVAL_19 & 32'h18000020;
  assign _EVAL_593 = _EVAL_1006 == 32'h4000;
  assign _EVAL_650 = _EVAL_547 == 32'h48;
  assign _EVAL_878 = _EVAL_1416 | _EVAL_994;
  assign _EVAL_661 = _EVAL_454 & _EVAL_948;
  assign _EVAL_671 = _EVAL_700 == 32'h0;
  assign _EVAL_603 = _EVAL_870 | _EVAL_1363;
  assign bpu__EVAL_12 = csr__EVAL_22;
  assign _EVAL_925 = _EVAL_1379 & _EVAL_1172;
  assign _EVAL_910 = _EVAL_907;
  assign _EVAL_656 = $signed(_EVAL_466) & -32'sh2;
  assign _EVAL_359 = _EVAL_687 == 32'h1000202f;
  assign _EVAL_1265 = _EVAL_377;
  assign bpu__EVAL_42 = csr__EVAL_100;
  assign _EVAL_531 = _EVAL_1374 | _EVAL_1344;
  assign _EVAL_413 = _EVAL_803 | _EVAL_495;
  assign _EVAL_1256 = _EVAL_295 | _EVAL_1166;
  assign _EVAL_489 = _EVAL_584 | _EVAL_596;
  assign _EVAL_856 = _EVAL_755 == 3'h5;
  assign csr__EVAL_27 = _EVAL_113;
  assign _EVAL_309 = _EVAL_729 == _EVAL_797;
  assign ibuf__EVAL_0 = _EVAL_107;
  assign _EVAL_494 = _EVAL_699 | _EVAL_287;
  assign _EVAL_381 = ~_EVAL_1147;
  assign _EVAL_397 = _EVAL_859 != 5'h0;
  assign _EVAL_1290 = _EVAL_835 | _EVAL_1061;
  assign _EVAL_264 = _EVAL_1417[19:12];
  assign _EVAL_1187 = _EVAL_342 | _EVAL_1395;
  assign _EVAL_711 = ibuf__EVAL_19 & 32'h3054;
  assign _EVAL_644 = ibuf__EVAL_19[13:12];
  assign _EVAL_502 = _EVAL_981 | _EVAL_1351;
  assign _EVAL_508 = _EVAL_841 == 32'h1;
  assign _EVAL_410 = _EVAL_956;
  assign _EVAL_1060 = _EVAL_880 | _EVAL_1081;
  assign _EVAL_130 = _EVAL_634;
  assign _EVAL_156 = csr__EVAL_87;
  assign _EVAL_282 = _EVAL_1228 | ibuf__EVAL_4;
  assign _EVAL_462 = _EVAL_1306 | _EVAL_849;
  assign _EVAL_387 = _EVAL_166 == 32'h20;
  assign _EVAL_9 = _EVAL_1337;
  assign _EVAL_457 = _EVAL_281 | _EVAL_1211;
  assign _EVAL_450 = _EVAL_1099 ? 2'h2 : 2'h3;
  assign _EVAL_778 = _EVAL_322 == 32'h2073;
  assign _EVAL_631 = _EVAL_511 ? 4'hd : {{1'd0}, _EVAL_1223};
  assign _EVAL_483 = _EVAL_2[0];
  assign _EVAL_1026 = _EVAL_1046 | _EVAL_926;
  assign _EVAL_1297 = _EVAL_804 | _EVAL_1106;
  assign _EVAL_167 = _EVAL_1333 ? _EVAL_963 : _EVAL_1230;
  assign csr__EVAL_73 = _EVAL_1377;
  assign _EVAL_262 = _EVAL_994 ? 4'h6 : _EVAL_223;
  assign _EVAL_635 = _EVAL_580 | _EVAL_1307;
  assign _EVAL_279 = _EVAL_602 == 5'h0;
  assign _EVAL_1212 = _EVAL_1177 | _EVAL_857;
  assign _EVAL_796 = _EVAL_1229 | _EVAL_588;
  assign _EVAL_683 = _EVAL_1007 | _EVAL_487;
  assign _EVAL_818 = _EVAL_1138 & _EVAL_1242;
  assign _EVAL_478 = ibuf__EVAL_19 & 32'h40003054;
  assign _EVAL_863 = _EVAL_280 == 4'h0;
  assign _EVAL_52 = _EVAL_1339;
  assign _EVAL_243 = _EVAL_751 ? 4'h0 : _EVAL_894;
  assign _EVAL_1264 = _EVAL_925 ? 4'h0 : _EVAL_1082;
  assign _EVAL_1274 = _EVAL_808 | _EVAL_1051;
  assign _EVAL_760 = _EVAL_685 | _EVAL_1222;
  assign _EVAL_581 = _EVAL_1197 & _EVAL_1162;
  assign csr__EVAL_151 = _EVAL_1364[31:20];
  assign _EVAL_1311 = _EVAL_703 == 5'h4;
  assign _EVAL_843 = _EVAL_551 | _EVAL_810;
  assign _EVAL_1288 = {_EVAL_424,_EVAL_362,_EVAL_1129,_EVAL_650,_EVAL_666,_EVAL_1031,_EVAL_345};
  assign _EVAL_936 = _EVAL_627 & _EVAL_309;
  assign _EVAL_811 = _EVAL_1205 | _EVAL_674;
  assign _EVAL_879 = ibuf__EVAL_19 & 32'hf800707f;
  assign _EVAL_568 = _EVAL_702 == 32'h2010;
  assign bpu__EVAL_22 = csr__EVAL_91;
  assign _EVAL_432 = _EVAL_209 == 32'h2010;
  assign _EVAL_853 = _EVAL_181[0];
  assign _EVAL_185 = _EVAL_273 ? 2'h2 : 2'h3;
  assign _EVAL_570 = ~_EVAL_1374;
  assign _EVAL_1018 = _EVAL_1417[11:8];
  assign _EVAL_686 = _EVAL_1185 | _EVAL_1368;
  assign _EVAL_873 = _EVAL_1417[30:25];
  assign _EVAL_369 = _EVAL_1379 & _EVAL_1348;
  assign _EVAL_986 = _EVAL_841 == 32'h5;
  assign _EVAL_509 = _EVAL_946 == 32'h2003033;
  assign _EVAL_246 = _EVAL_1182 == _EVAL_1261;
  assign _EVAL_532 = _EVAL_298 & _EVAL_1282;
  assign _EVAL_707 = _EVAL_816 | _EVAL_1213;
  assign _EVAL_828 = ibuf__EVAL_19 & 32'h20;
  assign _EVAL_651 = _EVAL_541 == 32'h2010;
  assign _EVAL_338 = _EVAL_987 & _EVAL_1037;
  assign _EVAL_609 = _EVAL_1254 | _EVAL_741;
  assign _EVAL_1298 = _EVAL_713 != ibuf__EVAL_15;
  assign _EVAL_812 = _EVAL_1395 & _EVAL_1079;
  assign _EVAL_482 = _EVAL_386 == 2'h3;
  assign _EVAL_1008 = _EVAL_1138 & _EVAL_397;
  assign _EVAL_345 = {_EVAL_507,_EVAL_800,_EVAL_866,_EVAL_1014,1'h0};
  assign _EVAL_1247 = ibuf__EVAL_19 & 32'h1048;
  assign bpu__EVAL_26 = csr__EVAL_182;
  assign _EVAL_1145 = _EVAL_1337 == 5'hf;
  assign _EVAL_507 = _EVAL_755 != 3'h0;
  assign _EVAL_202 = _EVAL_1216 | _EVAL_1203;
  assign _EVAL_1244 = _EVAL_1297 | _EVAL_964;
  assign _EVAL_175 = _EVAL_190 | _EVAL_768;
  assign _EVAL_702 = ibuf__EVAL_19 & 32'h2010;
  assign _EVAL_639 = _EVAL_560;
  assign _EVAL_1119 = |_EVAL_271;
  assign _EVAL_16 = 4'h0;
  assign _EVAL_26 = csr__EVAL_13;
  assign _EVAL_1067 = _EVAL_730 & _EVAL_1420;
  assign _EVAL_407 = _EVAL_951 ? _EVAL_1401 : _EVAL_713;
  assign div__EVAL_3 = _EVAL_1374 & _EVAL_1410;
  assign _EVAL_1127 = _EVAL_899[1:0];
  assign _EVAL_281 = _EVAL_608 | _EVAL_595;
  assign _EVAL_1150 = _EVAL_1417[24:21];
  assign _EVAL_1309 = ibuf__EVAL_23 ? {{16'd0}, _EVAL_586} : ibuf__EVAL_29;
  assign _EVAL_372 = _EVAL_1207 ? _EVAL_1029 : _EVAL_1150;
  assign _EVAL_197 = _EVAL_1008 & _EVAL_794;
  assign _EVAL_390 = _EVAL_229 | ibuf__EVAL_26;
  assign _EVAL_967 = _EVAL_1267 | _EVAL_370;
  assign _EVAL_846 = _EVAL_188 | _EVAL_1211;
  assign csr__EVAL_45 = _EVAL_157;
  assign _EVAL_339 = _EVAL_1278[15:0];
  assign _EVAL_566 = _EVAL_328 | _EVAL_1310;
  assign _EVAL_703 = {1'h0,_EVAL_357,_EVAL_861,_EVAL_318,_EVAL_834};
  assign _EVAL_356 = _EVAL_946 == 32'h2001033;
  assign _EVAL_842 = bpu__EVAL_9 ? 4'he : _EVAL_583;
  assign _EVAL_758 = _EVAL_1364[24:20];
  assign _EVAL_1040 = div__EVAL_10 & div__EVAL_11;
  assign _EVAL_1011 = ~_EVAL_57;
  assign _EVAL_647 = ~_EVAL_212;
  assign _EVAL_1230 = {_EVAL_1400,_EVAL_1358};
  assign bpu__EVAL_38 = csr__EVAL_16;
  assign _EVAL_401 = _EVAL_879 == 32'hc000202f;
  assign _EVAL_1178 = _EVAL_860 | _EVAL_268;
  assign _EVAL_451 = ibuf__EVAL_19 & 32'h2001074;
  assign _EVAL_374 = _EVAL_827 | _EVAL_1099;
  assign _EVAL_168 = _EVAL_1417[11:7];
  assign _EVAL_38 = csr__EVAL_160;
  assign csr__EVAL_57 = _EVAL_63;
  assign _EVAL_258 = _EVAL_729 == _EVAL_1261;
  assign _EVAL_62 = csr__EVAL_94;
  assign csr__EVAL_23 = _EVAL_12;
  assign _EVAL_555 = _EVAL_1140 >> _EVAL_797;
  assign _EVAL_404 = _EVAL_1043 == 32'h4;
  assign _EVAL_1271 = _EVAL_788 | _EVAL_219;
  assign _EVAL_753 = _EVAL_1008 & _EVAL_174;
  assign _EVAL_537 = ibuf__EVAL_19 & 32'h2034;
  assign _EVAL_1154 = _EVAL_1271 | _EVAL_1015;
  assign _EVAL_927 = _EVAL_1375 & _EVAL_1391;
  assign _EVAL_200 = _EVAL_700 == 32'h10;
  assign _EVAL_162 = _EVAL_717 & _EVAL_449;
  assign _EVAL_302 = _EVAL_1424[31];
  assign _EVAL_803 = _EVAL_210 | _EVAL_401;
  assign _EVAL_466 = _EVAL_1422 ? $signed(_EVAL_817) : $signed(_EVAL_1110);
  assign bpu__EVAL_40 = csr__EVAL_138;
  assign _EVAL_1087 = _EVAL_829 ? $signed(1'sh0) : $signed(_EVAL_363);
  assign _EVAL_781 = csr__EVAL_56[0];
  assign _EVAL_201 = alu__EVAL;
  assign _EVAL_1151 = csr__EVAL_71;
  assign _EVAL_36 = csr__EVAL_44;
  assign _EVAL_790 = {_EVAL_397,_EVAL_775};
  assign _EVAL_1118 = ~_EVAL_1368;
  assign _EVAL_625 = _EVAL_523 | _EVAL_941;
  assign _EVAL_467 = _EVAL_968[0];
  assign _EVAL_1077 = _EVAL_841 == 32'hf;
  assign _EVAL_1226 = _EVAL_1252;
  assign _EVAL_540 = _EVAL_454 & _EVAL_1281;
  assign _EVAL_956 = _EVAL_937;
  assign _EVAL_342 = _EVAL_292 | _EVAL_1387;
  assign _EVAL_253 = _EVAL_1337 == 5'hc;
  assign _EVAL_591 = _EVAL_1407 ? $signed(4'sh2) : $signed(4'sh4);
  assign _EVAL_229 = _EVAL_303 | bpu__EVAL_2;
  assign _EVAL_1017 = ibuf__EVAL_19 & 32'h4050;
  assign _EVAL_188 = _EVAL_617 | _EVAL_595;
  assign _EVAL_1064 = _EVAL_1072 ? $signed({{28{_EVAL_898[3]}},_EVAL_898}) : $signed(_EVAL_172);
  assign _EVAL_859 = ibuf__EVAL_11;
  assign _EVAL_1306 = _EVAL_461 | _EVAL_1279;
  assign ibuf__EVAL_21 = _EVAL_149;
  assign _EVAL_220 = _EVAL_703 == 5'h7;
  assign _EVAL_1262 = _EVAL_1358 == 2'h2;
  assign bpu__EVAL_36 = csr__EVAL_112;
  assign _EVAL_981 = _EVAL_369 & _EVAL_109;
  assign _EVAL_308 = _EVAL_347 & _EVAL_405;
  assign csr__EVAL_167 = _EVAL_90;
  assign _EVAL_464 = _EVAL_1067 & _EVAL_912;
  assign _EVAL_1123 = _EVAL_215;
  assign _EVAL_1138 = _EVAL_688 | _EVAL_387;
  assign _EVAL_607 = _EVAL_859 == _EVAL_525;
  assign _EVAL_1308 = _EVAL_708 == 32'h4010;
  assign _EVAL_60 = _EVAL_1365;
  assign _EVAL_1153 = _EVAL_1118 & _EVAL_594;
  assign _EVAL_1129 = _EVAL_1034 == 32'h4;
  assign _EVAL_573 = _EVAL_968 & _EVAL_406;
  assign _EVAL_1317 = ~_EVAL_528;
  assign _EVAL_903 = _EVAL_589 | _EVAL_1122;
  assign _EVAL_498 = _EVAL_20[1];
  assign _EVAL_820 = ibuf__EVAL_19 & 32'h6044;
  assign _EVAL_892 = _EVAL_1417[14];
  assign _EVAL_299 = _EVAL_627 | _EVAL_798;
  assign _EVAL_1188 = _EVAL_1353 & _EVAL_1180;
  assign _EVAL_717 = ~_EVAL_337;
  assign _EVAL_1015 = _EVAL_322 == 32'h7063;
  assign _EVAL_545 = _EVAL_1327 == 3'h1;
  assign _EVAL_11 = csr__EVAL_89;
  assign _EVAL_773 = _EVAL_729 == _EVAL_859;
  assign _EVAL_929 = _EVAL_813 == 32'h8;
  assign bpu__EVAL_1 = csr__EVAL_81;
  assign _EVAL_953 = ~_EVAL_945;
  assign _EVAL_97 = _EVAL_1379 & _EVAL_658;
  assign _EVAL_563 = _EVAL_615 == 32'h18000020;
  assign _EVAL_1282 = ibuf__EVAL_19[25];
  assign div__EVAL = gated_clock_rocket_clock_gate_out;
  assign _EVAL_287 = _EVAL_531 | _EVAL_1362;
  assign _EVAL_1296 = csr__EVAL_155;
  assign _EVAL_326 = _EVAL_1098 | _EVAL_368;
  assign bpu__EVAL_5 = csr__EVAL_32;
  assign _EVAL_898 = _EVAL_1388 ? $signed(4'sh2) : $signed(4'sh4);
  assign _EVAL_78 = csr__EVAL_38;
  assign bpu__EVAL_20 = csr__EVAL_58;
  assign _EVAL_1164 = _EVAL_1294 & 5'h1b;
  assign _EVAL_958 = _EVAL_1140 & _EVAL_1214;
  assign _EVAL_1246 = ~_EVAL_150;
  assign csr__EVAL_49 = _EVAL_115;
  assign csr__EVAL_66 = _EVAL_100;
  assign _EVAL_1095 = csr__EVAL_181 & _EVAL_706;
  assign _EVAL_999 = _EVAL_1381 ? m__EVAL : _EVAL_1377;
  assign _EVAL_553 = _EVAL_353 | _EVAL_162;
  assign _EVAL_870 = _EVAL_1387 & csr__EVAL_2;
  assign _EVAL_705 = _EVAL_278 | _EVAL_750;
  assign _EVAL_766 = _EVAL_1402 + _EVAL_334;
  assign _EVAL_1094 = _EVAL_879 == 32'h2000202f;
  assign _EVAL_68 = csr__EVAL_24;
  assign _EVAL_817 = _EVAL_1347;
  assign _EVAL_868 = _EVAL_270 | _EVAL_752;
  assign _EVAL_1111 = ~_EVAL_202;
  assign m__EVAL_4 = gated_clock_rocket_clock_gate_out;
  assign _EVAL_567 = _EVAL_643 & _EVAL_604;
  assign _EVAL_380 = _EVAL_462 | _EVAL_1266;
  assign _EVAL_975 = _EVAL_1117 | csr__EVAL_168;
  assign _EVAL_895 = _EVAL_1345;
  assign _EVAL_386 = csr__EVAL_118[1:0];
  assign _EVAL_665 = _EVAL_821 | _EVAL_987;
  assign csr__EVAL_88 = _EVAL_122;
  assign _EVAL_1139 = _EVAL_1327 == 3'h4;
  assign _EVAL_1132 = _EVAL_646 | _EVAL_184;
  assign _EVAL_341 = _EVAL_730 & _EVAL_1355;
  assign _EVAL_1025 = csr__EVAL_70;
  assign _EVAL_855 = _EVAL_1112 | _EVAL_206;
  assign _EVAL_499 = {_EVAL_689,_EVAL_549};
  assign _EVAL_139 = _EVAL_1374 & _EVAL_1395;
  assign _EVAL_1137 = _EVAL_1027 | _EVAL_889;
  assign csr__EVAL_51 = _EVAL_84;
  assign _EVAL_251 = _EVAL_1043 == 32'h40;
  assign _EVAL_453 = _EVAL_903 | _EVAL_924;
  assign _EVAL_1149 = _EVAL_1126;
  assign _EVAL_1240 = _EVAL_661 ? 2'h1 : _EVAL_185;
  assign bpu__EVAL_31 = csr__EVAL_158;
  assign _EVAL_729 = _EVAL_629 ? _EVAL_622 : div__EVAL_7;
  assign _EVAL_725 = _EVAL_322 == 32'hf;
  assign _EVAL_1148 = ~_EVAL_85;
  assign _EVAL_772 = _EVAL_1309[1:0];
  assign _EVAL_1172 = _EVAL_186 & _EVAL_915;
  assign _EVAL_426 = ~_EVAL_324;
  assign _EVAL_1304 = _EVAL_332 | _EVAL_545;
  assign _EVAL_1029 = _EVAL_1417[19:16];
  assign _EVAL_268 = _EVAL_885 == 32'h2008;
  assign _EVAL_155 = csr__EVAL_42;
  assign _EVAL_688 = _EVAL_1225 | _EVAL_488;
  assign _EVAL_377 = _EVAL_645 & _EVAL_868;
  assign _EVAL_963 = _EVAL_231 ? _EVAL_152 : _EVAL_230;
  assign _EVAL_1116 = _EVAL_1353 & _EVAL_1339;
  assign _EVAL_1156 = _EVAL_322 == 32'h100f;
  assign _EVAL_968 = csr__EVAL_104[31:8];
  assign _EVAL_444 = {ibuf__EVAL_26,ibuf__EVAL_6};
  assign _EVAL_1176 = _EVAL_854 == 32'h2050;
  assign _EVAL_915 = _EVAL_713[1];
  assign _EVAL_692 = _EVAL_1413 == 2'h2;
  assign _EVAL_564 = _EVAL_173 | _EVAL_1276;
  assign _EVAL_726 = _EVAL_620 | _EVAL_1380;
  assign _EVAL_761 = _EVAL_1132 | _EVAL_393;
  assign _EVAL_170 = _EVAL_205 & _EVAL_1037;
  assign _EVAL_436 = _EVAL_218 | _EVAL_1260;
  assign _EVAL_984 = _EVAL_228 | _EVAL_1023;
  assign _EVAL_1051 = _EVAL_927 & _EVAL_118;
  assign _EVAL_124 = csr__EVAL_179;
  assign csr__EVAL_84 = _EVAL_31;
  assign _EVAL_735 = _EVAL_1379 & _EVAL_1249;
  assign _EVAL_394 = _EVAL_1208 | _EVAL_365;
  assign _EVAL_1223 = _EVAL_810 ? 3'h7 : 3'h5;
  assign _EVAL_1189 = _EVAL_867 | _EVAL_759;
  assign _EVAL_415 = _EVAL_795 | _EVAL_570;
  assign _EVAL_412 = _EVAL_322 == 32'h1063;
  assign csr__EVAL_63 = _EVAL_0;
  assign _EVAL_469 = csr__EVAL_118[31:8];
  assign _EVAL_190 = _EVAL_648 | _EVAL_304;
  assign _EVAL_101 = _EVAL_287 ? _EVAL_527 : _EVAL_216;
  assign _EVAL_874 = ~_EVAL_769;
  assign _EVAL_584 = _EVAL_567 | _EVAL_970;
  assign bpu__EVAL_11 = csr__EVAL_2;
  assign _EVAL_510 = ibuf__EVAL_19 & 32'h58;
  assign _EVAL_1181 = _EVAL_929 | _EVAL_732;
  assign _EVAL_283 = _EVAL_1337 == 5'h0;
  assign _EVAL_797 = ibuf__EVAL_18;
  assign _EVAL_1086 = _EVAL_1424[19:12];
  assign _EVAL_1033 = _EVAL_305 | _EVAL_825;
  assign _EVAL_907 = {11{_EVAL_677}};
  assign _EVAL_1036 = _EVAL_1417[15];
  assign _EVAL_962 = _EVAL_300 | _EVAL_1044;
  assign _EVAL_1216 = _EVAL_1033 | _EVAL_222;
  assign _EVAL_611 = _EVAL_1350[1:0];
  assign _EVAL_865 = _EVAL_478 == 32'h40001010;
  assign _EVAL_1324 = _EVAL_92;
  assign _EVAL_1055 = _EVAL_1375 & _EVAL_486;
  assign _EVAL_346 = &_EVAL_611;
  assign _EVAL_234 = _EVAL_1313 & _EVAL_747;
  assign _EVAL_713 = _EVAL_225;
  assign _EVAL_1005 = ibuf__EVAL_19 & 32'h2002074;
  assign _EVAL_667 = _EVAL_1327 != 3'h3;
  assign _EVAL_30 = csr__EVAL_148;
  assign _EVAL_273 = _EVAL_982 & _EVAL_1056;
  assign div__EVAL_2 = _EVAL_955 & _EVAL_1411;
  assign ibuf__EVAL_24 = _EVAL_72;
  assign _EVAL_1253 = _EVAL_460 | _EVAL_1410;
  assign _EVAL_458 = _EVAL_1000 == 32'h8000008;
  assign bpu__EVAL_8 = csr__EVAL_4;
  assign _EVAL_284 = _EVAL_1413 == 2'h3;
  assign _EVAL_549 = _EVAL_837 | _EVAL_943;
  assign _EVAL_876 = _EVAL_946 == 32'h40005013;
  assign csr__EVAL_10 = _EVAL_8;
  assign _EVAL_738 = _EVAL_572 | _EVAL_1058;
  assign _EVAL_597 = _EVAL_887 ? _EVAL_1089 : _EVAL_1278;
  assign _EVAL_860 = _EVAL_792 | _EVAL_917;
  assign _EVAL_449 = ibuf__EVAL_22 | _EVAL_47;
  assign _EVAL_533 = _EVAL_167;
  assign _EVAL_759 = ~div__EVAL_0;
  assign _EVAL_265 = _EVAL_967 | _EVAL_503;
  assign _EVAL_577 = _EVAL_404 | _EVAL_294;
  assign _EVAL_173 = _EVAL_204 | _EVAL_986;
  assign _EVAL_142 = csr__EVAL_26;
  assign _EVAL_1108 = _EVAL_1409 & bpu__EVAL_25;
  assign _EVAL_261 = ibuf__EVAL_19[26];
  assign _EVAL_637 = _EVAL_525;
  assign _EVAL_1091 = _EVAL_1100;
  assign _EVAL_833 = _EVAL_1217 & _EVAL_259;
  assign _EVAL_867 = _EVAL_756 | _EVAL_448;
  assign _EVAL_930 = _EVAL_575 | _EVAL_1055;
  assign _EVAL_332 = _EVAL_1327 == 3'h0;
  assign bpu__EVAL_14 = csr__EVAL_109;
  assign _EVAL_205 = _EVAL_1379 & _EVAL_658;
  assign _EVAL_578 = _EVAL_703 == 5'h8;
  assign _EVAL_1115 = _EVAL_1165 | _EVAL_1289;
  assign _EVAL_422 = ibuf__EVAL_19 == 32'h73;
  assign _EVAL_618 = _EVAL_758;
  assign _EVAL_366 = _EVAL_362 | _EVAL_424;
  assign _EVAL_862 = _EVAL_1344 | _EVAL_514;
  assign _EVAL_529 = _EVAL_500 == 32'h0;
  assign _EVAL_481 = ibuf__EVAL_19 & 32'h20000020;
  assign _EVAL_368 = _EVAL_1083 & _EVAL_1393;
  assign _EVAL_821 = _EVAL_371 | _EVAL_1359;
  assign _EVAL_887 = _EVAL_1370 == 2'h1;
  assign _EVAL_720 = ~_EVAL_695;
  assign _EVAL_269 = ibuf__EVAL_19 & 32'h8;
  assign _EVAL_1195 = div__EVAL_0 | _EVAL_1263;
  assign _EVAL_830 = _EVAL_676 | _EVAL_1058;
  assign _EVAL_558 = _EVAL_1245 | _EVAL_796;
  assign _EVAL_58 = csr__EVAL_180;
  assign _EVAL_1209 = ~_EVAL_1117;
  assign _EVAL_1130 = _EVAL_1024 & _EVAL_1085;
  assign _EVAL_477 = ~_EVAL_15;
  assign csr__EVAL_113 = ibuf__EVAL_29[31:20];
  assign _EVAL_888 = _EVAL_946 == 32'h5013;
  assign _EVAL_280 = ibuf__EVAL_19[23:20];
  assign _EVAL_641 = ibuf__EVAL_19 & 32'h2002054;
  assign _EVAL_653 = |_EVAL_573;
  assign _EVAL_795 = _EVAL_665 | _EVAL_862;
  assign _EVAL_1242 = ~_EVAL_983;
  assign _EVAL_1035 = _EVAL_1155 | csr__EVAL_114;
  assign _EVAL_827 = _EVAL_574 | _EVAL_540;
  assign _EVAL_1006 = ibuf__EVAL_19 & 32'h4008;
  assign _EVAL_619 = _EVAL_1051 ? 4'hf : _EVAL_631;
  assign _EVAL_627 = _EVAL_629 | _EVAL_1040;
  assign _EVAL_1251 = _EVAL_559 | _EVAL_180;
  assign _EVAL_1022 = _EVAL_322 == 32'h4063;
  assign _EVAL_883 = _EVAL_1256 | _EVAL_200;
  assign _EVAL_292 = _EVAL_1340 != 3'h0;
  assign _EVAL_330 = _EVAL_1349 & _EVAL_1395;
  assign _EVAL_875 = ~csr__EVAL_155;
  assign _EVAL_1289 = ibuf__EVAL_19 == 32'h100073;
  assign _EVAL_398 = _EVAL_1327 == 3'h3;
  assign _EVAL_530 = _EVAL_974 | _EVAL_1156;
  assign _EVAL_646 = _EVAL_855 | _EVAL_359;
  assign _EVAL_245 = csr__EVAL_114 ? csr__EVAL_140 : {{28'd0}, _EVAL_842};
  assign _EVAL_513 = _EVAL_389 | _EVAL_247;
  assign _EVAL_954 = _EVAL_978 | _EVAL_1053;
  assign bpu__EVAL_43 = csr__EVAL_33;
  assign _EVAL_439 = _EVAL_612 == 32'h20;
  assign _EVAL_164 = _EVAL_477 | 32'h3;
  assign bpu__EVAL_33 = csr__EVAL_93;
  assign _EVAL_940 = _EVAL_1323 & csr__EVAL_77;
  assign csr__EVAL_134 = _EVAL_1335 & _EVAL_426;
  assign _EVAL_585 = _EVAL_283 | _EVAL_882;
  assign _EVAL_276 = _EVAL_1337 == 5'hd;
  assign bpu__EVAL_24 = csr__EVAL_74;
  assign _EVAL_1284 = _EVAL_335 & _EVAL_1273;
  assign _EVAL_848 = _EVAL_314 | _EVAL_356;
  assign _EVAL_275 = _EVAL_879 == 32'h202f;
  assign _EVAL_1028 = _EVAL_864[31:2];
  assign bpu__EVAL_32 = csr__EVAL_95;
  assign _EVAL_946 = ibuf__EVAL_19 & 32'hfe00707f;
  assign _EVAL_857 = _EVAL_441 == 32'h40000030;
  assign _EVAL_952 = _EVAL_428 ? _EVAL_1174 : _EVAL_520;
  assign _EVAL_54 = csr__EVAL_139;
  assign _EVAL_1030 = _EVAL_340 | _EVAL_557;
  assign _EVAL_28 = csr__EVAL_30;
  assign _EVAL_941 = _EVAL_946 == 32'h4033;
  assign _EVAL_518 = _EVAL_694[0];
  assign _EVAL_923 = ibuf__EVAL_19 & 32'h40004054;
  assign _EVAL_24 = _EVAL_821 | _EVAL_987;
  assign _EVAL_866 = _EVAL_347 & _EVAL_471;
  assign _EVAL_721 = 2'h1 == _EVAL_1386;
  assign _EVAL_41 = csr__EVAL_25;
  assign _EVAL_21 = csr__EVAL_172;
  assign _EVAL_1117 = _EVAL_843 | _EVAL_877;
  assign _EVAL_690 = _EVAL_1424[11:8];
  assign _EVAL_65 = _EVAL_1353;
  assign _EVAL_184 = _EVAL_879 == 32'h1800202f;
  assign _EVAL_231 = _EVAL_1358 == 2'h3;
  assign _EVAL_900 = _EVAL_322 == 32'h63;
  assign _EVAL_1249 = _EVAL_436 | _EVAL_1010;
  assign _EVAL_241 = _EVAL_1424[30:25];
  assign _EVAL_1312 = _EVAL_464;
  assign _EVAL_1096 = _EVAL_1005 == 32'h2002030;
  assign _EVAL_782 = _EVAL_846 | _EVAL_599;
  assign _EVAL_682 = ~_EVAL_1379;
  assign _EVAL_1081 = _EVAL_703 == 5'hd;
  assign _EVAL_479 = _EVAL_820 == 32'h6000;
  assign _EVAL_195 = _EVAL_1190 ? _EVAL_1347 : 32'h0;
  assign _EVAL_523 = _EVAL_1303 | _EVAL_947;
  assign _EVAL_1155 = _EVAL_517 | _EVAL_297;
  assign _EVAL_669 = _EVAL_841 == 32'hd;
  assign _EVAL_17 = csr__EVAL_98;
  assign _EVAL_232 = _EVAL_1302 & csr__EVAL_146;
  assign _EVAL_260 = _EVAL_1327 != 3'h2;
  assign _EVAL_95 = csr__EVAL_34;
  assign ibuf__EVAL_28 = _EVAL_71;
  assign _EVAL_501 = 2'h3 == _EVAL_1399;
  assign _EVAL_1280 = _EVAL_264;
  assign _EVAL_1222 = _EVAL_923 == 32'h4010;
  assign _EVAL_428 = _EVAL_1182 != 5'h0;
  assign _EVAL_1322 = _EVAL_1202 | _EVAL_1237;
  assign _EVAL_970 = _EVAL_1191 & _EVAL_838;
  assign _EVAL_904 = _EVAL_797 == _EVAL_181;
  assign _EVAL_443 = _EVAL_935 == 32'h0;
  assign _EVAL_244 = 32'h1 << _EVAL_729;
  assign _EVAL_1105 = _EVAL_627 & _EVAL_258;
  assign _EVAL_1093 = _EVAL_692 ? _EVAL_1377 : _EVAL_195;
  assign _EVAL_521 = ~_EVAL_539;
  assign _EVAL_813 = ibuf__EVAL_19 & 32'h2048;
  assign _EVAL_660 = _EVAL_260 & _EVAL_667;
  assign _EVAL_99 = csr__EVAL_2;
  assign _EVAL_951 = _EVAL_81 | _EVAL_1354;
  assign _EVAL_349 = _EVAL_958 | _EVAL_546;
  assign _EVAL_1075 = _EVAL_469 & _EVAL_406;
  assign _EVAL_556 = _EVAL_1420 & _EVAL_1244;
  assign _EVAL_1057 = _EVAL_1114 & ibuf__EVAL_22;
  assign _EVAL_807 = _EVAL_1143 | _EVAL_480;
  assign _EVAL_1295 = _EVAL_1251 | _EVAL_1290;
  assign _EVAL_899 = _EVAL_668 ? _EVAL_952 : _EVAL_520;
  assign _EVAL_704 = _EVAL_47 | _EVAL_1338;
  assign _EVAL_596 = _EVAL_1055 & _EVAL_1412;
  assign _EVAL_15 = _EVAL_766[31:0];
  assign _EVAL_1110 = _EVAL_906;
  assign _EVAL_340 = _EVAL_762 | _EVAL_1204;
  assign _EVAL_1098 = _EVAL_187 | _EVAL_207;
  assign _EVAL_1211 = _EVAL_322 == 32'h4003;
  assign _EVAL_1000 = ibuf__EVAL_19 & 32'h8000008;
  assign _EVAL_708 = ibuf__EVAL_19 & 32'h5054;
  assign _EVAL_599 = _EVAL_322 == 32'h5003;
  assign _EVAL_808 = _EVAL_878 | _EVAL_1062;
  assign _EVAL_1273 = ~_EVAL_1188;
  assign _EVAL_1278 = _EVAL_1415 ? _EVAL_1066 : _EVAL_998;
  assign _EVAL_974 = _EVAL_576 | _EVAL_919;
  assign _EVAL_459 = ibuf__EVAL_22 | ibuf__EVAL_5;
  assign _EVAL_503 = _EVAL_942 & _EVAL_754;
  assign _EVAL_314 = _EVAL_946 == 32'h2000033;
  assign _EVAL_411 = _EVAL_211 | _EVAL_273;
  assign _EVAL_146 = _EVAL_1325;
  assign _EVAL_61 = ~_EVAL_821;
  assign _EVAL_488 = _EVAL_698 == 32'h20;
  assign _EVAL_255 = _EVAL_942 & _EVAL_774;
  assign _EVAL_429 = _EVAL_966;
  assign _EVAL_335 = _EVAL_338 & _EVAL_539;
  assign _EVAL_734 = _EVAL_968 & _EVAL_1048;
  assign _EVAL_1002 = csr__EVAL_48 & _EVAL_875;
  assign _EVAL_919 = ibuf__EVAL_19 == 32'h70200073;
  assign _EVAL_1084 = csr__EVAL_108;
  assign _EVAL_550 = |_EVAL_831;
  assign _EVAL_676 = _EVAL_806 | _EVAL_1238;
  assign _EVAL_463 = _EVAL_1116 | _EVAL_1422;
  assign _EVAL_238 = ~_EVAL_645;
  assign bpu__EVAL_18 = csr__EVAL_92;
  assign _EVAL_1052 = ibuf__EVAL_27 ? 2'h1 : 2'h2;
  assign m__EVAL_1 = div__EVAL_4;
  assign _EVAL_172 = _EVAL_501 ? $signed(_EVAL_1149) : $signed(_EVAL_776);
  assign _EVAL_296 = _EVAL_987 & _EVAL_1188;
  assign _EVAL_746 = _EVAL_171 | _EVAL_876;
  assign _EVAL_586 = ibuf__EVAL_29[15:0];
  assign _EVAL_997 = _EVAL_1131 | _EVAL_893;
  assign _EVAL_1197 = _EVAL_1102 & _EVAL_775;
  assign _EVAL_497 = ~_EVAL_1239;
  assign _EVAL_825 = _EVAL_322 == 32'h5073;
  assign _EVAL_448 = _EVAL_20[2];
  assign _EVAL_748 = _EVAL_1337 == 5'h4;
  assign _EVAL_133 = csr__EVAL_144;
  assign _EVAL_490 = _EVAL_1366 | _EVAL_139;
  assign _EVAL_750 = _EVAL_310 == 32'h17;
  assign ibuf__EVAL_13 = ~_EVAL_297;
  assign _EVAL_289 = _EVAL_322 == 32'h2023;
  assign _EVAL_893 = _EVAL_946 == 32'h40005033;
  assign _EVAL_723 = {_EVAL_489,_EVAL_951,_EVAL_1359,_EVAL_1171,_EVAL_296,_EVAL_680,_EVAL_212,_EVAL_438,_EVAL_265,
    _EVAL_872};
  assign _EVAL_1038 = _EVAL_942 & _EVAL_904;
  assign _EVAL_222 = _EVAL_322 == 32'h6073;
  assign _EVAL_1269 = _EVAL_1137 | _EVAL_1361;
  assign _EVAL_836 = _EVAL_650 | _EVAL_1129;
  assign _EVAL_819 = _EVAL_453 | _EVAL_538;
  assign _EVAL_926 = _EVAL_946 == 32'h40000033;
  assign _EVAL_420 = _EVAL_1417[7];
  assign _EVAL_949 = ibuf__EVAL_19 & 32'h3044;
  assign _EVAL_1089 = {_EVAL_339,_EVAL_339};
  assign _EVAL_966 = _EVAL_1417[30:20];
  assign _EVAL_294 = _EVAL_269 == 32'h8;
  assign _EVAL_854 = ibuf__EVAL_19 & 32'h2050;
  assign _EVAL_1237 = ibuf__EVAL_19 == 32'h10500073;
  assign _EVAL_312 = _EVAL_332 ? _EVAL_420 : _EVAL_396;
  assign _EVAL_144 = ~_EVAL_892;
  assign bpu__EVAL_7 = csr__EVAL_162;
  assign _EVAL_885 = ibuf__EVAL_19 & 32'h2008;
  assign _EVAL_440 = _EVAL_585 | _EVAL_924;
  assign _EVAL_526 = _EVAL_1404[31:1];
  assign _EVAL_242 = _EVAL_976 | _EVAL_1077;
  assign _EVAL_628 = _EVAL_1197 & _EVAL_343;
  assign _EVAL_1109 = _EVAL_1367 | _EVAL_1422;
  assign _EVAL_736 = _EVAL_897 ? _EVAL_1332 : {{28'd0}, _EVAL_1264};
  assign _EVAL_209 = ibuf__EVAL_19 & 32'h2006054;
  assign _EVAL_352 = _EVAL_1370 == 2'h0;
  assign _EVAL_869 = _EVAL_1337 == 5'h8;
  assign _EVAL_787 = 2'h2 == _EVAL_1399;
  assign csr__EVAL_83 = _EVAL_74;
  assign _EVAL_1128 = _EVAL_1425 & bpu__EVAL_3;
  assign _EVAL_55 = csr__EVAL_119;
  assign _EVAL_1134 = _EVAL_624 & _EVAL_598;
  assign _EVAL_25 = csr__EVAL_163;
  assign _EVAL_214 = _EVAL_1002;
  assign _EVAL_1319 = ~csr__EVAL_115;
  assign _EVAL_385 = _EVAL_1379 & _EVAL_1373;
  assign _EVAL_1012 = _EVAL_1375 & _EVAL_1420;
  assign alu__EVAL_0 = _EVAL_1064;
  assign _EVAL_373 = div__EVAL_1;
  assign _EVAL_367 = 5'h0 == _EVAL_1261;
  assign _EVAL_145 = csr__EVAL_154;
  assign _EVAL_695 = _EVAL_411 | _EVAL_655;
  assign _EVAL_801 = _EVAL_547 == 32'h0;
  assign _EVAL_539 = _EVAL_319 | _EVAL_1367;
  assign _EVAL_1147 = _EVAL_955 | _EVAL_675;
  assign _EVAL_1171 = _EVAL_1284 & _EVAL_647;
  assign _EVAL_419 = _EVAL_770 | _EVAL_662;
  assign _EVAL_472 = _EVAL_417 | _EVAL_443;
  assign _EVAL_88 = csr__EVAL_131;
  assign _EVAL_433 = _EVAL_1295 | _EVAL_400;
  assign csr__EVAL_90 = _EVAL_147;
  assign _EVAL_937 = _EVAL_1424[20];
  assign _EVAL_20 = csr__EVAL_145;
  assign _EVAL_993 = {_EVAL_979,_EVAL_979,_EVAL_979,_EVAL_979};
  assign _EVAL_784 = _EVAL_1119 | ibuf__EVAL_23;
  assign _EVAL_108 = csr__EVAL_52;
  assign _EVAL_643 = _EVAL_1374 & _EVAL_891;
  assign _EVAL_288 = ~ibuf__EVAL_23;
  assign _EVAL_1136 = ~_EVAL_936;
  assign _EVAL_788 = _EVAL_664 | _EVAL_329;
  assign _EVAL_942 = _EVAL_194 & _EVAL_1221;
  assign _EVAL_217 = ~_EVAL_1035;
  assign _EVAL_616 = ibuf__EVAL_26 ? 4'hc : _EVAL_1016;
  assign _EVAL_789 = |_EVAL_1227;
  assign _EVAL_491 = _EVAL_700 == 32'h50;
  assign _EVAL_1292 = _EVAL_377;
  assign _EVAL_971 = _EVAL_322 == 32'h67;
  assign _EVAL_182 = _EVAL_516 | _EVAL_1416;
  assign _EVAL_194 = _EVAL_1178 | _EVAL_568;
  assign _EVAL_638 = _EVAL_841 == 32'h6;
  assign bpu__EVAL_35 = csr__EVAL_78;
  assign _EVAL_1305 = _EVAL_929 & _EVAL_863;
  assign _EVAL_1069 = _EVAL_419 | _EVAL_317;
  assign _EVAL_403 = _EVAL_705 | _EVAL_1307;
  assign _EVAL_998 = {_EVAL_1336,_EVAL_1413};
  assign _EVAL_213 = _EVAL_807 | _EVAL_401;
  assign _EVAL_913 = _EVAL_1116 ? $signed(_EVAL_786) : $signed(_EVAL_1218);
  assign _EVAL_1182 = _EVAL_627 ? _EVAL_729 : _EVAL_525;
  assign _EVAL_1301 = _EVAL_946 == 32'h2004033;
  assign _EVAL_34 = csr__EVAL_100;
  assign _EVAL_379 = _EVAL_703 == 5'h6;
  assign _EVAL_896 = _EVAL_930 | _EVAL_265;
  assign _EVAL_207 = _EVAL_1410 & _EVAL_759;
  assign _EVAL_914 = _EVAL_1358 == 2'h1;
  assign bpu__EVAL_13 = csr__EVAL_106;
  assign _EVAL_86 = csr__EVAL_2;
  assign _EVAL_889 = _EVAL_1357 & _EVAL_1394;
  assign _EVAL_370 = _EVAL_1008 & _EVAL_833;
  assign _EVAL_178 = _EVAL_717 & _EVAL_47;
  assign _EVAL_614 = _EVAL_1117 & _EVAL_1135;
  assign bpu__EVAL = csr__EVAL_46;
  assign _EVAL_663 = csr__EVAL_104[1:0];
  assign _EVAL_204 = _EVAL_1069 | _EVAL_638;
  assign _EVAL_1219 = _EVAL_1366 & _EVAL_747;
  assign _EVAL_765 = ibuf__EVAL_19 & 32'h4054;
  assign _EVAL_897 = _EVAL_1380 | _EVAL_1368;
  assign _EVAL_989 = _EVAL_310 == 32'h6f;
  assign _EVAL_431 = _EVAL_1375 & _EVAL_1257;
  assign _EVAL_1302 = _EVAL_624 & _EVAL_953;
  assign _EVAL_230 = _EVAL_1262 ? _EVAL_1377 : _EVAL_1101;
  assign _EVAL_829 = _EVAL_751 | _EVAL_1207;
  assign _EVAL_56 = _EVAL_552 & _EVAL_1319;
  assign _EVAL_365 = _EVAL_1323 | _EVAL_232;
  assign _EVAL_890 = _EVAL_369 & _EVAL_1152;
  assign _EVAL_336 = _EVAL_703 == 5'ha;
  assign csr__EVAL_130 = _EVAL_1401;
  assign _EVAL_994 = _EVAL_927 & _EVAL_23;
  assign _EVAL_1113 = _EVAL_946 == 32'h2007033;
  assign ibuf__EVAL_8 = _EVAL_105;
  assign _EVAL_916 = _EVAL_703 == 5'hc;
  assign _EVAL_357 = _EVAL_649 == 32'h8;
  assign _EVAL_1023 = _EVAL_946 == 32'h2002033;
  assign _EVAL_128 = _EVAL_1423;
  assign _EVAL_350 = _EVAL_1198;
  assign _EVAL_901 = ibuf__EVAL_7 ? 4'hc : {{2'd0}, _EVAL_1052};
  assign csr__EVAL_133 = _EVAL_44;
  assign _EVAL_447 = ibuf__EVAL_19 & 32'h1010;
  assign _EVAL_73 = csr__EVAL_17;
  assign _EVAL_924 = _EVAL_1337 == 5'h7;
  assign _EVAL_480 = _EVAL_879 == 32'h8000202f;
  assign _EVAL_800 = _EVAL_347 & _EVAL_433;
  assign _EVAL_395 = _EVAL_322 == 32'h1003;
  assign _EVAL_976 = _EVAL_465 | _EVAL_669;
  assign _EVAL_756 = _EVAL_933 | _EVAL_182;
  assign _EVAL_1320 = _EVAL_864[1:0];
  assign _EVAL_980 = _EVAL_1342 & _EVAL_601;
  assign _EVAL_680 = _EVAL_347 & _EVAL_1219;
  assign _EVAL_516 = _EVAL_1375 | _EVAL_1354;
  assign _EVAL_604 = _EVAL_1406 | _EVAL_1410;
  assign _EVAL_768 = _EVAL_879 == 32'h4000202f;
  assign _EVAL_132 = 1'h0;
  assign _EVAL_600 = _EVAL_420;
  assign _EVAL_1131 = _EVAL_822 | _EVAL_320;
  assign _EVAL_465 = _EVAL_564 | _EVAL_508;
  assign _EVAL_110 = _EVAL_1047 ? 2'h2 : _EVAL_824;
  assign _EVAL_396 = _EVAL_1139 ? _EVAL_215 : _EVAL_421;
  assign _EVAL_606 = _EVAL_252 | div__EVAL_3;
  assign _EVAL_677 = _EVAL_302;
  assign _EVAL_70 = csr__EVAL_24;
  assign _EVAL_762 = _EVAL_587 | _EVAL_680;
  assign _EVAL_583 = bpu__EVAL_2 ? 4'h3 : _EVAL_616;
  assign _EVAL_877 = _EVAL_927 & _EVAL_126;
  assign _EVAL_908 = _EVAL_721 ? $signed(_EVAL_533) : $signed(32'sh0);
  assign _EVAL_177 = _EVAL_1331;
  assign _EVAL_216 = _EVAL_459 ? _EVAL_1298 : 1'h1;
  assign _EVAL_442 = _EVAL_537 == 32'h2010;
  assign _EVAL_776 = _EVAL_787 ? $signed(_EVAL_1270) : $signed(32'sh0);
  assign _EVAL_657 = {{13'd0}, _EVAL_1288};
  assign _EVAL_301 = _EVAL_1337 == 5'h9;
  assign _EVAL_393 = _EVAL_946 == 32'h1013;
  assign _EVAL_835 = _EVAL_1060 | _EVAL_1074;
  assign _EVAL_935 = ibuf__EVAL_19 & 32'h30;
  assign _EVAL_1243 = _EVAL_1335 != 3'h0;
  assign bpu__EVAL_19 = csr__EVAL_14;
  assign _EVAL_504 = {_EVAL_472,_EVAL_577,_EVAL_1088};
  assign _EVAL_992 = _EVAL_566 | _EVAL_1145;
  assign _EVAL_274 = {_EVAL_1144,_EVAL_910,_EVAL_639,_EVAL_410,_EVAL_241,_EVAL_561,1'h0};
  assign _EVAL_228 = _EVAL_848 | _EVAL_509;
  assign _EVAL_10 = csr__EVAL_29;
  assign _EVAL_461 = _EVAL_445 | _EVAL_1004;
  assign _EVAL_1061 = _EVAL_703 == 5'hf;
  assign _EVAL_804 = _EVAL_1197 & _EVAL_1146;
  assign _EVAL_329 = _EVAL_322 == 32'h6063;
  assign _EVAL_1054 = csr__EVAL_115;
  assign csr__EVAL_120 = _EVAL_151;
  assign _EVAL_1315 = _EVAL_375 | _EVAL_865;
  assign _EVAL_1078 = ibuf__EVAL_19 & 32'h80000008;
  assign gated_clock_rocket_clock_gate_en = _EVAL_494 | _EVAL_178;
  assign _EVAL_519 = _EVAL_946 == 32'h1033;
  assign _EVAL_263 = _EVAL_1191 & _EVAL_1027;
  assign _EVAL_517 = _EVAL_282 | _EVAL_665;
  assign _EVAL_1146 = _EVAL_1261 == _EVAL_525;
  assign _EVAL_1202 = _EVAL_1115 | _EVAL_1168;
  assign _EVAL_304 = _EVAL_879 == 32'h6000202f;
  assign _EVAL_551 = _EVAL_1274 | _EVAL_511;
  assign _EVAL_5 = _EVAL_170 & _EVAL_582;
  assign _EVAL_582 = _EVAL_521 | _EVAL_727;
  assign _EVAL_324 = _EVAL_1375 ? 3'h0 : 3'h4;
  assign _EVAL_969 = ibuf__EVAL_19 & 32'h7044;
  assign _EVAL_894 = _EVAL_1304 ? _EVAL_1018 : _EVAL_372;
  assign _EVAL_655 = _EVAL_369 & _EVAL_1056;
  assign _EVAL_1167 = ~_EVAL_1357;
  assign _EVAL_780 = _EVAL_1370 < 2'h2;
  assign _EVAL_1193 = _EVAL_730 & _EVAL_1371;
  assign _EVAL_1270 = _EVAL_1278;
  assign _EVAL_884 = _EVAL_946 == 32'h3033;
  assign _EVAL_506 = _EVAL_946 == 32'h2005033;
  assign _EVAL_438 = _EVAL_1160 | _EVAL_536;
  assign _EVAL_405 = _EVAL_703 == 5'h14;
  assign _EVAL_1152 = _EVAL_181 == _EVAL_859;
  assign _EVAL_617 = _EVAL_635 | _EVAL_395;
  assign bpu__EVAL_39 = csr__EVAL_152;
  assign _EVAL_1198 = csr__EVAL_1;
  assign _EVAL_709 = ~_EVAL_1012;
  assign _EVAL_798 = _EVAL_605 & _EVAL_1067;
  assign _EVAL_256 = _EVAL_1186 | _EVAL_884;
  assign _EVAL_455 = _EVAL_545 ? $signed(_EVAL_600) : $signed(_EVAL_847);
  assign _EVAL_1079 = _EVAL_440 | _EVAL_538;
  assign _EVAL_414 = {_EVAL_621,_EVAL_1321};
  assign _EVAL_1255 = _EVAL_760 | _EVAL_1308;
  assign _EVAL_322 = ibuf__EVAL_19 & 32'h707f;
  assign _EVAL_672 = _EVAL_764 & _EVAL_840;
  assign _EVAL_210 = _EVAL_175 | _EVAL_480;
  assign _EVAL_166 = ibuf__EVAL_19 & 32'h34;
  assign _EVAL_732 = _EVAL_298 & _EVAL_261;
  assign _EVAL_1102 = _EVAL_1275 | _EVAL_327;
  assign _EVAL_1010 = _EVAL_1108 | _EVAL_1128;
  assign _EVAL_127 = _EVAL_955 | _EVAL_1249;
  assign _EVAL_1021 = _EVAL_755 == 3'h4;
  assign _EVAL_376 = _EVAL_851 == 32'h10000008;
  assign _EVAL_588 = _EVAL_288 & _EVAL_940;
  assign _EVAL_684 = _EVAL_439 | _EVAL_563;
  assign _EVAL_538 = _EVAL_193 | _EVAL_992;
  assign bpu__EVAL_10 = csr__EVAL_12;
  assign _EVAL_361 = ibuf__EVAL_19 & 32'h4058;
  assign _EVAL_912 = ~_EVAL_605;
  assign _EVAL_1261 = ibuf__EVAL_25;
  assign _EVAL_325 = 1'h0;
  assign _EVAL_741 = _EVAL_949 == 32'h3000;
  assign _EVAL_1043 = ibuf__EVAL_19 & 32'h44;
  assign _EVAL_793 = _EVAL_1309[31:2];
  assign _EVAL_364 = {{31'd0}, _EVAL_157};
  assign _EVAL_864 = _EVAL_668 ? _EVAL_266 : _EVAL_1071;
  assign _EVAL_743 = _EVAL_1402;
  assign _EVAL_837 = _EVAL_378 | _EVAL_763;
  assign _EVAL_278 = _EVAL_333 | _EVAL_971;
  assign _EVAL_917 = _EVAL_447 == 32'h1010;
  assign _EVAL_159 = csr__EVAL_8;
  assign _EVAL_318 = _EVAL_376 | _EVAL_1220;
  assign _EVAL_334 = {{30'd0}, _EVAL_950};
  assign _EVAL_49 = csr__EVAL_0;
  assign _EVAL_1037 = _EVAL_287 ? _EVAL_527 : _EVAL_216;
  assign _EVAL_211 = _EVAL_367 | _EVAL_661;
  assign _EVAL_1228 = ~ibuf__EVAL_22;
  assign _EVAL_623 = _EVAL_217 | csr__EVAL_114;
  assign _EVAL_693 = ~_EVAL_81;
  assign _EVAL_1042 = _EVAL_1215 | _EVAL_1038;
  assign _EVAL_920 = _EVAL_829 ? 6'h0 : _EVAL_873;
  assign ibuf__EVAL_1 = _EVAL_74;
  assign bpu__EVAL_34 = csr__EVAL_171;
  assign _EVAL_363 = _EVAL_398 ? $signed(_EVAL_1123) : $signed(_EVAL_455);
  assign _EVAL_620 = _EVAL_1379 | _EVAL_1351;
  assign _EVAL_174 = _EVAL_859 == _EVAL_168;
  assign _EVAL_430 = _EVAL_643 & _EVAL_292;
  assign _EVAL_552 = ibuf__EVAL_22 & _EVAL_347;
  assign _EVAL_642 = _EVAL_740 == 32'h1050;
  assign _EVAL_1020 = _EVAL_1024 & _EVAL_140;
  assign _EVAL_163 = 32'h1 << _EVAL_525;
  assign _EVAL_418 = _EVAL_405 | _EVAL_452;
  assign _EVAL_76 = {{1'd0}, _EVAL_957};
  assign _EVAL_1100 = {8{_EVAL_677}};
  assign _EVAL_645 = _EVAL_1011 | _EVAL_139;
  assign _EVAL_1310 = _EVAL_1337 == 5'he;
  assign _EVAL_354 = 2'h2 == _EVAL_1386;
  assign _EVAL_716 = _EVAL_1350[15:0];
  assign _EVAL_425 = _EVAL_902 == 32'h4;
  assign _EVAL_1063 = _EVAL_811 | _EVAL_771;
  assign _EVAL_1072 = 2'h1 == _EVAL_1399;
  assign bpu__EVAL_16 = csr__EVAL_186;
  assign _EVAL_1192 = _EVAL_627 ? _EVAL_244 : 32'h0;
  assign _EVAL_559 = _EVAL_475 | _EVAL_336;
  assign _EVAL_652 = _EVAL_221;
  assign _EVAL_343 = _EVAL_1261 == _EVAL_168;
  assign _EVAL_353 = _EVAL_1189 | _EVAL_109;
  assign _EVAL_1207 = _EVAL_1327 == 3'h5;
  assign _EVAL_94 = csr__EVAL_147;
  assign _EVAL_1238 = _EVAL_322 == 32'h23;
  assign _EVAL_102 = csr__EVAL_11;
  assign _EVAL_1034 = ibuf__EVAL_19 & 32'h1c;
  assign _EVAL_554 = _EVAL_899[31:2];
  assign _EVAL_1122 = _EVAL_1337 == 5'h11;
  assign _EVAL_408 = _EVAL_555[0];
  assign _EVAL_1203 = _EVAL_322 == 32'h7073;
  assign _EVAL_239 = _EVAL_386 == 2'h2;
  assign _EVAL_218 = _EVAL_1409 & bpu__EVAL_6;
  assign _EVAL_792 = _EVAL_883 | _EVAL_650;
  assign _EVAL_348 = _EVAL_1196;
  assign _EVAL_972 = _EVAL_663 == 2'h2;
  assign _EVAL_931 = _EVAL_515 | _EVAL_814;
  assign _EVAL_1229 = _EVAL_724 | _EVAL_1134;
  assign _EVAL_522 = ibuf__EVAL_19 & 32'h2004064;
  assign _EVAL_701 = _EVAL_1191 & _EVAL_1357;
  assign _EVAL_561 = _EVAL_1424[24:21];
  assign _EVAL_852 = _EVAL_1078 == 32'h80000008;
  assign _EVAL_851 = ibuf__EVAL_19 & 32'h10000008;
  assign _EVAL_1163 = _EVAL_354 ? $signed(_EVAL_959) : $signed(_EVAL_908);
  assign _EVAL_1204 = _EVAL_424 & _EVAL_606;
  assign _EVAL_630 = _EVAL_1300 & _EVAL_1357;
  assign _EVAL_180 = _EVAL_703 == 5'hb;
  assign _EVAL_1287 = {_EVAL_1315,_EVAL_697,_EVAL_785,_EVAL_1063};
  assign _EVAL_1121 = ibuf__EVAL_19 & 32'h40000008;
  assign _EVAL_382 = _EVAL_1362 | _EVAL_1397;
  assign _EVAL_237 = ibuf__EVAL_25 == 5'h0;
  assign _EVAL_689 = _EVAL_425 | _EVAL_650;
  assign _EVAL_880 = _EVAL_578 | _EVAL_916;
  assign _EVAL_1071 = _EVAL_1231__EVAL_1233_data;
  assign _EVAL_1307 = _EVAL_322 == 32'h3;
  assign _EVAL_826 = _EVAL_535;
  assign _EVAL_1074 = _EVAL_703 == 5'he;
  assign _EVAL_1142 = _EVAL_1087;
  assign _EVAL_574 = 5'h0 == _EVAL_859;
  assign csr__EVAL_50 = _EVAL_1416 ? _EVAL_1329 : {{28'd0}, _EVAL_262};
  assign _EVAL_794 = _EVAL_859 == _EVAL_181;
  assign _EVAL_933 = _EVAL_287 | _EVAL_726;
  assign _EVAL_96 = csr__EVAL_7;
  assign _EVAL_752 = _EVAL_1378 & _EVAL_347;
  assign _EVAL_745 = _EVAL_74;
  assign _EVAL_824 = _EVAL_850 ? 2'h3 : {{1'd0}, _EVAL_1109};
  assign _EVAL_1177 = _EVAL_226 | _EVAL_1096;
  assign alu__EVAL_3 = _EVAL_1376;
  assign _EVAL_400 = _EVAL_379 | _EVAL_220;
  assign csr__EVAL_20 = _EVAL_80;
  assign _EVAL_527 = _EVAL_713 != _EVAL_1356;
  assign _EVAL_1300 = _EVAL_1379 & _EVAL_764;
  assign _EVAL_64 = csr__EVAL_43;
  assign _EVAL_1103 = _EVAL_529 | _EVAL_763;
  assign _EVAL_546 = _EVAL_798 ? _EVAL_163 : 32'h0;
  assign _EVAL_1009 = _EVAL_714 | ibuf__EVAL_7;
  assign _EVAL_543 = _EVAL_663 == 2'h1;
  assign _EVAL_1104 = _EVAL_366 & _EVAL_874;
  assign csr__EVAL_141 = _EVAL_103;
  assign _EVAL_589 = _EVAL_1337 == 5'h1;
  assign _EVAL_557 = ~_EVAL_922;
  assign _EVAL_153 = 4'h0;
  assign _EVAL_515 = _EVAL_1175 | _EVAL_1094;
  assign _EVAL_722 = _EVAL_707 | _EVAL_1166;
  assign _EVAL_536 = _EVAL_1055 & _EVAL_1243;
  assign _EVAL_1047 = _EVAL_1109 & _EVAL_853;
  assign gated_clock_rocket_clock_gate_in = _EVAL_92;
  assign _EVAL_189 = _EVAL_836 | _EVAL_347;
  assign _EVAL_272 = ~_EVAL_699;
  assign _EVAL_77 = csr__EVAL_47;
  assign csr__EVAL_166 = _EVAL_1392;
  assign _EVAL_1215 = _EVAL_581 | _EVAL_197;
  assign _EVAL_1276 = _EVAL_841 == 32'h7;
  assign _EVAL_235 = _EVAL_623 | ibuf__EVAL_4;
  assign _EVAL_737 = ibuf__EVAL_19 & 32'hc;
  assign _EVAL_1208 = _EVAL_1247 == 32'h1008;
  assign ibuf__EVAL_5 = _EVAL_47;
  assign _EVAL_822 = _EVAL_625 | _EVAL_519;
  assign _EVAL_505 = _EVAL_962 | _EVAL_778;
  assign _EVAL_724 = _EVAL_683 | _EVAL_496;
  assign _EVAL_670 = ibuf__EVAL_19 == 32'h30500073;
  assign _EVAL_484 = _EVAL_953 & csr__EVAL_37;
  assign bpu__EVAL_17 = csr__EVAL_157;
  assign _EVAL_402 = _EVAL_845 | _EVAL_900;
  assign div__EVAL_6 = _EVAL_1333 ? _EVAL_963 : _EVAL_1230;
  assign _EVAL_266 = _EVAL_428 ? _EVAL_485 : _EVAL_1071;
  assign _EVAL_1032 = _EVAL_427;
  assign _EVAL_777 = 5'h1 == _EVAL_1164;
  assign div__EVAL_10 = _EVAL_629 ? 1'h0 : _EVAL_709;
  assign _EVAL_285 = ibuf__EVAL_19 & 32'h70;
  assign _EVAL_215 = _EVAL_1417[20];
  assign _EVAL_138 = csr__EVAL_40;
  assign _EVAL_1070 = _EVAL_951 | _EVAL_1117;
  assign _EVAL_525 = _EVAL_1364[11:7];
  assign _EVAL_964 = _EVAL_942 & _EVAL_749;
  assign csr__EVAL_126 = _EVAL_131;
  assign csr__EVAL_85 = gated_clock_rocket_clock_gate_out;
  assign _EVAL_754 = _EVAL_408 & _EVAL_1136;
  assign _EVAL_427 = _EVAL_751 ? $signed(_EVAL_429) : $signed({11{_EVAL_847}});
  assign _EVAL_50 = csr__EVAL_137;
  assign _EVAL_471 = _EVAL_703 == 5'h1;
  assign _EVAL_1258 = _EVAL_609 | _EVAL_479;
  assign _EVAL_918 = _EVAL_1182 == _EVAL_859;
  assign _EVAL_19 = csr__EVAL_164 & _EVAL_272;
  assign _EVAL_595 = _EVAL_322 == 32'h2003;
  assign _EVAL_165 = _EVAL_469[0];
  assign _EVAL_1184 = _EVAL_844 == 32'h40001010;
  assign _EVAL_733 = _EVAL_924 | _EVAL_780;
  assign _EVAL_148 = _EVAL_112;
  assign _EVAL_1263 = div__EVAL_11 & _EVAL_709;
  assign _EVAL_291 = _EVAL_711 == 32'h1010;
  assign _EVAL_770 = _EVAL_841 == 32'h2;
  assign _EVAL_13 = csr__EVAL_65;
  assign csr__EVAL_5 = _EVAL_82;
  assign _EVAL_1133 = _EVAL_310 == 32'h37;
  assign div__EVAL_5 = _EVAL_74;
  assign _EVAL_391 = _EVAL_1374 | _EVAL_1379;
  assign _EVAL_1286 = _EVAL_643 & _EVAL_1395;
  assign _EVAL_1248 = _EVAL_432 | _EVAL_651;
  assign csr__EVAL_41 = _EVAL_92;
  assign _EVAL_909 = {_EVAL_1144,_EVAL_910,_EVAL_1091,_EVAL_313,_EVAL_241,_EVAL_690,1'h0};
  assign csr__EVAL_86 = _EVAL_1390;
  assign _EVAL_328 = _EVAL_323 | _EVAL_276;
  assign _EVAL_406 = {{18'd0}, _EVAL_965};
  assign _EVAL_841 = _EVAL_1416 ? _EVAL_1329 : {{28'd0}, _EVAL_262};
  assign _EVAL_626 = _EVAL_1140 >> _EVAL_859;
  assign _EVAL_858 = _EVAL_755 == 3'h7;
  assign _EVAL_1281 = _EVAL_168 == _EVAL_859;
  assign m__EVAL_0 = div__EVAL_6;
  assign _EVAL_1161 = _EVAL_703 == 5'h9;
  assign _EVAL_219 = _EVAL_322 == 32'h5063;
  assign _EVAL_454 = _EVAL_1374 & _EVAL_1342;
  assign _EVAL_1185 = _EVAL_981 | _EVAL_821;
  assign _EVAL_840 = _EVAL_1269 | _EVAL_1421;
  assign _EVAL_14 = csr__EVAL_185;
  assign _EVAL_872 = _EVAL_562 | _EVAL_470;
  assign _EVAL_1257 = ~_EVAL_951;
  assign _EVAL_1213 = _EVAL_828 == 32'h0;
  assign _EVAL_134 = csr__EVAL_80;
  assign _EVAL_1090 = _EVAL_627 ? _EVAL_373 : _EVAL_1200;
  assign _EVAL_706 = _EVAL_391 | _EVAL_1375;
  assign _EVAL_1092 = |_EVAL_444;
  assign _EVAL_121 = _EVAL_319 | _EVAL_1367;
  assign _EVAL_612 = ibuf__EVAL_19 & 32'h28;
  assign csr__EVAL_21 = _EVAL_53;
  assign _EVAL_1014 = _EVAL_347 & _EVAL_985;
  assign _EVAL_1186 = _EVAL_1026 | _EVAL_512;
  assign _EVAL_978 = _EVAL_748 | _EVAL_301;
  assign _EVAL_79 = _EVAL_911 & _EVAL_693;
  assign _EVAL_1236 = _EVAL_275 | _EVAL_1094;
  assign _EVAL_186 = ~_EVAL_290;
  assign m__EVAL_5 = div__EVAL_9;
  assign _EVAL_640 = _EVAL_722 | _EVAL_650;
  assign _EVAL_580 = _EVAL_1241 | _EVAL_184;
  assign _EVAL_747 = ~_EVAL_32;
  assign ibuf__EVAL_3 = gated_clock_rocket_clock_gate_out;
  assign _EVAL_323 = _EVAL_869 | _EVAL_253;
  assign _EVAL_1114 = ~_EVAL_665;
  assign _EVAL_1159 = _EVAL_1248 | _EVAL_791;
  assign _EVAL_40 = 1'h0;
  assign _EVAL_221 = _EVAL_1424[7];
  assign _EVAL_297 = _EVAL_409 | _EVAL_473;
  assign _EVAL_327 = _EVAL_854 == 32'h2000;
  assign _EVAL_1321 = _EVAL_640 | _EVAL_344;
  assign _EVAL_1143 = _EVAL_534 | _EVAL_768;
  assign _EVAL_696 = ~_EVAL_415;
  assign m__EVAL_2 = _EVAL_1374 & _EVAL_1406;
  assign _EVAL_375 = _EVAL_1159 | _EVAL_857;
  assign _EVAL_233 = _EVAL_1285 | _EVAL_277;
  assign _EVAL_995 = _EVAL_322 == 32'h6013;
  assign _EVAL_785 = _EVAL_1212 | _EVAL_1184;
  assign _EVAL_1205 = _EVAL_291 | _EVAL_710;
  assign _EVAL_270 = _EVAL_532 | _EVAL_1208;
  assign _EVAL_1191 = _EVAL_1379 & _EVAL_672;
  assign ibuf__EVAL_16 = _EVAL_48;
  assign _EVAL_1166 = _EVAL_737 == 32'h4;
  assign _EVAL_1170 = _EVAL_481 == 32'h20000020;
  assign _EVAL_1200 = _EVAL_1243 ? csr__EVAL_103 : _EVAL_999;
  assign _EVAL_1066 = _EVAL_284 ? _EVAL_152 : _EVAL_1093;
  assign _EVAL_838 = _EVAL_1361 | _EVAL_1421;
  assign _EVAL_421 = _EVAL_1207 & _EVAL_1036;
  assign _EVAL_834 = _EVAL_684 | _EVAL_1170;
  assign _EVAL_181 = _EVAL_1424[11:7];
  assign _EVAL_602 = csr__EVAL_1[4:0];
  assign _EVAL_648 = _EVAL_1236 | _EVAL_814;
  assign _EVAL_66 = csr__EVAL_15;
  assign _EVAL_512 = _EVAL_946 == 32'h2033;
  assign _EVAL_542 = _EVAL_355 == 32'h6000;
  assign _EVAL_1227 = _EVAL_469 & _EVAL_1048;
  assign _EVAL_844 = ibuf__EVAL_19 & 32'h40001054;
  assign _EVAL_1260 = _EVAL_1425 & bpu__EVAL_28;
  assign _EVAL_675 = _EVAL_1073 | _EVAL_735;
  assign _EVAL_547 = ibuf__EVAL_19 & 32'h48;
  assign _EVAL_944 = _EVAL_274;
  assign _EVAL_664 = _EVAL_402 | _EVAL_1022;
  assign _EVAL_311 = _EVAL_641 == 32'h2010;
  assign _EVAL_786 = _EVAL_909;
  assign _EVAL_562 = _EVAL_1286 | _EVAL_701;
  assign _EVAL_579 = _EVAL_473 & _EVAL_497;
  assign _EVAL_441 = ibuf__EVAL_19 & 32'h40003034;
  assign _EVAL_143 = csr__EVAL_173;
  assign _EVAL_928 = ibuf__EVAL_19 & 32'h54;
  assign _EVAL_806 = _EVAL_457 | _EVAL_599;
  assign _EVAL_331 = _EVAL_1364[31:16];
  always @(posedge _EVAL_92) begin
    _EVAL_337 <= _EVAL_1054 | _EVAL_579;
    if (_EVAL_1239) begin
      _EVAL_473 <= 1'h0;
    end else if (_EVAL_217) begin
      _EVAL_473 <= _EVAL_613;
    end
    _EVAL_634 <= _EVAL_933 | _EVAL_498;
    _EVAL_699 <= _EVAL_74 | _EVAL_553;
  end
  always @(posedge gated_clock_rocket_clock_gate_out) begin
    if(_EVAL_1231__EVAL_1234_en & _EVAL_1231__EVAL_1234_mask) begin
      _EVAL_1231[_EVAL_1231__EVAL_1234_addr] <= _EVAL_1231__EVAL_1234_data;
    end
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        if (_EVAL_330) begin
          if (_EVAL_352) begin
            _EVAL_1325 <= _EVAL_993;
          end else begin
            _EVAL_1325 <= _EVAL_597;
          end
        end
      end
    end
    if (_EVAL_217) begin
      _EVAL_1326 <= _EVAL_394;
    end
    if (_EVAL_217) begin
      _EVAL_1327 <= _EVAL_504;
    end
    if (_EVAL_235) begin
      _EVAL_1328 <= ibuf__EVAL_12;
    end
    if (_EVAL_726) begin
      if (_EVAL_897) begin
        _EVAL_1329 <= _EVAL_1332;
      end else begin
        _EVAL_1329 <= {{28'd0}, _EVAL_1264};
      end
    end
    if (_EVAL_726) begin
      _EVAL_1330 <= _EVAL_1346;
    end
    _EVAL_1331 <= _EVAL_1414;
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        _EVAL_1332 <= _EVAL_1398;
      end
    end
    if (_EVAL_217) begin
      if (_EVAL_796) begin
        _EVAL_1333 <= 1'h0;
      end else begin
        _EVAL_1333 <= _EVAL_695;
      end
    end
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        _EVAL_1334 <= _EVAL_1405;
      end
    end
    if (_EVAL_726) begin
      _EVAL_1335 <= _EVAL_1403;
    end
    if (_EVAL_217) begin
      if (_EVAL_818) begin
        _EVAL_1336 <= _EVAL_1028;
      end
    end
    if (_EVAL_217) begin
      _EVAL_1337 <= _EVAL_703;
    end
    _EVAL_1338 <= _EVAL_47;
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        _EVAL_1339 <= alu__EVAL_1;
      end
    end
    if (_EVAL_217) begin
      if (_EVAL_945) begin
        _EVAL_1340 <= 3'h2;
      end else begin
        _EVAL_1340 <= _EVAL_755;
      end
    end
    if (_EVAL_287) begin
      _EVAL_1341 <= _EVAL_1372;
    end
    if (_EVAL_217) begin
      _EVAL_1342 <= _EVAL_194;
    end
    if (_EVAL_217) begin
      _EVAL_1343 <= _EVAL_550;
    end
    _EVAL_1344 <= _EVAL_1057 & ibuf__EVAL_4;
    _EVAL_1345 <= _EVAL_1418;
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        _EVAL_1346 <= _EVAL_603;
      end
    end
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        _EVAL_1347 <= _EVAL_201;
      end
    end
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        _EVAL_1348 <= _EVAL_1342;
      end
    end
    if (_EVAL_217) begin
      _EVAL_1349 <= _EVAL_1138;
    end
    if (_EVAL_726) begin
      _EVAL_1350 <= _EVAL_1419;
    end
    _EVAL_1351 <= _EVAL_1114 & _EVAL_862;
    if (_EVAL_217) begin
      _EVAL_1352 <= _EVAL_650;
    end
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        _EVAL_1353 <= _EVAL_1383;
      end
    end
    _EVAL_1354 <= _EVAL_502 & _EVAL_658;
    if (_EVAL_726) begin
      _EVAL_1355 <= _EVAL_1341;
    end
    if (_EVAL_235) begin
      _EVAL_1356 <= ibuf__EVAL_15;
    end
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        _EVAL_1357 <= _EVAL_1395;
      end
    end
    if (_EVAL_217) begin
      if (_EVAL_796) begin
        _EVAL_1358 <= _EVAL_772;
      end else if (_EVAL_1001) begin
        _EVAL_1358 <= _EVAL_1127;
      end else if (_EVAL_367) begin
        _EVAL_1358 <= 2'h0;
      end else begin
        _EVAL_1358 <= _EVAL_1240;
      end
    end
    _EVAL_1359 <= _EVAL_381 & _EVAL_1373;
    if (_EVAL_235) begin
      _EVAL_1360 <= ibuf__EVAL_29;
    end
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        _EVAL_1361 <= _EVAL_1406;
      end
    end
    _EVAL_1362 <= _EVAL_1057 & csr__EVAL_114;
    if (_EVAL_217) begin
      _EVAL_1363 <= _EVAL_1208;
    end
    if (_EVAL_726) begin
      _EVAL_1364 <= _EVAL_1424;
    end
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        _EVAL_1365 <= _EVAL_1384;
      end
    end
    _EVAL_1366 <= _EVAL_234 & _EVAL_1268;
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        _EVAL_1367 <= _EVAL_1352;
      end
    end
    _EVAL_1368 <= _EVAL_696 & _EVAL_382;
    if (_EVAL_287) begin
      _EVAL_1369 <= _EVAL_1343;
    end
    if (_EVAL_217) begin
      if (_EVAL_418) begin
        _EVAL_1370 <= _EVAL_790;
      end else begin
        _EVAL_1370 <= _EVAL_644;
      end
    end
    if (_EVAL_726) begin
      _EVAL_1371 <= _EVAL_1369;
    end
    if (_EVAL_217) begin
      _EVAL_1372 <= _EVAL_199;
    end
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        _EVAL_1373 <= _EVAL_1314;
      end
    end
    _EVAL_1374 <= ~_EVAL_1035;
    _EVAL_1375 <= ~_EVAL_1147;
    if (_EVAL_217) begin
      if (_EVAL_558) begin
        _EVAL_1376 <= 4'h0;
      end else begin
        _EVAL_1376 <= _EVAL_1287;
      end
    end
    if (_EVAL_726) begin
      _EVAL_1377 <= _EVAL_435;
    end
    if (_EVAL_74) begin
      _EVAL_1378 <= 1'h0;
    end else if (_EVAL_217) begin
      _EVAL_1378 <= _EVAL_203;
    end else if (_EVAL_238) begin
      _EVAL_1378 <= 1'h0;
    end
    _EVAL_1379 <= ~_EVAL_415;
    _EVAL_1380 <= _EVAL_1114 & _EVAL_1362;
    if (_EVAL_726) begin
      _EVAL_1381 <= _EVAL_1361;
    end
    if (_EVAL_217) begin
      _EVAL_1383 <= _EVAL_666;
    end
    if (_EVAL_235) begin
      _EVAL_1384 <= ibuf__EVAL_9;
    end
    if (_EVAL_217) begin
      if (_EVAL_558) begin
        if (_EVAL_1224) begin
          _EVAL_1386 <= 2'h2;
        end else if (_EVAL_1119) begin
          _EVAL_1386 <= 2'h2;
        end else begin
          _EVAL_1386 <= 2'h1;
        end
      end else begin
        _EVAL_1386 <= _EVAL_499;
      end
    end
    if (_EVAL_217) begin
      _EVAL_1387 <= _EVAL_1129;
    end
    if (_EVAL_217) begin
      if (_EVAL_558) begin
        _EVAL_1388 <= _EVAL_784;
      end else begin
        _EVAL_1388 <= ibuf__EVAL_23;
      end
    end
    if (_EVAL_973) begin
      _EVAL_1390 <= _EVAL_653;
    end else if (_EVAL_972) begin
      _EVAL_1390 <= _EVAL_653;
    end else if (_EVAL_543) begin
      _EVAL_1390 <= _EVAL_437;
    end else if (_EVAL_1117) begin
      _EVAL_1390 <= _EVAL_467;
    end else begin
      _EVAL_1390 <= _EVAL_1193;
    end
    if (_EVAL_726) begin
      _EVAL_1391 <= _EVAL_1357;
    end
    if (_EVAL_482) begin
      _EVAL_1392 <= _EVAL_1059;
    end else if (_EVAL_239) begin
      _EVAL_1392 <= _EVAL_1059;
    end else if (_EVAL_1272) begin
      _EVAL_1392 <= _EVAL_789;
    end else if (_EVAL_1117) begin
      _EVAL_1392 <= _EVAL_165;
    end else begin
      _EVAL_1392 <= _EVAL_341;
    end
    if (_EVAL_217) begin
      _EVAL_1393 <= _EVAL_630;
    end
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        _EVAL_1394 <= _EVAL_733;
      end
    end
    if (_EVAL_217) begin
      _EVAL_1395 <= _EVAL_347;
    end
    _EVAL_1397 <= _EVAL_217 & _EVAL_558;
    if (_EVAL_235) begin
      if (csr__EVAL_114) begin
        _EVAL_1398 <= csr__EVAL_140;
      end else begin
        _EVAL_1398 <= {{28'd0}, _EVAL_842};
      end
    end
    if (_EVAL_217) begin
      if (_EVAL_558) begin
        if (_EVAL_1224) begin
          _EVAL_1399 <= 2'h0;
        end else if (_EVAL_1119) begin
          _EVAL_1399 <= 2'h1;
        end else begin
          _EVAL_1399 <= 2'h0;
        end
      end else begin
        _EVAL_1399 <= _EVAL_414;
      end
    end
    if (_EVAL_217) begin
      if (_EVAL_796) begin
        _EVAL_1400 <= _EVAL_793;
      end else if (_EVAL_1001) begin
        _EVAL_1400 <= _EVAL_554;
      end
    end
    if (_EVAL_726) begin
      _EVAL_1401 <= _EVAL_1402;
    end
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        _EVAL_1402 <= _EVAL_1356;
      end
    end
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        _EVAL_1403 <= _EVAL_1340;
      end
    end
    if (_EVAL_74) begin
      _EVAL_1404 <= 32'h0;
    end else if (_EVAL_299) begin
      _EVAL_1404 <= _EVAL_349;
    end else if (_EVAL_627) begin
      _EVAL_1404 <= _EVAL_958;
    end
    if (_EVAL_235) begin
      _EVAL_1405 <= ibuf__EVAL_20;
    end
    if (_EVAL_217) begin
      _EVAL_1406 <= _EVAL_362;
    end
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        _EVAL_1407 <= _EVAL_1388;
      end
    end
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        _EVAL_1409 <= _EVAL_812;
      end
    end
    if (_EVAL_217) begin
      _EVAL_1410 <= _EVAL_424;
    end
    _EVAL_1411 <= div__EVAL_0 & div__EVAL_3;
    if (_EVAL_726) begin
      _EVAL_1412 <= _EVAL_1421;
    end
    if (_EVAL_217) begin
      if (_EVAL_818) begin
        _EVAL_1413 <= _EVAL_1320;
      end else if (_EVAL_574) begin
        _EVAL_1413 <= 2'h0;
      end else if (_EVAL_540) begin
        _EVAL_1413 <= 2'h1;
      end else begin
        _EVAL_1413 <= _EVAL_450;
      end
    end
    if (_EVAL_1333) begin
      if (_EVAL_231) begin
        _EVAL_1414 <= _EVAL_152;
      end else if (_EVAL_1262) begin
        _EVAL_1414 <= _EVAL_1377;
      end else if (_EVAL_914) begin
        _EVAL_1414 <= _EVAL_1347;
      end else begin
        _EVAL_1414 <= 32'h0;
      end
    end else begin
      _EVAL_1414 <= _EVAL_1230;
    end
    if (_EVAL_217) begin
      _EVAL_1415 <= _EVAL_983;
    end
    _EVAL_1416 <= _EVAL_675 & _EVAL_658;
    if (_EVAL_235) begin
      _EVAL_1417 <= ibuf__EVAL_19;
    end
    if (_EVAL_1415) begin
      if (_EVAL_284) begin
        _EVAL_1418 <= _EVAL_152;
      end else if (_EVAL_692) begin
        _EVAL_1418 <= _EVAL_1377;
      end else if (_EVAL_1190) begin
        _EVAL_1418 <= _EVAL_1347;
      end else begin
        _EVAL_1418 <= 32'h0;
      end
    end else begin
      _EVAL_1418 <= _EVAL_998;
    end
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        _EVAL_1419 <= _EVAL_1360;
      end
    end
    if (_EVAL_726) begin
      _EVAL_1420 <= _EVAL_1348;
    end
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        _EVAL_1421 <= _EVAL_1410;
      end
    end
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        _EVAL_1422 <= _EVAL_1387;
      end
    end
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        _EVAL_1423 <= _EVAL_1328;
      end
    end
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        _EVAL_1424 <= _EVAL_1417;
      end
    end
    if (!(_EVAL_385)) begin
      if (_EVAL_287) begin
        _EVAL_1425 <= _EVAL_1076;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_5 = {1{`RANDOM}};
  _RAND_6 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 31; initvar = initvar+1)
    _EVAL_1231[initvar] = _RAND_4[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_337 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_473 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_634 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_699 = _RAND_3[0:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_1325 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_1326 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_1327 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_1328 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_1329 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_1330 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_1331 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_1332 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_1333 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_1334 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _EVAL_1335 = _RAND_17[2:0];
  _RAND_18 = {1{`RANDOM}};
  _EVAL_1336 = _RAND_18[29:0];
  _RAND_19 = {1{`RANDOM}};
  _EVAL_1337 = _RAND_19[4:0];
  _RAND_20 = {1{`RANDOM}};
  _EVAL_1338 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _EVAL_1339 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  _EVAL_1340 = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  _EVAL_1341 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  _EVAL_1342 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  _EVAL_1343 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  _EVAL_1344 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  _EVAL_1345 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  _EVAL_1346 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  _EVAL_1347 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  _EVAL_1348 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  _EVAL_1349 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  _EVAL_1350 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  _EVAL_1351 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  _EVAL_1352 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  _EVAL_1353 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  _EVAL_1354 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  _EVAL_1355 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  _EVAL_1356 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  _EVAL_1357 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  _EVAL_1358 = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  _EVAL_1359 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  _EVAL_1360 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  _EVAL_1361 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  _EVAL_1362 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  _EVAL_1363 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  _EVAL_1364 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  _EVAL_1365 = _RAND_47[4:0];
  _RAND_48 = {1{`RANDOM}};
  _EVAL_1366 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  _EVAL_1367 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  _EVAL_1368 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  _EVAL_1369 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  _EVAL_1370 = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  _EVAL_1371 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  _EVAL_1372 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  _EVAL_1373 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  _EVAL_1374 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  _EVAL_1375 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  _EVAL_1376 = _RAND_58[3:0];
  _RAND_59 = {1{`RANDOM}};
  _EVAL_1377 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  _EVAL_1378 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  _EVAL_1379 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  _EVAL_1380 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  _EVAL_1381 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  _EVAL_1383 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  _EVAL_1384 = _RAND_65[4:0];
  _RAND_66 = {1{`RANDOM}};
  _EVAL_1386 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  _EVAL_1387 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  _EVAL_1388 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  _EVAL_1390 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  _EVAL_1391 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  _EVAL_1392 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  _EVAL_1393 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  _EVAL_1394 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  _EVAL_1395 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  _EVAL_1397 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  _EVAL_1398 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  _EVAL_1399 = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  _EVAL_1400 = _RAND_78[29:0];
  _RAND_79 = {1{`RANDOM}};
  _EVAL_1401 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  _EVAL_1402 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  _EVAL_1403 = _RAND_81[2:0];
  _RAND_82 = {1{`RANDOM}};
  _EVAL_1404 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  _EVAL_1405 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  _EVAL_1406 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  _EVAL_1407 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  _EVAL_1409 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  _EVAL_1410 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  _EVAL_1411 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  _EVAL_1412 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  _EVAL_1413 = _RAND_90[1:0];
  _RAND_91 = {1{`RANDOM}};
  _EVAL_1414 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  _EVAL_1415 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  _EVAL_1416 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  _EVAL_1417 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  _EVAL_1418 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  _EVAL_1419 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  _EVAL_1420 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  _EVAL_1421 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  _EVAL_1422 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  _EVAL_1423 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  _EVAL_1424 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  _EVAL_1425 = _RAND_102[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
