//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module SiFive_CoreIPSubsystem(
  input          clock,
  input          reset,
  input          external_source_for_core_0_clock,
  input          external_source_for_core_0_reset,
  output         halt_from_tile_0,
  output         wfi_from_tile_0,
  output         cease_from_tile_0,
  output         debug_from_tile_0,
  input          psd_test_clock_enable,
  input          resetctrl_hartIsInReset_0,
  input          debug_clock,
  input          debug_reset,
  input          debug_systemjtag_jtag_TCK,
  input          debug_systemjtag_jtag_TMS,
  input          debug_systemjtag_jtag_TDI,
  output         debug_systemjtag_jtag_TDO_data,
  output         debug_systemjtag_jtag_TDO_driven,
  input          debug_systemjtag_reset,
  input  [10:0]  debug_systemjtag_mfr_id,
  input  [15:0]  debug_systemjtag_part_number,
  input  [3:0]   debug_systemjtag_version,
  output         debug_ndreset,
  output         debug_dmactive,
  input          debug_dmactiveAck,
  input  [31:0]  reset_vector_0,
  input          nmi_0_rnmi,
  input  [31:0]  nmi_0_rnmi_interrupt_vector,
  input  [31:0]  nmi_0_rnmi_exception_vector,
  input          rtc_toggle,
  input  [126:0] global_interrupts,
  input  [15:0]  local_interrupts_0,
  output         sys_port_ahb_0_hmastlock,
  input          sys_port_ahb_0_hready,
  output [1:0]   sys_port_ahb_0_htrans,
  output [2:0]   sys_port_ahb_0_hsize,
  output [2:0]   sys_port_ahb_0_hburst,
  output         sys_port_ahb_0_hwrite,
  output [3:0]   sys_port_ahb_0_hprot,
  output [30:0]  sys_port_ahb_0_haddr,
  output [31:0]  sys_port_ahb_0_hwdata,
  input          sys_port_ahb_0_hresp,
  input  [31:0]  sys_port_ahb_0_hrdata,
  output         periph_port_ahb_0_hmastlock,
  input          periph_port_ahb_0_hready,
  output [1:0]   periph_port_ahb_0_htrans,
  output [2:0]   periph_port_ahb_0_hsize,
  output [2:0]   periph_port_ahb_0_hburst,
  output         periph_port_ahb_0_hwrite,
  output [3:0]   periph_port_ahb_0_hprot,
  output [29:0]  periph_port_ahb_0_haddr,
  output [31:0]  periph_port_ahb_0_hwdata,
  input          periph_port_ahb_0_hresp,
  input  [31:0]  periph_port_ahb_0_hrdata,
  input          front_port_ahb_0_hmastlock,
  input          front_port_ahb_0_hsel,
  input          front_port_ahb_0_hready,
  output         front_port_ahb_0_hreadyout,
  input  [1:0]   front_port_ahb_0_htrans,
  input  [2:0]   front_port_ahb_0_hsize,
  input  [2:0]   front_port_ahb_0_hburst,
  input          front_port_ahb_0_hwrite,
  input  [3:0]   front_port_ahb_0_hprot,
  input  [31:0]  front_port_ahb_0_haddr,
  input  [31:0]  front_port_ahb_0_hwdata,
  output         front_port_ahb_0_hresp,
  output [31:0]  front_port_ahb_0_hrdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL;
  wire  _EVAL_0;
  wire  _EVAL_1;
  wire  _EVAL_2;
  wire  _EVAL_3;
  wire  _EVAL_4;
  wire  _EVAL_5;
  wire  _EVAL_7;
  wire [31:0] _EVAL_8;
  wire [4:0] _EVAL_10;
  wire  _EVAL_11;
  wire [1:0] _EVAL_12;
  wire  _EVAL_13;
  wire [3:0] _EVAL_14;
  wire  _EVAL_15;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire [2:0] _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire [2:0] _EVAL_25;
  wire  _EVAL_26;
  wire [3:0] _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  plicDomainWrapper__EVAL;
  wire  plicDomainWrapper__EVAL_0;
  wire  plicDomainWrapper__EVAL_1;
  wire  plicDomainWrapper__EVAL_2;
  wire [3:0] plicDomainWrapper__EVAL_3;
  wire  plicDomainWrapper__EVAL_4;
  wire  plicDomainWrapper__EVAL_5;
  wire  plicDomainWrapper__EVAL_6;
  wire  plicDomainWrapper__EVAL_7;
  wire  plicDomainWrapper__EVAL_8;
  wire  plicDomainWrapper__EVAL_9;
  wire  plicDomainWrapper__EVAL_10;
  wire [2:0] plicDomainWrapper__EVAL_11;
  wire  plicDomainWrapper__EVAL_12;
  wire  plicDomainWrapper__EVAL_13;
  wire  plicDomainWrapper__EVAL_14;
  wire  plicDomainWrapper__EVAL_15;
  wire  plicDomainWrapper__EVAL_16;
  wire  plicDomainWrapper__EVAL_17;
  wire  plicDomainWrapper__EVAL_18;
  wire  plicDomainWrapper__EVAL_19;
  wire  plicDomainWrapper__EVAL_20;
  wire  plicDomainWrapper__EVAL_21;
  wire  plicDomainWrapper__EVAL_22;
  wire  plicDomainWrapper__EVAL_23;
  wire  plicDomainWrapper__EVAL_24;
  wire  plicDomainWrapper__EVAL_25;
  wire  plicDomainWrapper__EVAL_26;
  wire  plicDomainWrapper__EVAL_27;
  wire  plicDomainWrapper__EVAL_28;
  wire  plicDomainWrapper__EVAL_29;
  wire  plicDomainWrapper__EVAL_30;
  wire [31:0] plicDomainWrapper__EVAL_31;
  wire  plicDomainWrapper__EVAL_32;
  wire  plicDomainWrapper__EVAL_33;
  wire  plicDomainWrapper__EVAL_34;
  wire  plicDomainWrapper__EVAL_35;
  wire  plicDomainWrapper__EVAL_36;
  wire  plicDomainWrapper__EVAL_37;
  wire  plicDomainWrapper__EVAL_38;
  wire  plicDomainWrapper__EVAL_39;
  wire  plicDomainWrapper__EVAL_40;
  wire  plicDomainWrapper__EVAL_41;
  wire  plicDomainWrapper__EVAL_42;
  wire [27:0] plicDomainWrapper__EVAL_43;
  wire [9:0] plicDomainWrapper__EVAL_44;
  wire  plicDomainWrapper__EVAL_45;
  wire  plicDomainWrapper__EVAL_46;
  wire  plicDomainWrapper__EVAL_47;
  wire  plicDomainWrapper__EVAL_48;
  wire  plicDomainWrapper__EVAL_49;
  wire  plicDomainWrapper__EVAL_50;
  wire  plicDomainWrapper__EVAL_51;
  wire  plicDomainWrapper__EVAL_52;
  wire  plicDomainWrapper__EVAL_53;
  wire  plicDomainWrapper__EVAL_54;
  wire  plicDomainWrapper__EVAL_55;
  wire  plicDomainWrapper__EVAL_56;
  wire  plicDomainWrapper__EVAL_57;
  wire  plicDomainWrapper__EVAL_58;
  wire  plicDomainWrapper__EVAL_59;
  wire  plicDomainWrapper__EVAL_60;
  wire  plicDomainWrapper__EVAL_61;
  wire  plicDomainWrapper__EVAL_62;
  wire  plicDomainWrapper__EVAL_63;
  wire  plicDomainWrapper__EVAL_64;
  wire  plicDomainWrapper__EVAL_65;
  wire  plicDomainWrapper__EVAL_66;
  wire  plicDomainWrapper__EVAL_67;
  wire  plicDomainWrapper__EVAL_68;
  wire  plicDomainWrapper__EVAL_69;
  wire  plicDomainWrapper__EVAL_70;
  wire  plicDomainWrapper__EVAL_71;
  wire  plicDomainWrapper__EVAL_72;
  wire  plicDomainWrapper__EVAL_73;
  wire  plicDomainWrapper__EVAL_74;
  wire  plicDomainWrapper__EVAL_75;
  wire  plicDomainWrapper__EVAL_76;
  wire  plicDomainWrapper__EVAL_77;
  wire  plicDomainWrapper__EVAL_78;
  wire  plicDomainWrapper__EVAL_79;
  wire [2:0] plicDomainWrapper__EVAL_80;
  wire  plicDomainWrapper__EVAL_81;
  wire  plicDomainWrapper__EVAL_82;
  wire  plicDomainWrapper__EVAL_83;
  wire  plicDomainWrapper__EVAL_84;
  wire  plicDomainWrapper__EVAL_85;
  wire  plicDomainWrapper__EVAL_86;
  wire  plicDomainWrapper__EVAL_87;
  wire  plicDomainWrapper__EVAL_88;
  wire  plicDomainWrapper__EVAL_89;
  wire  plicDomainWrapper__EVAL_90;
  wire  plicDomainWrapper__EVAL_91;
  wire  plicDomainWrapper__EVAL_92;
  wire  plicDomainWrapper__EVAL_93;
  wire  plicDomainWrapper__EVAL_94;
  wire  plicDomainWrapper__EVAL_95;
  wire  plicDomainWrapper__EVAL_96;
  wire  plicDomainWrapper__EVAL_97;
  wire  plicDomainWrapper__EVAL_98;
  wire  plicDomainWrapper__EVAL_99;
  wire  plicDomainWrapper__EVAL_100;
  wire  plicDomainWrapper__EVAL_101;
  wire [2:0] plicDomainWrapper__EVAL_102;
  wire  plicDomainWrapper__EVAL_103;
  wire  plicDomainWrapper__EVAL_104;
  wire  plicDomainWrapper__EVAL_105;
  wire  plicDomainWrapper__EVAL_106;
  wire  plicDomainWrapper__EVAL_107;
  wire  plicDomainWrapper__EVAL_108;
  wire  plicDomainWrapper__EVAL_109;
  wire  plicDomainWrapper__EVAL_110;
  wire  plicDomainWrapper__EVAL_111;
  wire  plicDomainWrapper__EVAL_112;
  wire  plicDomainWrapper__EVAL_113;
  wire  plicDomainWrapper__EVAL_114;
  wire  plicDomainWrapper__EVAL_115;
  wire  plicDomainWrapper__EVAL_116;
  wire [9:0] plicDomainWrapper__EVAL_117;
  wire  plicDomainWrapper__EVAL_118;
  wire  plicDomainWrapper__EVAL_119;
  wire  plicDomainWrapper__EVAL_120;
  wire  plicDomainWrapper__EVAL_121;
  wire  plicDomainWrapper__EVAL_122;
  wire  plicDomainWrapper__EVAL_123;
  wire  plicDomainWrapper__EVAL_124;
  wire  plicDomainWrapper__EVAL_125;
  wire  plicDomainWrapper__EVAL_126;
  wire  plicDomainWrapper__EVAL_127;
  wire [1:0] plicDomainWrapper__EVAL_128;
  wire  plicDomainWrapper__EVAL_129;
  wire  plicDomainWrapper__EVAL_130;
  wire  plicDomainWrapper__EVAL_131;
  wire  plicDomainWrapper__EVAL_132;
  wire  plicDomainWrapper__EVAL_133;
  wire  plicDomainWrapper__EVAL_134;
  wire  plicDomainWrapper__EVAL_135;
  wire  plicDomainWrapper__EVAL_136;
  wire  plicDomainWrapper__EVAL_137;
  wire  plicDomainWrapper__EVAL_138;
  wire  plicDomainWrapper__EVAL_139;
  wire [31:0] plicDomainWrapper__EVAL_140;
  wire [1:0] plicDomainWrapper__EVAL_141;
  wire  plicDomainWrapper__EVAL_142;
  wire  plicDomainWrapper__EVAL_143;
  wire  plicDomainWrapper__EVAL_144;
  wire  _EVAL_31;
  wire [4:0] _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire [3:0] _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire [31:0] subsystem_cbus__EVAL;
  wire [31:0] subsystem_cbus__EVAL_0;
  wire [31:0] subsystem_cbus__EVAL_1;
  wire [4:0] subsystem_cbus__EVAL_2;
  wire  subsystem_cbus__EVAL_3;
  wire [2:0] subsystem_cbus__EVAL_4;
  wire [4:0] subsystem_cbus__EVAL_5;
  wire [2:0] subsystem_cbus__EVAL_6;
  wire [1:0] subsystem_cbus__EVAL_7;
  wire [11:0] subsystem_cbus__EVAL_8;
  wire [1:0] subsystem_cbus__EVAL_9;
  wire [1:0] subsystem_cbus__EVAL_10;
  wire  subsystem_cbus__EVAL_11;
  wire [3:0] subsystem_cbus__EVAL_12;
  wire  subsystem_cbus__EVAL_13;
  wire [31:0] subsystem_cbus__EVAL_14;
  wire  subsystem_cbus__EVAL_15;
  wire  subsystem_cbus__EVAL_16;
  wire  subsystem_cbus__EVAL_17;
  wire  subsystem_cbus__EVAL_18;
  wire [31:0] subsystem_cbus__EVAL_19;
  wire [3:0] subsystem_cbus__EVAL_20;
  wire [9:0] subsystem_cbus__EVAL_21;
  wire [1:0] subsystem_cbus__EVAL_22;
  wire [2:0] subsystem_cbus__EVAL_23;
  wire [31:0] subsystem_cbus__EVAL_24;
  wire [1:0] subsystem_cbus__EVAL_25;
  wire [3:0] subsystem_cbus__EVAL_26;
  wire  subsystem_cbus__EVAL_27;
  wire [2:0] subsystem_cbus__EVAL_28;
  wire [2:0] subsystem_cbus__EVAL_29;
  wire [2:0] subsystem_cbus__EVAL_30;
  wire [2:0] subsystem_cbus__EVAL_31;
  wire [31:0] subsystem_cbus__EVAL_32;
  wire [9:0] subsystem_cbus__EVAL_33;
  wire [4:0] subsystem_cbus__EVAL_34;
  wire  subsystem_cbus__EVAL_35;
  wire [31:0] subsystem_cbus__EVAL_36;
  wire [2:0] subsystem_cbus__EVAL_37;
  wire [2:0] subsystem_cbus__EVAL_38;
  wire  subsystem_cbus__EVAL_39;
  wire  subsystem_cbus__EVAL_40;
  wire [2:0] subsystem_cbus__EVAL_41;
  wire [2:0] subsystem_cbus__EVAL_42;
  wire  subsystem_cbus__EVAL_43;
  wire [4:0] subsystem_cbus__EVAL_44;
  wire [14:0] subsystem_cbus__EVAL_45;
  wire  subsystem_cbus__EVAL_46;
  wire  subsystem_cbus__EVAL_47;
  wire [2:0] subsystem_cbus__EVAL_48;
  wire [31:0] subsystem_cbus__EVAL_49;
  wire  subsystem_cbus__EVAL_50;
  wire [9:0] subsystem_cbus__EVAL_51;
  wire [3:0] subsystem_cbus__EVAL_52;
  wire [9:0] subsystem_cbus__EVAL_53;
  wire [2:0] subsystem_cbus__EVAL_54;
  wire  subsystem_cbus__EVAL_55;
  wire  subsystem_cbus__EVAL_56;
  wire [1:0] subsystem_cbus__EVAL_57;
  wire  subsystem_cbus__EVAL_58;
  wire  subsystem_cbus__EVAL_59;
  wire [1:0] subsystem_cbus__EVAL_60;
  wire [3:0] subsystem_cbus__EVAL_61;
  wire [1:0] subsystem_cbus__EVAL_62;
  wire [2:0] subsystem_cbus__EVAL_63;
  wire  subsystem_cbus__EVAL_64;
  wire  subsystem_cbus__EVAL_65;
  wire  subsystem_cbus__EVAL_66;
  wire [2:0] subsystem_cbus__EVAL_67;
  wire [31:0] subsystem_cbus__EVAL_68;
  wire [4:0] subsystem_cbus__EVAL_69;
  wire  subsystem_cbus__EVAL_70;
  wire  subsystem_cbus__EVAL_71;
  wire [1:0] subsystem_cbus__EVAL_72;
  wire [1:0] subsystem_cbus__EVAL_73;
  wire [9:0] subsystem_cbus__EVAL_74;
  wire  subsystem_cbus__EVAL_75;
  wire  subsystem_cbus__EVAL_76;
  wire [25:0] subsystem_cbus__EVAL_77;
  wire  subsystem_cbus__EVAL_78;
  wire [31:0] subsystem_cbus__EVAL_79;
  wire  subsystem_cbus__EVAL_80;
  wire [27:0] subsystem_cbus__EVAL_81;
  wire  subsystem_cbus__EVAL_82;
  wire [31:0] subsystem_cbus__EVAL_83;
  wire [3:0] subsystem_cbus__EVAL_84;
  wire [4:0] subsystem_cbus__EVAL_85;
  wire  subsystem_cbus__EVAL_86;
  wire [2:0] subsystem_cbus__EVAL_87;
  wire [2:0] subsystem_cbus__EVAL_88;
  wire  subsystem_cbus__EVAL_89;
  wire [2:0] subsystem_cbus__EVAL_90;
  wire  subsystem_cbus__EVAL_91;
  wire [31:0] subsystem_cbus__EVAL_92;
  wire [3:0] subsystem_cbus__EVAL_93;
  wire [2:0] subsystem_cbus__EVAL_94;
  wire  subsystem_cbus__EVAL_95;
  wire  subsystem_cbus__EVAL_96;
  wire  subsystem_cbus__EVAL_97;
  wire [1:0] subsystem_cbus__EVAL_98;
  wire  subsystem_cbus__EVAL_99;
  wire [2:0] subsystem_cbus__EVAL_100;
  wire [31:0] subsystem_cbus__EVAL_101;
  wire  subsystem_cbus__EVAL_102;
  wire [31:0] subsystem_cbus__EVAL_103;
  wire [1:0] subsystem_cbus__EVAL_104;
  wire [29:0] subsystem_cbus__EVAL_105;
  wire [1:0] subsystem_cbus__EVAL_106;
  wire [1:0] subsystem_cbus__EVAL_107;
  wire [2:0] subsystem_cbus__EVAL_108;
  wire  subsystem_cbus__EVAL_109;
  wire [31:0] subsystem_cbus__EVAL_110;
  wire [2:0] subsystem_cbus__EVAL_111;
  wire  subsystem_cbus__EVAL_112;
  wire  subsystem_cbus__EVAL_113;
  wire [2:0] subsystem_cbus__EVAL_114;
  wire [31:0] subsystem_cbus__EVAL_115;
  wire [2:0] subsystem_cbus__EVAL_116;
  wire [3:0] subsystem_cbus__EVAL_117;
  wire [9:0] subsystem_cbus__EVAL_118;
  wire [31:0] subsystem_cbus__EVAL_119;
  wire  subsystem_cbus__EVAL_120;
  wire [3:0] subsystem_cbus__EVAL_121;
  wire [2:0] subsystem_cbus__EVAL_122;
  wire [9:0] subsystem_cbus__EVAL_123;
  wire [9:0] subsystem_cbus__EVAL_124;
  wire  subsystem_cbus__EVAL_125;
  wire [31:0] subsystem_cbus__EVAL_126;
  wire [3:0] subsystem_cbus__EVAL_127;
  wire  subsystem_cbus__EVAL_128;
  wire  subsystem_cbus__EVAL_129;
  wire  subsystem_cbus__EVAL_130;
  wire [2:0] subsystem_cbus__EVAL_131;
  wire  subsystem_cbus__EVAL_132;
  wire  subsystem_cbus__EVAL_133;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire [3:0] _EVAL_49;
  wire  _EVAL_51;
  wire [3:0] _EVAL_52;
  wire  intsource__EVAL;
  wire  intsource__EVAL_0;
  wire  intsource__EVAL_1;
  wire  intsource__EVAL_2;
  wire  intsource__EVAL_3;
  wire  intsource__EVAL_4;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire [2:0] _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire [3:0] _EVAL_61;
  wire  xbar_1__EVAL;
  wire  xbar_1__EVAL_0;
  wire [2:0] _EVAL_62;
  wire [3:0] _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_67;
  wire [4:0] _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_81;
  wire [31:0] _EVAL_82;
  wire  xbar__EVAL;
  wire  xbar__EVAL_0;
  wire  _EVAL_83;
  wire [2:0] _EVAL_84;
  wire [4:0] _EVAL_85;
  wire [31:0] _EVAL_86;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire [31:0] _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire [4:0] _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire [3:0] _EVAL_108;
  wire [3:0] _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire [31:0] _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  intsource_1__EVAL;
  wire  intsource_1__EVAL_0;
  wire  intsource_1__EVAL_1;
  wire  intsource_1__EVAL_2;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire [2:0] _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire [3:0] _EVAL_160;
  reg  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire [3:0] _EVAL_170;
  wire  _EVAL_171;
  wire [31:0] _EVAL_172;
  wire  intsink_3__EVAL;
  wire  intsink_3__EVAL_0;
  wire  _EVAL_174;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire [3:0] _EVAL_178;
  wire [31:0] _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire [1:0] _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire [4:0] _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire [4:0] _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire [1:0] _EVAL_195;
  wire [4:0] tile_prci_domain__EVAL;
  wire [2:0] tile_prci_domain__EVAL_0;
  wire  tile_prci_domain__EVAL_1;
  wire [31:0] tile_prci_domain__EVAL_2;
  wire  tile_prci_domain__EVAL_3;
  wire  tile_prci_domain__EVAL_4;
  wire [2:0] tile_prci_domain__EVAL_5;
  wire  tile_prci_domain__EVAL_6;
  wire [2:0] tile_prci_domain__EVAL_7;
  wire [31:0] tile_prci_domain__EVAL_8;
  wire [31:0] tile_prci_domain__EVAL_9;
  wire [1:0] tile_prci_domain__EVAL_10;
  wire [2:0] tile_prci_domain__EVAL_11;
  wire  tile_prci_domain__EVAL_12;
  wire [2:0] tile_prci_domain__EVAL_13;
  wire [3:0] tile_prci_domain__EVAL_14;
  wire [2:0] tile_prci_domain__EVAL_15;
  wire  tile_prci_domain__EVAL_16;
  wire [31:0] tile_prci_domain__EVAL_17;
  wire [31:0] tile_prci_domain__EVAL_18;
  wire  tile_prci_domain__EVAL_19;
  wire  tile_prci_domain__EVAL_20;
  wire  tile_prci_domain__EVAL_21;
  wire  tile_prci_domain__EVAL_22;
  wire [4:0] tile_prci_domain__EVAL_23;
  wire  tile_prci_domain__EVAL_24;
  wire [1:0] tile_prci_domain__EVAL_25;
  wire [2:0] tile_prci_domain__EVAL_26;
  wire [31:0] tile_prci_domain__EVAL_27;
  wire  tile_prci_domain__EVAL_28;
  wire  tile_prci_domain__EVAL_29;
  wire [2:0] tile_prci_domain__EVAL_30;
  wire [3:0] tile_prci_domain__EVAL_31;
  wire  tile_prci_domain__EVAL_32;
  wire [3:0] tile_prci_domain__EVAL_33;
  wire [31:0] tile_prci_domain__EVAL_34;
  wire  tile_prci_domain__EVAL_35;
  wire  tile_prci_domain__EVAL_36;
  wire  tile_prci_domain__EVAL_37;
  wire [3:0] tile_prci_domain__EVAL_38;
  wire  tile_prci_domain__EVAL_39;
  wire  tile_prci_domain__EVAL_40;
  wire [4:0] tile_prci_domain__EVAL_41;
  wire  tile_prci_domain__EVAL_42;
  wire  tile_prci_domain__EVAL_43;
  wire  tile_prci_domain__EVAL_44;
  wire  tile_prci_domain__EVAL_45;
  wire  tile_prci_domain__EVAL_46;
  wire [3:0] tile_prci_domain__EVAL_47;
  wire  tile_prci_domain__EVAL_48;
  wire [1:0] tile_prci_domain__EVAL_49;
  wire  tile_prci_domain__EVAL_50;
  wire [3:0] tile_prci_domain__EVAL_51;
  wire  tile_prci_domain__EVAL_52;
  wire  tile_prci_domain__EVAL_53;
  wire [2:0] tile_prci_domain__EVAL_54;
  wire [31:0] tile_prci_domain__EVAL_55;
  wire  tile_prci_domain__EVAL_56;
  wire  tile_prci_domain__EVAL_57;
  wire [2:0] tile_prci_domain__EVAL_58;
  wire  tile_prci_domain__EVAL_59;
  wire [2:0] tile_prci_domain__EVAL_60;
  wire  tile_prci_domain__EVAL_61;
  wire [1:0] tile_prci_domain__EVAL_62;
  wire  tile_prci_domain__EVAL_63;
  wire  tile_prci_domain__EVAL_64;
  wire [3:0] tile_prci_domain__EVAL_65;
  wire [2:0] tile_prci_domain__EVAL_66;
  wire [3:0] tile_prci_domain__EVAL_67;
  wire  tile_prci_domain__EVAL_68;
  wire [1:0] tile_prci_domain__EVAL_69;
  wire  tile_prci_domain__EVAL_70;
  wire [2:0] tile_prci_domain__EVAL_71;
  wire [3:0] tile_prci_domain__EVAL_72;
  wire  tile_prci_domain__EVAL_73;
  wire  tile_prci_domain__EVAL_74;
  wire [1:0] tile_prci_domain__EVAL_75;
  wire  tile_prci_domain__EVAL_76;
  wire  tile_prci_domain__EVAL_77;
  wire [3:0] tile_prci_domain__EVAL_78;
  wire [1:0] tile_prci_domain__EVAL_79;
  wire  tile_prci_domain__EVAL_80;
  wire [31:0] tile_prci_domain__EVAL_81;
  wire [2:0] tile_prci_domain__EVAL_82;
  wire [1:0] tile_prci_domain__EVAL_83;
  wire  tile_prci_domain__EVAL_84;
  wire  tile_prci_domain__EVAL_85;
  wire [31:0] tile_prci_domain__EVAL_86;
  wire [31:0] tile_prci_domain__EVAL_87;
  wire [31:0] tile_prci_domain__EVAL_88;
  wire  tile_prci_domain__EVAL_89;
  wire  tile_prci_domain__EVAL_90;
  wire [31:0] tile_prci_domain__EVAL_91;
  wire [1:0] tile_prci_domain__EVAL_92;
  wire  tile_prci_domain__EVAL_93;
  wire  tile_prci_domain__EVAL_94;
  wire  tile_prci_domain__EVAL_95;
  wire  tile_prci_domain__EVAL_96;
  wire [3:0] tile_prci_domain__EVAL_97;
  wire [1:0] tile_prci_domain__EVAL_98;
  wire  tile_prci_domain__EVAL_99;
  wire  tile_prci_domain__EVAL_100;
  wire [31:0] tile_prci_domain__EVAL_101;
  wire [3:0] tile_prci_domain__EVAL_102;
  wire [2:0] tile_prci_domain__EVAL_103;
  wire  tile_prci_domain__EVAL_104;
  wire [4:0] tile_prci_domain__EVAL_105;
  wire [2:0] tile_prci_domain__EVAL_106;
  wire  tile_prci_domain__EVAL_107;
  wire [31:0] tile_prci_domain__EVAL_108;
  wire [4:0] _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire [4:0] _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire [31:0] _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  reg  _EVAL_209;
  wire  _EVAL_210;
  wire  rtc_sync_chain__EVAL;
  wire  rtc_sync_chain__EVAL_0;
  wire  rtc_sync_chain__EVAL_1;
  wire  rtc_sync_chain__EVAL_2;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire [3:0] _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire [31:0] _EVAL_230;
  wire  _EVAL_231;
  wire [1:0] _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_236;
  wire  _EVAL_238;
  wire  tileHartIdNexusNode__EVAL;
  wire [4:0] _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_243;
  wire  _EVAL_245;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire [4:0] _EVAL_249;
  wire  intsink_2__EVAL;
  wire  intsink_2__EVAL_0;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire [3:0] _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire  subsystem_fbus__EVAL;
  wire [7:0] subsystem_fbus__EVAL_0;
  wire  subsystem_fbus__EVAL_1;
  wire  subsystem_fbus__EVAL_2;
  wire  subsystem_fbus__EVAL_3;
  wire  subsystem_fbus__EVAL_4;
  wire [2:0] subsystem_fbus__EVAL_5;
  wire  subsystem_fbus__EVAL_6;
  wire [3:0] subsystem_fbus__EVAL_7;
  wire  subsystem_fbus__EVAL_8;
  wire  subsystem_fbus__EVAL_9;
  wire  subsystem_fbus__EVAL_10;
  wire [31:0] subsystem_fbus__EVAL_11;
  wire  subsystem_fbus__EVAL_12;
  wire [31:0] subsystem_fbus__EVAL_13;
  wire  subsystem_fbus__EVAL_14;
  wire  subsystem_fbus__EVAL_15;
  wire [3:0] subsystem_fbus__EVAL_16;
  wire [2:0] subsystem_fbus__EVAL_17;
  wire  subsystem_fbus__EVAL_18;
  wire [2:0] subsystem_fbus__EVAL_19;
  wire [2:0] subsystem_fbus__EVAL_20;
  wire [3:0] subsystem_fbus__EVAL_21;
  wire  subsystem_fbus__EVAL_22;
  wire  subsystem_fbus__EVAL_23;
  wire [7:0] subsystem_fbus__EVAL_24;
  wire  subsystem_fbus__EVAL_25;
  wire  subsystem_fbus__EVAL_26;
  wire [3:0] subsystem_fbus__EVAL_27;
  wire [1:0] subsystem_fbus__EVAL_28;
  wire  subsystem_fbus__EVAL_29;
  wire  subsystem_fbus__EVAL_30;
  wire  subsystem_fbus__EVAL_31;
  wire [31:0] subsystem_fbus__EVAL_32;
  wire  subsystem_fbus__EVAL_33;
  wire  subsystem_fbus__EVAL_34;
  wire [31:0] subsystem_fbus__EVAL_35;
  wire  subsystem_fbus__EVAL_36;
  wire [2:0] subsystem_fbus__EVAL_37;
  wire [1:0] subsystem_fbus__EVAL_38;
  wire [31:0] subsystem_fbus__EVAL_39;
  wire [31:0] subsystem_fbus__EVAL_40;
  wire  subsystem_fbus__EVAL_41;
  wire [2:0] subsystem_fbus__EVAL_42;
  wire  subsystem_fbus__EVAL_43;
  wire [3:0] subsystem_fbus__EVAL_44;
  wire  subsystem_fbus__EVAL_45;
  wire [31:0] subsystem_fbus__EVAL_46;
  wire  subsystem_fbus__EVAL_47;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire [3:0] _EVAL_270;
  wire  _EVAL_271;
  wire [2:0] _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire [2:0] _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire [1:0] _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire [31:0] _EVAL_287;
  wire [31:0] _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_293;
  wire [2:0] _EVAL_294;
  wire  _EVAL_295;
  wire  ibus_int_bus__EVAL;
  wire  ibus_int_bus__EVAL_0;
  wire  ibus_int_bus__EVAL_1;
  wire  ibus_int_bus__EVAL_2;
  wire  ibus_int_bus__EVAL_3;
  wire  ibus_int_bus__EVAL_4;
  wire  ibus_int_bus__EVAL_5;
  wire  ibus_int_bus__EVAL_6;
  wire  ibus_int_bus__EVAL_7;
  wire  ibus_int_bus__EVAL_8;
  wire  ibus_int_bus__EVAL_9;
  wire  ibus_int_bus__EVAL_10;
  wire  ibus_int_bus__EVAL_11;
  wire  ibus_int_bus__EVAL_12;
  wire  ibus_int_bus__EVAL_13;
  wire  ibus_int_bus__EVAL_14;
  wire  ibus_int_bus__EVAL_15;
  wire  ibus_int_bus__EVAL_16;
  wire  ibus_int_bus__EVAL_17;
  wire  ibus_int_bus__EVAL_18;
  wire  ibus_int_bus__EVAL_19;
  wire  ibus_int_bus__EVAL_20;
  wire  ibus_int_bus__EVAL_21;
  wire  ibus_int_bus__EVAL_22;
  wire  ibus_int_bus__EVAL_23;
  wire  ibus_int_bus__EVAL_24;
  wire  ibus_int_bus__EVAL_25;
  wire  ibus_int_bus__EVAL_26;
  wire  ibus_int_bus__EVAL_27;
  wire  ibus_int_bus__EVAL_28;
  wire  ibus_int_bus__EVAL_29;
  wire  ibus_int_bus__EVAL_30;
  wire  ibus_int_bus__EVAL_31;
  wire  ibus_int_bus__EVAL_32;
  wire  ibus_int_bus__EVAL_33;
  wire  ibus_int_bus__EVAL_34;
  wire  ibus_int_bus__EVAL_35;
  wire  ibus_int_bus__EVAL_36;
  wire  ibus_int_bus__EVAL_37;
  wire  ibus_int_bus__EVAL_38;
  wire  ibus_int_bus__EVAL_39;
  wire  ibus_int_bus__EVAL_40;
  wire  ibus_int_bus__EVAL_41;
  wire  ibus_int_bus__EVAL_42;
  wire  ibus_int_bus__EVAL_43;
  wire  ibus_int_bus__EVAL_44;
  wire  ibus_int_bus__EVAL_45;
  wire  ibus_int_bus__EVAL_46;
  wire  ibus_int_bus__EVAL_47;
  wire  ibus_int_bus__EVAL_48;
  wire  ibus_int_bus__EVAL_49;
  wire  ibus_int_bus__EVAL_50;
  wire  ibus_int_bus__EVAL_51;
  wire  ibus_int_bus__EVAL_52;
  wire  ibus_int_bus__EVAL_53;
  wire  ibus_int_bus__EVAL_54;
  wire  ibus_int_bus__EVAL_55;
  wire  ibus_int_bus__EVAL_56;
  wire  ibus_int_bus__EVAL_57;
  wire  ibus_int_bus__EVAL_58;
  wire  ibus_int_bus__EVAL_59;
  wire  ibus_int_bus__EVAL_60;
  wire  ibus_int_bus__EVAL_61;
  wire  ibus_int_bus__EVAL_62;
  wire  ibus_int_bus__EVAL_63;
  wire  ibus_int_bus__EVAL_64;
  wire  ibus_int_bus__EVAL_65;
  wire  ibus_int_bus__EVAL_66;
  wire  ibus_int_bus__EVAL_67;
  wire  ibus_int_bus__EVAL_68;
  wire  ibus_int_bus__EVAL_69;
  wire  ibus_int_bus__EVAL_70;
  wire  ibus_int_bus__EVAL_71;
  wire  ibus_int_bus__EVAL_72;
  wire  ibus_int_bus__EVAL_73;
  wire  ibus_int_bus__EVAL_74;
  wire  ibus_int_bus__EVAL_75;
  wire  ibus_int_bus__EVAL_76;
  wire  ibus_int_bus__EVAL_77;
  wire  ibus_int_bus__EVAL_78;
  wire  ibus_int_bus__EVAL_79;
  wire  ibus_int_bus__EVAL_80;
  wire  ibus_int_bus__EVAL_81;
  wire  ibus_int_bus__EVAL_82;
  wire  ibus_int_bus__EVAL_83;
  wire  ibus_int_bus__EVAL_84;
  wire  ibus_int_bus__EVAL_85;
  wire  ibus_int_bus__EVAL_86;
  wire  ibus_int_bus__EVAL_87;
  wire  ibus_int_bus__EVAL_88;
  wire  ibus_int_bus__EVAL_89;
  wire  ibus_int_bus__EVAL_90;
  wire  ibus_int_bus__EVAL_91;
  wire  ibus_int_bus__EVAL_92;
  wire  ibus_int_bus__EVAL_93;
  wire  ibus_int_bus__EVAL_94;
  wire  ibus_int_bus__EVAL_95;
  wire  ibus_int_bus__EVAL_96;
  wire  ibus_int_bus__EVAL_97;
  wire  ibus_int_bus__EVAL_98;
  wire  ibus_int_bus__EVAL_99;
  wire  ibus_int_bus__EVAL_100;
  wire  ibus_int_bus__EVAL_101;
  wire  ibus_int_bus__EVAL_102;
  wire  ibus_int_bus__EVAL_103;
  wire  ibus_int_bus__EVAL_104;
  wire  ibus_int_bus__EVAL_105;
  wire  ibus_int_bus__EVAL_106;
  wire  ibus_int_bus__EVAL_107;
  wire  ibus_int_bus__EVAL_108;
  wire  ibus_int_bus__EVAL_109;
  wire  ibus_int_bus__EVAL_110;
  wire  ibus_int_bus__EVAL_111;
  wire  ibus_int_bus__EVAL_112;
  wire  ibus_int_bus__EVAL_113;
  wire  ibus_int_bus__EVAL_114;
  wire  ibus_int_bus__EVAL_115;
  wire  ibus_int_bus__EVAL_116;
  wire  ibus_int_bus__EVAL_117;
  wire  ibus_int_bus__EVAL_118;
  wire  ibus_int_bus__EVAL_119;
  wire  ibus_int_bus__EVAL_120;
  wire  ibus_int_bus__EVAL_121;
  wire  ibus_int_bus__EVAL_122;
  wire  ibus_int_bus__EVAL_123;
  wire  ibus_int_bus__EVAL_124;
  wire  ibus_int_bus__EVAL_125;
  wire  ibus_int_bus__EVAL_126;
  wire  ibus_int_bus__EVAL_127;
  wire  ibus_int_bus__EVAL_128;
  wire  ibus_int_bus__EVAL_129;
  wire  ibus_int_bus__EVAL_130;
  wire  ibus_int_bus__EVAL_131;
  wire  ibus_int_bus__EVAL_132;
  wire  ibus_int_bus__EVAL_133;
  wire  ibus_int_bus__EVAL_134;
  wire  ibus_int_bus__EVAL_135;
  wire  ibus_int_bus__EVAL_136;
  wire  ibus_int_bus__EVAL_137;
  wire  ibus_int_bus__EVAL_138;
  wire  ibus_int_bus__EVAL_139;
  wire  ibus_int_bus__EVAL_140;
  wire  ibus_int_bus__EVAL_141;
  wire  ibus_int_bus__EVAL_142;
  wire  ibus_int_bus__EVAL_143;
  wire  ibus_int_bus__EVAL_144;
  wire  ibus_int_bus__EVAL_145;
  wire  ibus_int_bus__EVAL_146;
  wire  ibus_int_bus__EVAL_147;
  wire  ibus_int_bus__EVAL_148;
  wire  ibus_int_bus__EVAL_149;
  wire  ibus_int_bus__EVAL_150;
  wire  ibus_int_bus__EVAL_151;
  wire  ibus_int_bus__EVAL_152;
  wire  ibus_int_bus__EVAL_153;
  wire  ibus_int_bus__EVAL_154;
  wire  ibus_int_bus__EVAL_155;
  wire  ibus_int_bus__EVAL_156;
  wire  ibus_int_bus__EVAL_157;
  wire  ibus_int_bus__EVAL_158;
  wire  ibus_int_bus__EVAL_159;
  wire  ibus_int_bus__EVAL_160;
  wire  ibus_int_bus__EVAL_161;
  wire  ibus_int_bus__EVAL_162;
  wire  ibus_int_bus__EVAL_163;
  wire  ibus_int_bus__EVAL_164;
  wire  ibus_int_bus__EVAL_165;
  wire  ibus_int_bus__EVAL_166;
  wire  ibus_int_bus__EVAL_167;
  wire  ibus_int_bus__EVAL_168;
  wire  ibus_int_bus__EVAL_169;
  wire  ibus_int_bus__EVAL_170;
  wire  ibus_int_bus__EVAL_171;
  wire  ibus_int_bus__EVAL_172;
  wire  ibus_int_bus__EVAL_173;
  wire  ibus_int_bus__EVAL_174;
  wire  ibus_int_bus__EVAL_175;
  wire  ibus_int_bus__EVAL_176;
  wire  ibus_int_bus__EVAL_177;
  wire  ibus_int_bus__EVAL_178;
  wire  ibus_int_bus__EVAL_179;
  wire  ibus_int_bus__EVAL_180;
  wire  ibus_int_bus__EVAL_181;
  wire  ibus_int_bus__EVAL_182;
  wire  ibus_int_bus__EVAL_183;
  wire  ibus_int_bus__EVAL_184;
  wire  ibus_int_bus__EVAL_185;
  wire  ibus_int_bus__EVAL_186;
  wire  ibus_int_bus__EVAL_187;
  wire  ibus_int_bus__EVAL_188;
  wire  ibus_int_bus__EVAL_189;
  wire  ibus_int_bus__EVAL_190;
  wire  ibus_int_bus__EVAL_191;
  wire  ibus_int_bus__EVAL_192;
  wire  ibus_int_bus__EVAL_193;
  wire  ibus_int_bus__EVAL_194;
  wire  ibus_int_bus__EVAL_195;
  wire  ibus_int_bus__EVAL_196;
  wire  ibus_int_bus__EVAL_197;
  wire  ibus_int_bus__EVAL_198;
  wire  ibus_int_bus__EVAL_199;
  wire  ibus_int_bus__EVAL_200;
  wire  ibus_int_bus__EVAL_201;
  wire  ibus_int_bus__EVAL_202;
  wire  ibus_int_bus__EVAL_203;
  wire  ibus_int_bus__EVAL_204;
  wire  ibus_int_bus__EVAL_205;
  wire  ibus_int_bus__EVAL_206;
  wire  ibus_int_bus__EVAL_207;
  wire  ibus_int_bus__EVAL_208;
  wire  ibus_int_bus__EVAL_209;
  wire  ibus_int_bus__EVAL_210;
  wire  ibus_int_bus__EVAL_211;
  wire  ibus_int_bus__EVAL_212;
  wire  ibus_int_bus__EVAL_213;
  wire  ibus_int_bus__EVAL_214;
  wire  ibus_int_bus__EVAL_215;
  wire  ibus_int_bus__EVAL_216;
  wire  ibus_int_bus__EVAL_217;
  wire  ibus_int_bus__EVAL_218;
  wire  ibus_int_bus__EVAL_219;
  wire  ibus_int_bus__EVAL_220;
  wire  ibus_int_bus__EVAL_221;
  wire  ibus_int_bus__EVAL_222;
  wire  ibus_int_bus__EVAL_223;
  wire  ibus_int_bus__EVAL_224;
  wire  ibus_int_bus__EVAL_225;
  wire  ibus_int_bus__EVAL_226;
  wire  ibus_int_bus__EVAL_227;
  wire  ibus_int_bus__EVAL_228;
  wire  ibus_int_bus__EVAL_229;
  wire  ibus_int_bus__EVAL_230;
  wire  ibus_int_bus__EVAL_231;
  wire  ibus_int_bus__EVAL_232;
  wire  ibus_int_bus__EVAL_233;
  wire  ibus_int_bus__EVAL_234;
  wire  ibus_int_bus__EVAL_235;
  wire  ibus_int_bus__EVAL_236;
  wire  ibus_int_bus__EVAL_237;
  wire  ibus_int_bus__EVAL_238;
  wire  ibus_int_bus__EVAL_239;
  wire  ibus_int_bus__EVAL_240;
  wire  ibus_int_bus__EVAL_241;
  wire  ibus_int_bus__EVAL_242;
  wire  ibus_int_bus__EVAL_243;
  wire  ibus_int_bus__EVAL_244;
  wire  ibus_int_bus__EVAL_245;
  wire  ibus_int_bus__EVAL_246;
  wire  ibus_int_bus__EVAL_247;
  wire  ibus_int_bus__EVAL_248;
  wire  ibus_int_bus__EVAL_249;
  wire  ibus_int_bus__EVAL_250;
  wire  ibus_int_bus__EVAL_251;
  wire  ibus_int_bus__EVAL_252;
  wire  _EVAL_296;
  wire  _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire  debug_1__EVAL;
  wire  debug_1__EVAL_0;
  wire  debug_1__EVAL_1;
  wire  debug_1__EVAL_2;
  wire  debug_1__EVAL_3;
  wire  debug_1__EVAL_4;
  wire [3:0] debug_1__EVAL_5;
  wire [1:0] debug_1__EVAL_6;
  wire  debug_1__EVAL_7;
  wire [3:0] debug_1__EVAL_8;
  wire  debug_1__EVAL_9;
  wire [2:0] debug_1__EVAL_10;
  wire  debug_1__EVAL_11;
  wire  debug_1__EVAL_12;
  wire  debug_1__EVAL_13;
  wire  debug_1__EVAL_14;
  wire [1:0] debug_1__EVAL_15;
  wire [9:0] debug_1__EVAL_16;
  wire [31:0] debug_1__EVAL_17;
  wire  debug_1__EVAL_18;
  wire  debug_1__EVAL_19;
  wire  debug_1__EVAL_20;
  wire  debug_1__EVAL_21;
  wire [7:0] debug_1__EVAL_22;
  wire [31:0] debug_1__EVAL_23;
  wire [2:0] debug_1__EVAL_24;
  wire [6:0] debug_1__EVAL_25;
  wire  debug_1__EVAL_26;
  wire [31:0] debug_1__EVAL_27;
  wire  debug_1__EVAL_28;
  wire [1:0] debug_1__EVAL_29;
  wire  debug_1__EVAL_30;
  wire [31:0] debug_1__EVAL_31;
  wire  debug_1__EVAL_32;
  wire  debug_1__EVAL_33;
  wire  debug_1__EVAL_34;
  wire [11:0] debug_1__EVAL_35;
  wire  debug_1__EVAL_36;
  wire  debug_1__EVAL_37;
  wire [2:0] debug_1__EVAL_38;
  wire [7:0] debug_1__EVAL_39;
  wire [2:0] debug_1__EVAL_40;
  wire [1:0] debug_1__EVAL_41;
  wire  debug_1__EVAL_42;
  wire  debug_1__EVAL_43;
  wire [9:0] debug_1__EVAL_44;
  wire [31:0] debug_1__EVAL_45;
  wire  _EVAL_302;
  wire  _EVAL_303;
  wire [2:0] _EVAL_304;
  wire  _EVAL_305;
  wire [2:0] _EVAL_307;
  wire  _EVAL_308;
  wire  _EVAL_309;
  wire  _EVAL_310;
  wire  _EVAL_311;
  wire  _EVAL_313;
  wire  _EVAL_314;
  wire [31:0] _EVAL_316;
  wire  _EVAL_317;
  wire  _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_320;
  wire  _EVAL_321;
  wire  _EVAL_322;
  wire  _EVAL_324;
  wire  _EVAL_325;
  wire  _EVAL_326;
  wire  _EVAL_327;
  wire  _EVAL_328;
  wire  _EVAL_329;
  wire  _EVAL_330;
  wire  _EVAL_331;
  wire  _EVAL_332;
  wire  _EVAL_334;
  wire  _EVAL_335;
  wire  _EVAL_337;
  wire [2:0] _EVAL_338;
  wire [4:0] _EVAL_340;
  wire  _EVAL_341;
  wire  _EVAL_342;
  wire  _EVAL_343;
  wire  _EVAL_344;
  wire  intsink_1__EVAL;
  wire  intsink_1__EVAL_0;
  wire  _EVAL_345;
  wire  _EVAL_346;
  wire  _EVAL_347;
  wire  _EVAL_349;
  wire [31:0] _EVAL_350;
  wire  _EVAL_351;
  wire  _EVAL_352;
  wire  _EVAL_353;
  wire [3:0] subsystem_sbus__EVAL;
  wire [1:0] subsystem_sbus__EVAL_0;
  wire  subsystem_sbus__EVAL_1;
  wire [1:0] subsystem_sbus__EVAL_2;
  wire  subsystem_sbus__EVAL_3;
  wire  subsystem_sbus__EVAL_4;
  wire  subsystem_sbus__EVAL_5;
  wire  subsystem_sbus__EVAL_6;
  wire [3:0] subsystem_sbus__EVAL_7;
  wire [3:0] subsystem_sbus__EVAL_8;
  wire  subsystem_sbus__EVAL_9;
  wire  subsystem_sbus__EVAL_10;
  wire [31:0] subsystem_sbus__EVAL_11;
  wire  subsystem_sbus__EVAL_12;
  wire  subsystem_sbus__EVAL_13;
  wire [31:0] subsystem_sbus__EVAL_14;
  wire [3:0] subsystem_sbus__EVAL_15;
  wire [30:0] subsystem_sbus__EVAL_16;
  wire [1:0] subsystem_sbus__EVAL_17;
  wire [31:0] subsystem_sbus__EVAL_18;
  wire  subsystem_sbus__EVAL_19;
  wire  subsystem_sbus__EVAL_20;
  wire [2:0] subsystem_sbus__EVAL_21;
  wire  subsystem_sbus__EVAL_22;
  wire  subsystem_sbus__EVAL_23;
  wire  subsystem_sbus__EVAL_24;
  wire [31:0] subsystem_sbus__EVAL_25;
  wire  subsystem_sbus__EVAL_26;
  wire  subsystem_sbus__EVAL_27;
  wire [3:0] subsystem_sbus__EVAL_28;
  wire [2:0] subsystem_sbus__EVAL_29;
  wire  subsystem_sbus__EVAL_30;
  wire  subsystem_sbus__EVAL_31;
  wire [1:0] subsystem_sbus__EVAL_32;
  wire  subsystem_sbus__EVAL_33;
  wire  subsystem_sbus__EVAL_34;
  wire  subsystem_sbus__EVAL_35;
  wire  subsystem_sbus__EVAL_36;
  wire [31:0] subsystem_sbus__EVAL_37;
  wire [1:0] subsystem_sbus__EVAL_38;
  wire [31:0] subsystem_sbus__EVAL_39;
  wire  subsystem_sbus__EVAL_40;
  wire [2:0] subsystem_sbus__EVAL_41;
  wire  subsystem_sbus__EVAL_42;
  wire  subsystem_sbus__EVAL_43;
  wire  subsystem_sbus__EVAL_44;
  wire  subsystem_sbus__EVAL_45;
  wire [1:0] subsystem_sbus__EVAL_46;
  wire [31:0] subsystem_sbus__EVAL_47;
  wire  subsystem_sbus__EVAL_48;
  wire [31:0] subsystem_sbus__EVAL_49;
  wire [2:0] subsystem_sbus__EVAL_50;
  wire [2:0] subsystem_sbus__EVAL_51;
  wire  subsystem_sbus__EVAL_52;
  wire  subsystem_sbus__EVAL_53;
  wire  subsystem_sbus__EVAL_54;
  wire [1:0] subsystem_sbus__EVAL_55;
  wire  subsystem_sbus__EVAL_56;
  wire  subsystem_sbus__EVAL_57;
  wire [1:0] subsystem_sbus__EVAL_58;
  wire [2:0] subsystem_sbus__EVAL_59;
  wire [3:0] subsystem_sbus__EVAL_60;
  wire  subsystem_sbus__EVAL_61;
  wire [3:0] subsystem_sbus__EVAL_62;
  wire  subsystem_sbus__EVAL_63;
  wire  subsystem_sbus__EVAL_64;
  wire [2:0] subsystem_sbus__EVAL_65;
  wire  subsystem_sbus__EVAL_66;
  wire  subsystem_sbus__EVAL_67;
  wire [4:0] subsystem_sbus__EVAL_68;
  wire  subsystem_sbus__EVAL_69;
  wire  subsystem_sbus__EVAL_70;
  wire  subsystem_sbus__EVAL_71;
  wire  subsystem_sbus__EVAL_72;
  wire [2:0] subsystem_sbus__EVAL_73;
  wire [3:0] subsystem_sbus__EVAL_74;
  wire  subsystem_sbus__EVAL_75;
  wire  subsystem_sbus__EVAL_76;
  wire [2:0] subsystem_sbus__EVAL_77;
  wire [2:0] subsystem_sbus__EVAL_78;
  wire [31:0] subsystem_sbus__EVAL_79;
  wire  subsystem_sbus__EVAL_80;
  wire [31:0] subsystem_sbus__EVAL_81;
  wire [3:0] subsystem_sbus__EVAL_82;
  wire [1:0] subsystem_sbus__EVAL_83;
  wire  subsystem_sbus__EVAL_84;
  wire  subsystem_sbus__EVAL_85;
  wire [31:0] subsystem_sbus__EVAL_86;
  wire  subsystem_sbus__EVAL_87;
  wire [3:0] subsystem_sbus__EVAL_88;
  wire  subsystem_sbus__EVAL_89;
  wire [31:0] subsystem_sbus__EVAL_90;
  wire  subsystem_sbus__EVAL_91;
  wire [3:0] subsystem_sbus__EVAL_92;
  wire [2:0] subsystem_sbus__EVAL_93;
  wire [3:0] subsystem_sbus__EVAL_94;
  wire  subsystem_sbus__EVAL_95;
  wire  subsystem_sbus__EVAL_96;
  wire [3:0] subsystem_sbus__EVAL_97;
  wire [3:0] subsystem_sbus__EVAL_98;
  wire [31:0] subsystem_sbus__EVAL_99;
  wire  subsystem_sbus__EVAL_100;
  wire [2:0] subsystem_sbus__EVAL_101;
  wire  subsystem_sbus__EVAL_102;
  wire  subsystem_sbus__EVAL_103;
  wire  subsystem_sbus__EVAL_104;
  wire  subsystem_sbus__EVAL_105;
  wire  subsystem_sbus__EVAL_106;
  wire  subsystem_sbus__EVAL_107;
  wire [2:0] subsystem_sbus__EVAL_108;
  wire [3:0] subsystem_sbus__EVAL_109;
  wire [2:0] subsystem_sbus__EVAL_110;
  wire  subsystem_sbus__EVAL_111;
  wire [3:0] subsystem_sbus__EVAL_112;
  wire  subsystem_sbus__EVAL_113;
  wire [3:0] subsystem_sbus__EVAL_114;
  wire [4:0] subsystem_sbus__EVAL_115;
  wire  subsystem_sbus__EVAL_116;
  wire [31:0] subsystem_sbus__EVAL_117;
  wire  subsystem_sbus__EVAL_118;
  wire [2:0] _EVAL_354;
  wire  _EVAL_355;
  wire [2:0] _EVAL_356;
  wire [2:0] _EVAL_357;
  wire  xbar_2__EVAL;
  wire  xbar_2__EVAL_0;
  wire  _EVAL_358;
  wire [3:0] _EVAL_359;
  wire  _EVAL_361;
  wire  _EVAL_362;
  wire [2:0] _EVAL_363;
  wire  _EVAL_364;
  wire  _EVAL_365;
  wire  _EVAL_366;
  wire [4:0] _EVAL_367;
  wire  _EVAL_368;
  wire  _EVAL_369;
  wire  _EVAL_370;
  wire  _EVAL_371;
  wire [31:0] dtm__EVAL;
  wire  dtm__EVAL_0;
  wire  dtm__EVAL_1;
  wire  dtm__EVAL_2;
  wire  dtm__EVAL_3;
  wire  dtm__EVAL_4;
  wire [6:0] dtm__EVAL_5;
  wire  dtm__EVAL_6;
  wire  dtm__EVAL_7;
  wire [10:0] dtm__EVAL_8;
  wire  dtm__EVAL_9;
  wire  dtm__EVAL_10;
  wire  dtm__EVAL_11;
  wire [1:0] dtm__EVAL_12;
  wire [31:0] dtm__EVAL_13;
  wire [3:0] dtm__EVAL_14;
  wire [15:0] dtm__EVAL_15;
  wire [1:0] dtm__EVAL_16;
  wire  _EVAL_372;
  wire  _EVAL_373;
  wire  _EVAL_374;
  wire  _EVAL_375;
  wire  _EVAL_376;
  wire [3:0] _EVAL_377;
  wire [31:0] _EVAL_378;
  wire  _EVAL_379;
  wire  _EVAL_380;
  wire  _EVAL_381;
  wire  _EVAL_382;
  wire  _EVAL_383;
  wire  _EVAL_384;
  wire  _EVAL_385;
  wire [3:0] _EVAL_386;
  wire  _EVAL_387;
  wire [31:0] _EVAL_388;
  wire  _EVAL_389;
  wire  _EVAL_391;
  wire  _EVAL_392;
  wire  _EVAL_393;
  wire  _EVAL_394;
  wire  _EVAL_395;
  wire  testIndicator_auto_control_xing_in_a_ready;
  wire  testIndicator_auto_control_xing_in_a_valid;
  wire [2:0] testIndicator_auto_control_xing_in_a_bits_opcode;
  wire [2:0] testIndicator_auto_control_xing_in_a_bits_param;
  wire [1:0] testIndicator_auto_control_xing_in_a_bits_size;
  wire [9:0] testIndicator_auto_control_xing_in_a_bits_source;
  wire [14:0] testIndicator_auto_control_xing_in_a_bits_address;
  wire [3:0] testIndicator_auto_control_xing_in_a_bits_mask;
  wire [31:0] testIndicator_auto_control_xing_in_a_bits_data;
  wire  testIndicator_auto_control_xing_in_a_bits_corrupt;
  wire  testIndicator_auto_control_xing_in_d_ready;
  wire  testIndicator_auto_control_xing_in_d_valid;
  wire [2:0] testIndicator_auto_control_xing_in_d_bits_opcode;
  wire [1:0] testIndicator_auto_control_xing_in_d_bits_size;
  wire [9:0] testIndicator_auto_control_xing_in_d_bits_source;
  wire [31:0] testIndicator_auto_control_xing_in_d_bits_data;
  wire  testIndicator_clock;
  wire  testIndicator_reset;
  wire [4:0] _EVAL_396;
  wire [31:0] _EVAL_397;
  wire [31:0] _EVAL_398;
  wire  _EVAL_399;
  wire  _EVAL_400;
  wire  _EVAL_401;
  wire  _EVAL_402;
  wire  _EVAL_403;
  wire  _EVAL_404;
  wire [2:0] _EVAL_405;
  wire  _EVAL_406;
  wire  xbar_3__EVAL;
  wire  xbar_3__EVAL_0;
  wire [2:0] _EVAL_407;
  wire [3:0] _EVAL_408;
  wire  _EVAL_409;
  wire [31:0] _EVAL_410;
  wire [31:0] _EVAL_411;
  wire  _EVAL_412;
  wire [31:0] _EVAL_413;
  wire [3:0] _EVAL_414;
  wire  _EVAL_415;
  wire  _EVAL_416;
  wire [2:0] _EVAL_418;
  wire  _EVAL_419;
  wire  _EVAL_420;
  wire [3:0] _EVAL_421;
  wire [31:0] _EVAL_422;
  wire  _EVAL_423;
  wire [1:0] _EVAL_424;
  wire  _EVAL_425;
  wire  _EVAL_426;
  wire [1:0] clint__EVAL;
  wire [3:0] clint__EVAL_0;
  wire [2:0] clint__EVAL_1;
  wire [9:0] clint__EVAL_2;
  wire [1:0] clint__EVAL_3;
  wire [31:0] clint__EVAL_4;
  wire  clint__EVAL_5;
  wire  clint__EVAL_6;
  wire [9:0] clint__EVAL_7;
  wire [31:0] clint__EVAL_8;
  wire  clint__EVAL_9;
  wire  clint__EVAL_10;
  wire [25:0] clint__EVAL_11;
  wire  clint__EVAL_12;
  wire  clint__EVAL_13;
  wire [2:0] clint__EVAL_14;
  wire  clint__EVAL_15;
  wire [2:0] clint__EVAL_16;
  wire  clint__EVAL_17;
  wire  clint__EVAL_18;
  wire  clint__EVAL_19;
  wire [4:0] _EVAL_429;
  wire  _EVAL_430;
  wire  _EVAL_431;
  wire [2:0] _EVAL_432;
  wire  _EVAL_434;
  wire  _EVAL_436;
  wire  _EVAL_437;
  wire  _EVAL_438;
  wire [4:0] _EVAL_440;
  wire  _EVAL_441;
  wire [2:0] _EVAL_442;
  wire  _EVAL_443;
  wire  _EVAL_444;
  wire  _EVAL_445;
  wire  _EVAL_446;
  wire  _EVAL_448;
  wire  _EVAL_449;
  wire  _EVAL_450;
  wire [2:0] _EVAL_451;
  wire  intsource_2__EVAL;
  wire  intsource_2__EVAL_0;
  wire  intsource_2__EVAL_1;
  wire  intsource_2__EVAL_2;
  wire  intsource_2__EVAL_3;
  wire  intsource_2__EVAL_4;
  wire  intsource_2__EVAL_5;
  wire  intsource_2__EVAL_6;
  wire  intsource_2__EVAL_7;
  wire  intsource_2__EVAL_8;
  wire  intsource_2__EVAL_9;
  wire  intsource_2__EVAL_10;
  wire  intsource_2__EVAL_11;
  wire  intsource_2__EVAL_12;
  wire  intsource_2__EVAL_13;
  wire  intsource_2__EVAL_14;
  wire  intsource_2__EVAL_15;
  wire  intsource_2__EVAL_16;
  wire  intsource_2__EVAL_17;
  wire  intsource_2__EVAL_18;
  wire  intsource_2__EVAL_19;
  wire  intsource_2__EVAL_20;
  wire  intsource_2__EVAL_21;
  wire  intsource_2__EVAL_22;
  wire  intsource_2__EVAL_23;
  wire  intsource_2__EVAL_24;
  wire  intsource_2__EVAL_25;
  wire  intsource_2__EVAL_26;
  wire  intsource_2__EVAL_27;
  wire  intsource_2__EVAL_28;
  wire  intsource_2__EVAL_29;
  wire  intsource_2__EVAL_30;
  wire  _EVAL_452;
  wire  _EVAL_453;
  wire  _EVAL_454;
  wire  _EVAL_455;
  wire [2:0] _EVAL_456;
  wire  intsink_4__EVAL;
  wire  intsink_4__EVAL_0;
  wire  _EVAL_458;
  wire  _EVAL_460;
  wire [31:0] _EVAL_461;
  wire [1:0] _EVAL_462;
  wire [31:0] _EVAL_463;
  wire  _EVAL_464;
  wire  _EVAL_465;
  wire  _EVAL_466;
  wire  _EVAL_467;
  wire  _EVAL_468;
  wire  _EVAL_469;
  wire  _EVAL_471;
  wire  _EVAL_472;
  wire  _EVAL_473;
  wire  _EVAL_474;
  wire  _EVAL_475;
  wire  _EVAL_476;
  wire  _EVAL_477;
  wire  _EVAL_478;
  wire  _EVAL_479;
  wire  _EVAL_480;
  wire [3:0] _EVAL_481;
  wire [3:0] _EVAL_482;
  wire  _EVAL_483;
  wire  _EVAL_484;
  wire  _EVAL_485;
  wire  _EVAL_486;
  wire  _EVAL_487;
  wire  _EVAL_488;
  wire  _EVAL_489;
  wire  _EVAL_490;
  wire  _EVAL_491;
  wire [31:0] _EVAL_492;
  wire  _EVAL_493;
  wire  _EVAL_494;
  wire  _EVAL_496;
  wire  _EVAL_497;
  wire  _EVAL_498;
  wire  _EVAL_499;
  wire  _EVAL_500;
  wire  _EVAL_502;
  wire  _EVAL_503;
  wire  _EVAL_504;
  wire  _EVAL_505;
  wire [3:0] _EVAL_506;
  wire [2:0] _EVAL_507;
  wire [1:0] _EVAL_508;
  wire  _EVAL_509;
  wire  _EVAL_510;
  wire  _EVAL_511;
  _EVAL_100 plicDomainWrapper (
    ._EVAL(plicDomainWrapper__EVAL),
    ._EVAL_0(plicDomainWrapper__EVAL_0),
    ._EVAL_1(plicDomainWrapper__EVAL_1),
    ._EVAL_2(plicDomainWrapper__EVAL_2),
    ._EVAL_3(plicDomainWrapper__EVAL_3),
    ._EVAL_4(plicDomainWrapper__EVAL_4),
    ._EVAL_5(plicDomainWrapper__EVAL_5),
    ._EVAL_6(plicDomainWrapper__EVAL_6),
    ._EVAL_7(plicDomainWrapper__EVAL_7),
    ._EVAL_8(plicDomainWrapper__EVAL_8),
    ._EVAL_9(plicDomainWrapper__EVAL_9),
    ._EVAL_10(plicDomainWrapper__EVAL_10),
    ._EVAL_11(plicDomainWrapper__EVAL_11),
    ._EVAL_12(plicDomainWrapper__EVAL_12),
    ._EVAL_13(plicDomainWrapper__EVAL_13),
    ._EVAL_14(plicDomainWrapper__EVAL_14),
    ._EVAL_15(plicDomainWrapper__EVAL_15),
    ._EVAL_16(plicDomainWrapper__EVAL_16),
    ._EVAL_17(plicDomainWrapper__EVAL_17),
    ._EVAL_18(plicDomainWrapper__EVAL_18),
    ._EVAL_19(plicDomainWrapper__EVAL_19),
    ._EVAL_20(plicDomainWrapper__EVAL_20),
    ._EVAL_21(plicDomainWrapper__EVAL_21),
    ._EVAL_22(plicDomainWrapper__EVAL_22),
    ._EVAL_23(plicDomainWrapper__EVAL_23),
    ._EVAL_24(plicDomainWrapper__EVAL_24),
    ._EVAL_25(plicDomainWrapper__EVAL_25),
    ._EVAL_26(plicDomainWrapper__EVAL_26),
    ._EVAL_27(plicDomainWrapper__EVAL_27),
    ._EVAL_28(plicDomainWrapper__EVAL_28),
    ._EVAL_29(plicDomainWrapper__EVAL_29),
    ._EVAL_30(plicDomainWrapper__EVAL_30),
    ._EVAL_31(plicDomainWrapper__EVAL_31),
    ._EVAL_32(plicDomainWrapper__EVAL_32),
    ._EVAL_33(plicDomainWrapper__EVAL_33),
    ._EVAL_34(plicDomainWrapper__EVAL_34),
    ._EVAL_35(plicDomainWrapper__EVAL_35),
    ._EVAL_36(plicDomainWrapper__EVAL_36),
    ._EVAL_37(plicDomainWrapper__EVAL_37),
    ._EVAL_38(plicDomainWrapper__EVAL_38),
    ._EVAL_39(plicDomainWrapper__EVAL_39),
    ._EVAL_40(plicDomainWrapper__EVAL_40),
    ._EVAL_41(plicDomainWrapper__EVAL_41),
    ._EVAL_42(plicDomainWrapper__EVAL_42),
    ._EVAL_43(plicDomainWrapper__EVAL_43),
    ._EVAL_44(plicDomainWrapper__EVAL_44),
    ._EVAL_45(plicDomainWrapper__EVAL_45),
    ._EVAL_46(plicDomainWrapper__EVAL_46),
    ._EVAL_47(plicDomainWrapper__EVAL_47),
    ._EVAL_48(plicDomainWrapper__EVAL_48),
    ._EVAL_49(plicDomainWrapper__EVAL_49),
    ._EVAL_50(plicDomainWrapper__EVAL_50),
    ._EVAL_51(plicDomainWrapper__EVAL_51),
    ._EVAL_52(plicDomainWrapper__EVAL_52),
    ._EVAL_53(plicDomainWrapper__EVAL_53),
    ._EVAL_54(plicDomainWrapper__EVAL_54),
    ._EVAL_55(plicDomainWrapper__EVAL_55),
    ._EVAL_56(plicDomainWrapper__EVAL_56),
    ._EVAL_57(plicDomainWrapper__EVAL_57),
    ._EVAL_58(plicDomainWrapper__EVAL_58),
    ._EVAL_59(plicDomainWrapper__EVAL_59),
    ._EVAL_60(plicDomainWrapper__EVAL_60),
    ._EVAL_61(plicDomainWrapper__EVAL_61),
    ._EVAL_62(plicDomainWrapper__EVAL_62),
    ._EVAL_63(plicDomainWrapper__EVAL_63),
    ._EVAL_64(plicDomainWrapper__EVAL_64),
    ._EVAL_65(plicDomainWrapper__EVAL_65),
    ._EVAL_66(plicDomainWrapper__EVAL_66),
    ._EVAL_67(plicDomainWrapper__EVAL_67),
    ._EVAL_68(plicDomainWrapper__EVAL_68),
    ._EVAL_69(plicDomainWrapper__EVAL_69),
    ._EVAL_70(plicDomainWrapper__EVAL_70),
    ._EVAL_71(plicDomainWrapper__EVAL_71),
    ._EVAL_72(plicDomainWrapper__EVAL_72),
    ._EVAL_73(plicDomainWrapper__EVAL_73),
    ._EVAL_74(plicDomainWrapper__EVAL_74),
    ._EVAL_75(plicDomainWrapper__EVAL_75),
    ._EVAL_76(plicDomainWrapper__EVAL_76),
    ._EVAL_77(plicDomainWrapper__EVAL_77),
    ._EVAL_78(plicDomainWrapper__EVAL_78),
    ._EVAL_79(plicDomainWrapper__EVAL_79),
    ._EVAL_80(plicDomainWrapper__EVAL_80),
    ._EVAL_81(plicDomainWrapper__EVAL_81),
    ._EVAL_82(plicDomainWrapper__EVAL_82),
    ._EVAL_83(plicDomainWrapper__EVAL_83),
    ._EVAL_84(plicDomainWrapper__EVAL_84),
    ._EVAL_85(plicDomainWrapper__EVAL_85),
    ._EVAL_86(plicDomainWrapper__EVAL_86),
    ._EVAL_87(plicDomainWrapper__EVAL_87),
    ._EVAL_88(plicDomainWrapper__EVAL_88),
    ._EVAL_89(plicDomainWrapper__EVAL_89),
    ._EVAL_90(plicDomainWrapper__EVAL_90),
    ._EVAL_91(plicDomainWrapper__EVAL_91),
    ._EVAL_92(plicDomainWrapper__EVAL_92),
    ._EVAL_93(plicDomainWrapper__EVAL_93),
    ._EVAL_94(plicDomainWrapper__EVAL_94),
    ._EVAL_95(plicDomainWrapper__EVAL_95),
    ._EVAL_96(plicDomainWrapper__EVAL_96),
    ._EVAL_97(plicDomainWrapper__EVAL_97),
    ._EVAL_98(plicDomainWrapper__EVAL_98),
    ._EVAL_99(plicDomainWrapper__EVAL_99),
    ._EVAL_100(plicDomainWrapper__EVAL_100),
    ._EVAL_101(plicDomainWrapper__EVAL_101),
    ._EVAL_102(plicDomainWrapper__EVAL_102),
    ._EVAL_103(plicDomainWrapper__EVAL_103),
    ._EVAL_104(plicDomainWrapper__EVAL_104),
    ._EVAL_105(plicDomainWrapper__EVAL_105),
    ._EVAL_106(plicDomainWrapper__EVAL_106),
    ._EVAL_107(plicDomainWrapper__EVAL_107),
    ._EVAL_108(plicDomainWrapper__EVAL_108),
    ._EVAL_109(plicDomainWrapper__EVAL_109),
    ._EVAL_110(plicDomainWrapper__EVAL_110),
    ._EVAL_111(plicDomainWrapper__EVAL_111),
    ._EVAL_112(plicDomainWrapper__EVAL_112),
    ._EVAL_113(plicDomainWrapper__EVAL_113),
    ._EVAL_114(plicDomainWrapper__EVAL_114),
    ._EVAL_115(plicDomainWrapper__EVAL_115),
    ._EVAL_116(plicDomainWrapper__EVAL_116),
    ._EVAL_117(plicDomainWrapper__EVAL_117),
    ._EVAL_118(plicDomainWrapper__EVAL_118),
    ._EVAL_119(plicDomainWrapper__EVAL_119),
    ._EVAL_120(plicDomainWrapper__EVAL_120),
    ._EVAL_121(plicDomainWrapper__EVAL_121),
    ._EVAL_122(plicDomainWrapper__EVAL_122),
    ._EVAL_123(plicDomainWrapper__EVAL_123),
    ._EVAL_124(plicDomainWrapper__EVAL_124),
    ._EVAL_125(plicDomainWrapper__EVAL_125),
    ._EVAL_126(plicDomainWrapper__EVAL_126),
    ._EVAL_127(plicDomainWrapper__EVAL_127),
    ._EVAL_128(plicDomainWrapper__EVAL_128),
    ._EVAL_129(plicDomainWrapper__EVAL_129),
    ._EVAL_130(plicDomainWrapper__EVAL_130),
    ._EVAL_131(plicDomainWrapper__EVAL_131),
    ._EVAL_132(plicDomainWrapper__EVAL_132),
    ._EVAL_133(plicDomainWrapper__EVAL_133),
    ._EVAL_134(plicDomainWrapper__EVAL_134),
    ._EVAL_135(plicDomainWrapper__EVAL_135),
    ._EVAL_136(plicDomainWrapper__EVAL_136),
    ._EVAL_137(plicDomainWrapper__EVAL_137),
    ._EVAL_138(plicDomainWrapper__EVAL_138),
    ._EVAL_139(plicDomainWrapper__EVAL_139),
    ._EVAL_140(plicDomainWrapper__EVAL_140),
    ._EVAL_141(plicDomainWrapper__EVAL_141),
    ._EVAL_142(plicDomainWrapper__EVAL_142),
    ._EVAL_143(plicDomainWrapper__EVAL_143),
    ._EVAL_144(plicDomainWrapper__EVAL_144)
  );
  _EVAL_94 subsystem_cbus (
    ._EVAL(subsystem_cbus__EVAL),
    ._EVAL_0(subsystem_cbus__EVAL_0),
    ._EVAL_1(subsystem_cbus__EVAL_1),
    ._EVAL_2(subsystem_cbus__EVAL_2),
    ._EVAL_3(subsystem_cbus__EVAL_3),
    ._EVAL_4(subsystem_cbus__EVAL_4),
    ._EVAL_5(subsystem_cbus__EVAL_5),
    ._EVAL_6(subsystem_cbus__EVAL_6),
    ._EVAL_7(subsystem_cbus__EVAL_7),
    ._EVAL_8(subsystem_cbus__EVAL_8),
    ._EVAL_9(subsystem_cbus__EVAL_9),
    ._EVAL_10(subsystem_cbus__EVAL_10),
    ._EVAL_11(subsystem_cbus__EVAL_11),
    ._EVAL_12(subsystem_cbus__EVAL_12),
    ._EVAL_13(subsystem_cbus__EVAL_13),
    ._EVAL_14(subsystem_cbus__EVAL_14),
    ._EVAL_15(subsystem_cbus__EVAL_15),
    ._EVAL_16(subsystem_cbus__EVAL_16),
    ._EVAL_17(subsystem_cbus__EVAL_17),
    ._EVAL_18(subsystem_cbus__EVAL_18),
    ._EVAL_19(subsystem_cbus__EVAL_19),
    ._EVAL_20(subsystem_cbus__EVAL_20),
    ._EVAL_21(subsystem_cbus__EVAL_21),
    ._EVAL_22(subsystem_cbus__EVAL_22),
    ._EVAL_23(subsystem_cbus__EVAL_23),
    ._EVAL_24(subsystem_cbus__EVAL_24),
    ._EVAL_25(subsystem_cbus__EVAL_25),
    ._EVAL_26(subsystem_cbus__EVAL_26),
    ._EVAL_27(subsystem_cbus__EVAL_27),
    ._EVAL_28(subsystem_cbus__EVAL_28),
    ._EVAL_29(subsystem_cbus__EVAL_29),
    ._EVAL_30(subsystem_cbus__EVAL_30),
    ._EVAL_31(subsystem_cbus__EVAL_31),
    ._EVAL_32(subsystem_cbus__EVAL_32),
    ._EVAL_33(subsystem_cbus__EVAL_33),
    ._EVAL_34(subsystem_cbus__EVAL_34),
    ._EVAL_35(subsystem_cbus__EVAL_35),
    ._EVAL_36(subsystem_cbus__EVAL_36),
    ._EVAL_37(subsystem_cbus__EVAL_37),
    ._EVAL_38(subsystem_cbus__EVAL_38),
    ._EVAL_39(subsystem_cbus__EVAL_39),
    ._EVAL_40(subsystem_cbus__EVAL_40),
    ._EVAL_41(subsystem_cbus__EVAL_41),
    ._EVAL_42(subsystem_cbus__EVAL_42),
    ._EVAL_43(subsystem_cbus__EVAL_43),
    ._EVAL_44(subsystem_cbus__EVAL_44),
    ._EVAL_45(subsystem_cbus__EVAL_45),
    ._EVAL_46(subsystem_cbus__EVAL_46),
    ._EVAL_47(subsystem_cbus__EVAL_47),
    ._EVAL_48(subsystem_cbus__EVAL_48),
    ._EVAL_49(subsystem_cbus__EVAL_49),
    ._EVAL_50(subsystem_cbus__EVAL_50),
    ._EVAL_51(subsystem_cbus__EVAL_51),
    ._EVAL_52(subsystem_cbus__EVAL_52),
    ._EVAL_53(subsystem_cbus__EVAL_53),
    ._EVAL_54(subsystem_cbus__EVAL_54),
    ._EVAL_55(subsystem_cbus__EVAL_55),
    ._EVAL_56(subsystem_cbus__EVAL_56),
    ._EVAL_57(subsystem_cbus__EVAL_57),
    ._EVAL_58(subsystem_cbus__EVAL_58),
    ._EVAL_59(subsystem_cbus__EVAL_59),
    ._EVAL_60(subsystem_cbus__EVAL_60),
    ._EVAL_61(subsystem_cbus__EVAL_61),
    ._EVAL_62(subsystem_cbus__EVAL_62),
    ._EVAL_63(subsystem_cbus__EVAL_63),
    ._EVAL_64(subsystem_cbus__EVAL_64),
    ._EVAL_65(subsystem_cbus__EVAL_65),
    ._EVAL_66(subsystem_cbus__EVAL_66),
    ._EVAL_67(subsystem_cbus__EVAL_67),
    ._EVAL_68(subsystem_cbus__EVAL_68),
    ._EVAL_69(subsystem_cbus__EVAL_69),
    ._EVAL_70(subsystem_cbus__EVAL_70),
    ._EVAL_71(subsystem_cbus__EVAL_71),
    ._EVAL_72(subsystem_cbus__EVAL_72),
    ._EVAL_73(subsystem_cbus__EVAL_73),
    ._EVAL_74(subsystem_cbus__EVAL_74),
    ._EVAL_75(subsystem_cbus__EVAL_75),
    ._EVAL_76(subsystem_cbus__EVAL_76),
    ._EVAL_77(subsystem_cbus__EVAL_77),
    ._EVAL_78(subsystem_cbus__EVAL_78),
    ._EVAL_79(subsystem_cbus__EVAL_79),
    ._EVAL_80(subsystem_cbus__EVAL_80),
    ._EVAL_81(subsystem_cbus__EVAL_81),
    ._EVAL_82(subsystem_cbus__EVAL_82),
    ._EVAL_83(subsystem_cbus__EVAL_83),
    ._EVAL_84(subsystem_cbus__EVAL_84),
    ._EVAL_85(subsystem_cbus__EVAL_85),
    ._EVAL_86(subsystem_cbus__EVAL_86),
    ._EVAL_87(subsystem_cbus__EVAL_87),
    ._EVAL_88(subsystem_cbus__EVAL_88),
    ._EVAL_89(subsystem_cbus__EVAL_89),
    ._EVAL_90(subsystem_cbus__EVAL_90),
    ._EVAL_91(subsystem_cbus__EVAL_91),
    ._EVAL_92(subsystem_cbus__EVAL_92),
    ._EVAL_93(subsystem_cbus__EVAL_93),
    ._EVAL_94(subsystem_cbus__EVAL_94),
    ._EVAL_95(subsystem_cbus__EVAL_95),
    ._EVAL_96(subsystem_cbus__EVAL_96),
    ._EVAL_97(subsystem_cbus__EVAL_97),
    ._EVAL_98(subsystem_cbus__EVAL_98),
    ._EVAL_99(subsystem_cbus__EVAL_99),
    ._EVAL_100(subsystem_cbus__EVAL_100),
    ._EVAL_101(subsystem_cbus__EVAL_101),
    ._EVAL_102(subsystem_cbus__EVAL_102),
    ._EVAL_103(subsystem_cbus__EVAL_103),
    ._EVAL_104(subsystem_cbus__EVAL_104),
    ._EVAL_105(subsystem_cbus__EVAL_105),
    ._EVAL_106(subsystem_cbus__EVAL_106),
    ._EVAL_107(subsystem_cbus__EVAL_107),
    ._EVAL_108(subsystem_cbus__EVAL_108),
    ._EVAL_109(subsystem_cbus__EVAL_109),
    ._EVAL_110(subsystem_cbus__EVAL_110),
    ._EVAL_111(subsystem_cbus__EVAL_111),
    ._EVAL_112(subsystem_cbus__EVAL_112),
    ._EVAL_113(subsystem_cbus__EVAL_113),
    ._EVAL_114(subsystem_cbus__EVAL_114),
    ._EVAL_115(subsystem_cbus__EVAL_115),
    ._EVAL_116(subsystem_cbus__EVAL_116),
    ._EVAL_117(subsystem_cbus__EVAL_117),
    ._EVAL_118(subsystem_cbus__EVAL_118),
    ._EVAL_119(subsystem_cbus__EVAL_119),
    ._EVAL_120(subsystem_cbus__EVAL_120),
    ._EVAL_121(subsystem_cbus__EVAL_121),
    ._EVAL_122(subsystem_cbus__EVAL_122),
    ._EVAL_123(subsystem_cbus__EVAL_123),
    ._EVAL_124(subsystem_cbus__EVAL_124),
    ._EVAL_125(subsystem_cbus__EVAL_125),
    ._EVAL_126(subsystem_cbus__EVAL_126),
    ._EVAL_127(subsystem_cbus__EVAL_127),
    ._EVAL_128(subsystem_cbus__EVAL_128),
    ._EVAL_129(subsystem_cbus__EVAL_129),
    ._EVAL_130(subsystem_cbus__EVAL_130),
    ._EVAL_131(subsystem_cbus__EVAL_131),
    ._EVAL_132(subsystem_cbus__EVAL_132),
    ._EVAL_133(subsystem_cbus__EVAL_133)
  );
  _EVAL_189 intsource (
    ._EVAL(intsource__EVAL),
    ._EVAL_0(intsource__EVAL_0),
    ._EVAL_1(intsource__EVAL_1),
    ._EVAL_2(intsource__EVAL_2),
    ._EVAL_3(intsource__EVAL_3),
    ._EVAL_4(intsource__EVAL_4)
  );
  _EVAL_186 xbar_1 (
    ._EVAL(xbar_1__EVAL),
    ._EVAL_0(xbar_1__EVAL_0)
  );
  _EVAL_186 xbar (
    ._EVAL(xbar__EVAL),
    ._EVAL_0(xbar__EVAL_0)
  );
  _EVAL_191 intsource_1 (
    ._EVAL(intsource_1__EVAL),
    ._EVAL_0(intsource_1__EVAL_0),
    ._EVAL_1(intsource_1__EVAL_1),
    ._EVAL_2(intsource_1__EVAL_2)
  );
  _EVAL_193 intsink_3 (
    ._EVAL(intsink_3__EVAL),
    ._EVAL_0(intsink_3__EVAL_0)
  );
  _EVAL_149 tile_prci_domain (
    ._EVAL(tile_prci_domain__EVAL),
    ._EVAL_0(tile_prci_domain__EVAL_0),
    ._EVAL_1(tile_prci_domain__EVAL_1),
    ._EVAL_2(tile_prci_domain__EVAL_2),
    ._EVAL_3(tile_prci_domain__EVAL_3),
    ._EVAL_4(tile_prci_domain__EVAL_4),
    ._EVAL_5(tile_prci_domain__EVAL_5),
    ._EVAL_6(tile_prci_domain__EVAL_6),
    ._EVAL_7(tile_prci_domain__EVAL_7),
    ._EVAL_8(tile_prci_domain__EVAL_8),
    ._EVAL_9(tile_prci_domain__EVAL_9),
    ._EVAL_10(tile_prci_domain__EVAL_10),
    ._EVAL_11(tile_prci_domain__EVAL_11),
    ._EVAL_12(tile_prci_domain__EVAL_12),
    ._EVAL_13(tile_prci_domain__EVAL_13),
    ._EVAL_14(tile_prci_domain__EVAL_14),
    ._EVAL_15(tile_prci_domain__EVAL_15),
    ._EVAL_16(tile_prci_domain__EVAL_16),
    ._EVAL_17(tile_prci_domain__EVAL_17),
    ._EVAL_18(tile_prci_domain__EVAL_18),
    ._EVAL_19(tile_prci_domain__EVAL_19),
    ._EVAL_20(tile_prci_domain__EVAL_20),
    ._EVAL_21(tile_prci_domain__EVAL_21),
    ._EVAL_22(tile_prci_domain__EVAL_22),
    ._EVAL_23(tile_prci_domain__EVAL_23),
    ._EVAL_24(tile_prci_domain__EVAL_24),
    ._EVAL_25(tile_prci_domain__EVAL_25),
    ._EVAL_26(tile_prci_domain__EVAL_26),
    ._EVAL_27(tile_prci_domain__EVAL_27),
    ._EVAL_28(tile_prci_domain__EVAL_28),
    ._EVAL_29(tile_prci_domain__EVAL_29),
    ._EVAL_30(tile_prci_domain__EVAL_30),
    ._EVAL_31(tile_prci_domain__EVAL_31),
    ._EVAL_32(tile_prci_domain__EVAL_32),
    ._EVAL_33(tile_prci_domain__EVAL_33),
    ._EVAL_34(tile_prci_domain__EVAL_34),
    ._EVAL_35(tile_prci_domain__EVAL_35),
    ._EVAL_36(tile_prci_domain__EVAL_36),
    ._EVAL_37(tile_prci_domain__EVAL_37),
    ._EVAL_38(tile_prci_domain__EVAL_38),
    ._EVAL_39(tile_prci_domain__EVAL_39),
    ._EVAL_40(tile_prci_domain__EVAL_40),
    ._EVAL_41(tile_prci_domain__EVAL_41),
    ._EVAL_42(tile_prci_domain__EVAL_42),
    ._EVAL_43(tile_prci_domain__EVAL_43),
    ._EVAL_44(tile_prci_domain__EVAL_44),
    ._EVAL_45(tile_prci_domain__EVAL_45),
    ._EVAL_46(tile_prci_domain__EVAL_46),
    ._EVAL_47(tile_prci_domain__EVAL_47),
    ._EVAL_48(tile_prci_domain__EVAL_48),
    ._EVAL_49(tile_prci_domain__EVAL_49),
    ._EVAL_50(tile_prci_domain__EVAL_50),
    ._EVAL_51(tile_prci_domain__EVAL_51),
    ._EVAL_52(tile_prci_domain__EVAL_52),
    ._EVAL_53(tile_prci_domain__EVAL_53),
    ._EVAL_54(tile_prci_domain__EVAL_54),
    ._EVAL_55(tile_prci_domain__EVAL_55),
    ._EVAL_56(tile_prci_domain__EVAL_56),
    ._EVAL_57(tile_prci_domain__EVAL_57),
    ._EVAL_58(tile_prci_domain__EVAL_58),
    ._EVAL_59(tile_prci_domain__EVAL_59),
    ._EVAL_60(tile_prci_domain__EVAL_60),
    ._EVAL_61(tile_prci_domain__EVAL_61),
    ._EVAL_62(tile_prci_domain__EVAL_62),
    ._EVAL_63(tile_prci_domain__EVAL_63),
    ._EVAL_64(tile_prci_domain__EVAL_64),
    ._EVAL_65(tile_prci_domain__EVAL_65),
    ._EVAL_66(tile_prci_domain__EVAL_66),
    ._EVAL_67(tile_prci_domain__EVAL_67),
    ._EVAL_68(tile_prci_domain__EVAL_68),
    ._EVAL_69(tile_prci_domain__EVAL_69),
    ._EVAL_70(tile_prci_domain__EVAL_70),
    ._EVAL_71(tile_prci_domain__EVAL_71),
    ._EVAL_72(tile_prci_domain__EVAL_72),
    ._EVAL_73(tile_prci_domain__EVAL_73),
    ._EVAL_74(tile_prci_domain__EVAL_74),
    ._EVAL_75(tile_prci_domain__EVAL_75),
    ._EVAL_76(tile_prci_domain__EVAL_76),
    ._EVAL_77(tile_prci_domain__EVAL_77),
    ._EVAL_78(tile_prci_domain__EVAL_78),
    ._EVAL_79(tile_prci_domain__EVAL_79),
    ._EVAL_80(tile_prci_domain__EVAL_80),
    ._EVAL_81(tile_prci_domain__EVAL_81),
    ._EVAL_82(tile_prci_domain__EVAL_82),
    ._EVAL_83(tile_prci_domain__EVAL_83),
    ._EVAL_84(tile_prci_domain__EVAL_84),
    ._EVAL_85(tile_prci_domain__EVAL_85),
    ._EVAL_86(tile_prci_domain__EVAL_86),
    ._EVAL_87(tile_prci_domain__EVAL_87),
    ._EVAL_88(tile_prci_domain__EVAL_88),
    ._EVAL_89(tile_prci_domain__EVAL_89),
    ._EVAL_90(tile_prci_domain__EVAL_90),
    ._EVAL_91(tile_prci_domain__EVAL_91),
    ._EVAL_92(tile_prci_domain__EVAL_92),
    ._EVAL_93(tile_prci_domain__EVAL_93),
    ._EVAL_94(tile_prci_domain__EVAL_94),
    ._EVAL_95(tile_prci_domain__EVAL_95),
    ._EVAL_96(tile_prci_domain__EVAL_96),
    ._EVAL_97(tile_prci_domain__EVAL_97),
    ._EVAL_98(tile_prci_domain__EVAL_98),
    ._EVAL_99(tile_prci_domain__EVAL_99),
    ._EVAL_100(tile_prci_domain__EVAL_100),
    ._EVAL_101(tile_prci_domain__EVAL_101),
    ._EVAL_102(tile_prci_domain__EVAL_102),
    ._EVAL_103(tile_prci_domain__EVAL_103),
    ._EVAL_104(tile_prci_domain__EVAL_104),
    ._EVAL_105(tile_prci_domain__EVAL_105),
    ._EVAL_106(tile_prci_domain__EVAL_106),
    ._EVAL_107(tile_prci_domain__EVAL_107),
    ._EVAL_108(tile_prci_domain__EVAL_108)
  );
  _EVAL_206 rtc_sync_chain (
    ._EVAL(rtc_sync_chain__EVAL),
    ._EVAL_0(rtc_sync_chain__EVAL_0),
    ._EVAL_1(rtc_sync_chain__EVAL_1),
    ._EVAL_2(rtc_sync_chain__EVAL_2)
  );
  _EVAL_187 tileHartIdNexusNode (
    ._EVAL(tileHartIdNexusNode__EVAL)
  );
  _EVAL_193 intsink_2 (
    ._EVAL(intsink_2__EVAL),
    ._EVAL_0(intsink_2__EVAL_0)
  );
  _EVAL_41 subsystem_fbus (
    ._EVAL(subsystem_fbus__EVAL),
    ._EVAL_0(subsystem_fbus__EVAL_0),
    ._EVAL_1(subsystem_fbus__EVAL_1),
    ._EVAL_2(subsystem_fbus__EVAL_2),
    ._EVAL_3(subsystem_fbus__EVAL_3),
    ._EVAL_4(subsystem_fbus__EVAL_4),
    ._EVAL_5(subsystem_fbus__EVAL_5),
    ._EVAL_6(subsystem_fbus__EVAL_6),
    ._EVAL_7(subsystem_fbus__EVAL_7),
    ._EVAL_8(subsystem_fbus__EVAL_8),
    ._EVAL_9(subsystem_fbus__EVAL_9),
    ._EVAL_10(subsystem_fbus__EVAL_10),
    ._EVAL_11(subsystem_fbus__EVAL_11),
    ._EVAL_12(subsystem_fbus__EVAL_12),
    ._EVAL_13(subsystem_fbus__EVAL_13),
    ._EVAL_14(subsystem_fbus__EVAL_14),
    ._EVAL_15(subsystem_fbus__EVAL_15),
    ._EVAL_16(subsystem_fbus__EVAL_16),
    ._EVAL_17(subsystem_fbus__EVAL_17),
    ._EVAL_18(subsystem_fbus__EVAL_18),
    ._EVAL_19(subsystem_fbus__EVAL_19),
    ._EVAL_20(subsystem_fbus__EVAL_20),
    ._EVAL_21(subsystem_fbus__EVAL_21),
    ._EVAL_22(subsystem_fbus__EVAL_22),
    ._EVAL_23(subsystem_fbus__EVAL_23),
    ._EVAL_24(subsystem_fbus__EVAL_24),
    ._EVAL_25(subsystem_fbus__EVAL_25),
    ._EVAL_26(subsystem_fbus__EVAL_26),
    ._EVAL_27(subsystem_fbus__EVAL_27),
    ._EVAL_28(subsystem_fbus__EVAL_28),
    ._EVAL_29(subsystem_fbus__EVAL_29),
    ._EVAL_30(subsystem_fbus__EVAL_30),
    ._EVAL_31(subsystem_fbus__EVAL_31),
    ._EVAL_32(subsystem_fbus__EVAL_32),
    ._EVAL_33(subsystem_fbus__EVAL_33),
    ._EVAL_34(subsystem_fbus__EVAL_34),
    ._EVAL_35(subsystem_fbus__EVAL_35),
    ._EVAL_36(subsystem_fbus__EVAL_36),
    ._EVAL_37(subsystem_fbus__EVAL_37),
    ._EVAL_38(subsystem_fbus__EVAL_38),
    ._EVAL_39(subsystem_fbus__EVAL_39),
    ._EVAL_40(subsystem_fbus__EVAL_40),
    ._EVAL_41(subsystem_fbus__EVAL_41),
    ._EVAL_42(subsystem_fbus__EVAL_42),
    ._EVAL_43(subsystem_fbus__EVAL_43),
    ._EVAL_44(subsystem_fbus__EVAL_44),
    ._EVAL_45(subsystem_fbus__EVAL_45),
    ._EVAL_46(subsystem_fbus__EVAL_46),
    ._EVAL_47(subsystem_fbus__EVAL_47)
  );
  _EVAL ibus_int_bus (
    ._EVAL(ibus_int_bus__EVAL),
    ._EVAL_0(ibus_int_bus__EVAL_0),
    ._EVAL_1(ibus_int_bus__EVAL_1),
    ._EVAL_2(ibus_int_bus__EVAL_2),
    ._EVAL_3(ibus_int_bus__EVAL_3),
    ._EVAL_4(ibus_int_bus__EVAL_4),
    ._EVAL_5(ibus_int_bus__EVAL_5),
    ._EVAL_6(ibus_int_bus__EVAL_6),
    ._EVAL_7(ibus_int_bus__EVAL_7),
    ._EVAL_8(ibus_int_bus__EVAL_8),
    ._EVAL_9(ibus_int_bus__EVAL_9),
    ._EVAL_10(ibus_int_bus__EVAL_10),
    ._EVAL_11(ibus_int_bus__EVAL_11),
    ._EVAL_12(ibus_int_bus__EVAL_12),
    ._EVAL_13(ibus_int_bus__EVAL_13),
    ._EVAL_14(ibus_int_bus__EVAL_14),
    ._EVAL_15(ibus_int_bus__EVAL_15),
    ._EVAL_16(ibus_int_bus__EVAL_16),
    ._EVAL_17(ibus_int_bus__EVAL_17),
    ._EVAL_18(ibus_int_bus__EVAL_18),
    ._EVAL_19(ibus_int_bus__EVAL_19),
    ._EVAL_20(ibus_int_bus__EVAL_20),
    ._EVAL_21(ibus_int_bus__EVAL_21),
    ._EVAL_22(ibus_int_bus__EVAL_22),
    ._EVAL_23(ibus_int_bus__EVAL_23),
    ._EVAL_24(ibus_int_bus__EVAL_24),
    ._EVAL_25(ibus_int_bus__EVAL_25),
    ._EVAL_26(ibus_int_bus__EVAL_26),
    ._EVAL_27(ibus_int_bus__EVAL_27),
    ._EVAL_28(ibus_int_bus__EVAL_28),
    ._EVAL_29(ibus_int_bus__EVAL_29),
    ._EVAL_30(ibus_int_bus__EVAL_30),
    ._EVAL_31(ibus_int_bus__EVAL_31),
    ._EVAL_32(ibus_int_bus__EVAL_32),
    ._EVAL_33(ibus_int_bus__EVAL_33),
    ._EVAL_34(ibus_int_bus__EVAL_34),
    ._EVAL_35(ibus_int_bus__EVAL_35),
    ._EVAL_36(ibus_int_bus__EVAL_36),
    ._EVAL_37(ibus_int_bus__EVAL_37),
    ._EVAL_38(ibus_int_bus__EVAL_38),
    ._EVAL_39(ibus_int_bus__EVAL_39),
    ._EVAL_40(ibus_int_bus__EVAL_40),
    ._EVAL_41(ibus_int_bus__EVAL_41),
    ._EVAL_42(ibus_int_bus__EVAL_42),
    ._EVAL_43(ibus_int_bus__EVAL_43),
    ._EVAL_44(ibus_int_bus__EVAL_44),
    ._EVAL_45(ibus_int_bus__EVAL_45),
    ._EVAL_46(ibus_int_bus__EVAL_46),
    ._EVAL_47(ibus_int_bus__EVAL_47),
    ._EVAL_48(ibus_int_bus__EVAL_48),
    ._EVAL_49(ibus_int_bus__EVAL_49),
    ._EVAL_50(ibus_int_bus__EVAL_50),
    ._EVAL_51(ibus_int_bus__EVAL_51),
    ._EVAL_52(ibus_int_bus__EVAL_52),
    ._EVAL_53(ibus_int_bus__EVAL_53),
    ._EVAL_54(ibus_int_bus__EVAL_54),
    ._EVAL_55(ibus_int_bus__EVAL_55),
    ._EVAL_56(ibus_int_bus__EVAL_56),
    ._EVAL_57(ibus_int_bus__EVAL_57),
    ._EVAL_58(ibus_int_bus__EVAL_58),
    ._EVAL_59(ibus_int_bus__EVAL_59),
    ._EVAL_60(ibus_int_bus__EVAL_60),
    ._EVAL_61(ibus_int_bus__EVAL_61),
    ._EVAL_62(ibus_int_bus__EVAL_62),
    ._EVAL_63(ibus_int_bus__EVAL_63),
    ._EVAL_64(ibus_int_bus__EVAL_64),
    ._EVAL_65(ibus_int_bus__EVAL_65),
    ._EVAL_66(ibus_int_bus__EVAL_66),
    ._EVAL_67(ibus_int_bus__EVAL_67),
    ._EVAL_68(ibus_int_bus__EVAL_68),
    ._EVAL_69(ibus_int_bus__EVAL_69),
    ._EVAL_70(ibus_int_bus__EVAL_70),
    ._EVAL_71(ibus_int_bus__EVAL_71),
    ._EVAL_72(ibus_int_bus__EVAL_72),
    ._EVAL_73(ibus_int_bus__EVAL_73),
    ._EVAL_74(ibus_int_bus__EVAL_74),
    ._EVAL_75(ibus_int_bus__EVAL_75),
    ._EVAL_76(ibus_int_bus__EVAL_76),
    ._EVAL_77(ibus_int_bus__EVAL_77),
    ._EVAL_78(ibus_int_bus__EVAL_78),
    ._EVAL_79(ibus_int_bus__EVAL_79),
    ._EVAL_80(ibus_int_bus__EVAL_80),
    ._EVAL_81(ibus_int_bus__EVAL_81),
    ._EVAL_82(ibus_int_bus__EVAL_82),
    ._EVAL_83(ibus_int_bus__EVAL_83),
    ._EVAL_84(ibus_int_bus__EVAL_84),
    ._EVAL_85(ibus_int_bus__EVAL_85),
    ._EVAL_86(ibus_int_bus__EVAL_86),
    ._EVAL_87(ibus_int_bus__EVAL_87),
    ._EVAL_88(ibus_int_bus__EVAL_88),
    ._EVAL_89(ibus_int_bus__EVAL_89),
    ._EVAL_90(ibus_int_bus__EVAL_90),
    ._EVAL_91(ibus_int_bus__EVAL_91),
    ._EVAL_92(ibus_int_bus__EVAL_92),
    ._EVAL_93(ibus_int_bus__EVAL_93),
    ._EVAL_94(ibus_int_bus__EVAL_94),
    ._EVAL_95(ibus_int_bus__EVAL_95),
    ._EVAL_96(ibus_int_bus__EVAL_96),
    ._EVAL_97(ibus_int_bus__EVAL_97),
    ._EVAL_98(ibus_int_bus__EVAL_98),
    ._EVAL_99(ibus_int_bus__EVAL_99),
    ._EVAL_100(ibus_int_bus__EVAL_100),
    ._EVAL_101(ibus_int_bus__EVAL_101),
    ._EVAL_102(ibus_int_bus__EVAL_102),
    ._EVAL_103(ibus_int_bus__EVAL_103),
    ._EVAL_104(ibus_int_bus__EVAL_104),
    ._EVAL_105(ibus_int_bus__EVAL_105),
    ._EVAL_106(ibus_int_bus__EVAL_106),
    ._EVAL_107(ibus_int_bus__EVAL_107),
    ._EVAL_108(ibus_int_bus__EVAL_108),
    ._EVAL_109(ibus_int_bus__EVAL_109),
    ._EVAL_110(ibus_int_bus__EVAL_110),
    ._EVAL_111(ibus_int_bus__EVAL_111),
    ._EVAL_112(ibus_int_bus__EVAL_112),
    ._EVAL_113(ibus_int_bus__EVAL_113),
    ._EVAL_114(ibus_int_bus__EVAL_114),
    ._EVAL_115(ibus_int_bus__EVAL_115),
    ._EVAL_116(ibus_int_bus__EVAL_116),
    ._EVAL_117(ibus_int_bus__EVAL_117),
    ._EVAL_118(ibus_int_bus__EVAL_118),
    ._EVAL_119(ibus_int_bus__EVAL_119),
    ._EVAL_120(ibus_int_bus__EVAL_120),
    ._EVAL_121(ibus_int_bus__EVAL_121),
    ._EVAL_122(ibus_int_bus__EVAL_122),
    ._EVAL_123(ibus_int_bus__EVAL_123),
    ._EVAL_124(ibus_int_bus__EVAL_124),
    ._EVAL_125(ibus_int_bus__EVAL_125),
    ._EVAL_126(ibus_int_bus__EVAL_126),
    ._EVAL_127(ibus_int_bus__EVAL_127),
    ._EVAL_128(ibus_int_bus__EVAL_128),
    ._EVAL_129(ibus_int_bus__EVAL_129),
    ._EVAL_130(ibus_int_bus__EVAL_130),
    ._EVAL_131(ibus_int_bus__EVAL_131),
    ._EVAL_132(ibus_int_bus__EVAL_132),
    ._EVAL_133(ibus_int_bus__EVAL_133),
    ._EVAL_134(ibus_int_bus__EVAL_134),
    ._EVAL_135(ibus_int_bus__EVAL_135),
    ._EVAL_136(ibus_int_bus__EVAL_136),
    ._EVAL_137(ibus_int_bus__EVAL_137),
    ._EVAL_138(ibus_int_bus__EVAL_138),
    ._EVAL_139(ibus_int_bus__EVAL_139),
    ._EVAL_140(ibus_int_bus__EVAL_140),
    ._EVAL_141(ibus_int_bus__EVAL_141),
    ._EVAL_142(ibus_int_bus__EVAL_142),
    ._EVAL_143(ibus_int_bus__EVAL_143),
    ._EVAL_144(ibus_int_bus__EVAL_144),
    ._EVAL_145(ibus_int_bus__EVAL_145),
    ._EVAL_146(ibus_int_bus__EVAL_146),
    ._EVAL_147(ibus_int_bus__EVAL_147),
    ._EVAL_148(ibus_int_bus__EVAL_148),
    ._EVAL_149(ibus_int_bus__EVAL_149),
    ._EVAL_150(ibus_int_bus__EVAL_150),
    ._EVAL_151(ibus_int_bus__EVAL_151),
    ._EVAL_152(ibus_int_bus__EVAL_152),
    ._EVAL_153(ibus_int_bus__EVAL_153),
    ._EVAL_154(ibus_int_bus__EVAL_154),
    ._EVAL_155(ibus_int_bus__EVAL_155),
    ._EVAL_156(ibus_int_bus__EVAL_156),
    ._EVAL_157(ibus_int_bus__EVAL_157),
    ._EVAL_158(ibus_int_bus__EVAL_158),
    ._EVAL_159(ibus_int_bus__EVAL_159),
    ._EVAL_160(ibus_int_bus__EVAL_160),
    ._EVAL_161(ibus_int_bus__EVAL_161),
    ._EVAL_162(ibus_int_bus__EVAL_162),
    ._EVAL_163(ibus_int_bus__EVAL_163),
    ._EVAL_164(ibus_int_bus__EVAL_164),
    ._EVAL_165(ibus_int_bus__EVAL_165),
    ._EVAL_166(ibus_int_bus__EVAL_166),
    ._EVAL_167(ibus_int_bus__EVAL_167),
    ._EVAL_168(ibus_int_bus__EVAL_168),
    ._EVAL_169(ibus_int_bus__EVAL_169),
    ._EVAL_170(ibus_int_bus__EVAL_170),
    ._EVAL_171(ibus_int_bus__EVAL_171),
    ._EVAL_172(ibus_int_bus__EVAL_172),
    ._EVAL_173(ibus_int_bus__EVAL_173),
    ._EVAL_174(ibus_int_bus__EVAL_174),
    ._EVAL_175(ibus_int_bus__EVAL_175),
    ._EVAL_176(ibus_int_bus__EVAL_176),
    ._EVAL_177(ibus_int_bus__EVAL_177),
    ._EVAL_178(ibus_int_bus__EVAL_178),
    ._EVAL_179(ibus_int_bus__EVAL_179),
    ._EVAL_180(ibus_int_bus__EVAL_180),
    ._EVAL_181(ibus_int_bus__EVAL_181),
    ._EVAL_182(ibus_int_bus__EVAL_182),
    ._EVAL_183(ibus_int_bus__EVAL_183),
    ._EVAL_184(ibus_int_bus__EVAL_184),
    ._EVAL_185(ibus_int_bus__EVAL_185),
    ._EVAL_186(ibus_int_bus__EVAL_186),
    ._EVAL_187(ibus_int_bus__EVAL_187),
    ._EVAL_188(ibus_int_bus__EVAL_188),
    ._EVAL_189(ibus_int_bus__EVAL_189),
    ._EVAL_190(ibus_int_bus__EVAL_190),
    ._EVAL_191(ibus_int_bus__EVAL_191),
    ._EVAL_192(ibus_int_bus__EVAL_192),
    ._EVAL_193(ibus_int_bus__EVAL_193),
    ._EVAL_194(ibus_int_bus__EVAL_194),
    ._EVAL_195(ibus_int_bus__EVAL_195),
    ._EVAL_196(ibus_int_bus__EVAL_196),
    ._EVAL_197(ibus_int_bus__EVAL_197),
    ._EVAL_198(ibus_int_bus__EVAL_198),
    ._EVAL_199(ibus_int_bus__EVAL_199),
    ._EVAL_200(ibus_int_bus__EVAL_200),
    ._EVAL_201(ibus_int_bus__EVAL_201),
    ._EVAL_202(ibus_int_bus__EVAL_202),
    ._EVAL_203(ibus_int_bus__EVAL_203),
    ._EVAL_204(ibus_int_bus__EVAL_204),
    ._EVAL_205(ibus_int_bus__EVAL_205),
    ._EVAL_206(ibus_int_bus__EVAL_206),
    ._EVAL_207(ibus_int_bus__EVAL_207),
    ._EVAL_208(ibus_int_bus__EVAL_208),
    ._EVAL_209(ibus_int_bus__EVAL_209),
    ._EVAL_210(ibus_int_bus__EVAL_210),
    ._EVAL_211(ibus_int_bus__EVAL_211),
    ._EVAL_212(ibus_int_bus__EVAL_212),
    ._EVAL_213(ibus_int_bus__EVAL_213),
    ._EVAL_214(ibus_int_bus__EVAL_214),
    ._EVAL_215(ibus_int_bus__EVAL_215),
    ._EVAL_216(ibus_int_bus__EVAL_216),
    ._EVAL_217(ibus_int_bus__EVAL_217),
    ._EVAL_218(ibus_int_bus__EVAL_218),
    ._EVAL_219(ibus_int_bus__EVAL_219),
    ._EVAL_220(ibus_int_bus__EVAL_220),
    ._EVAL_221(ibus_int_bus__EVAL_221),
    ._EVAL_222(ibus_int_bus__EVAL_222),
    ._EVAL_223(ibus_int_bus__EVAL_223),
    ._EVAL_224(ibus_int_bus__EVAL_224),
    ._EVAL_225(ibus_int_bus__EVAL_225),
    ._EVAL_226(ibus_int_bus__EVAL_226),
    ._EVAL_227(ibus_int_bus__EVAL_227),
    ._EVAL_228(ibus_int_bus__EVAL_228),
    ._EVAL_229(ibus_int_bus__EVAL_229),
    ._EVAL_230(ibus_int_bus__EVAL_230),
    ._EVAL_231(ibus_int_bus__EVAL_231),
    ._EVAL_232(ibus_int_bus__EVAL_232),
    ._EVAL_233(ibus_int_bus__EVAL_233),
    ._EVAL_234(ibus_int_bus__EVAL_234),
    ._EVAL_235(ibus_int_bus__EVAL_235),
    ._EVAL_236(ibus_int_bus__EVAL_236),
    ._EVAL_237(ibus_int_bus__EVAL_237),
    ._EVAL_238(ibus_int_bus__EVAL_238),
    ._EVAL_239(ibus_int_bus__EVAL_239),
    ._EVAL_240(ibus_int_bus__EVAL_240),
    ._EVAL_241(ibus_int_bus__EVAL_241),
    ._EVAL_242(ibus_int_bus__EVAL_242),
    ._EVAL_243(ibus_int_bus__EVAL_243),
    ._EVAL_244(ibus_int_bus__EVAL_244),
    ._EVAL_245(ibus_int_bus__EVAL_245),
    ._EVAL_246(ibus_int_bus__EVAL_246),
    ._EVAL_247(ibus_int_bus__EVAL_247),
    ._EVAL_248(ibus_int_bus__EVAL_248),
    ._EVAL_249(ibus_int_bus__EVAL_249),
    ._EVAL_250(ibus_int_bus__EVAL_250),
    ._EVAL_251(ibus_int_bus__EVAL_251),
    ._EVAL_252(ibus_int_bus__EVAL_252)
  );
  _EVAL_185 debug_1 (
    ._EVAL(debug_1__EVAL),
    ._EVAL_0(debug_1__EVAL_0),
    ._EVAL_1(debug_1__EVAL_1),
    ._EVAL_2(debug_1__EVAL_2),
    ._EVAL_3(debug_1__EVAL_3),
    ._EVAL_4(debug_1__EVAL_4),
    ._EVAL_5(debug_1__EVAL_5),
    ._EVAL_6(debug_1__EVAL_6),
    ._EVAL_7(debug_1__EVAL_7),
    ._EVAL_8(debug_1__EVAL_8),
    ._EVAL_9(debug_1__EVAL_9),
    ._EVAL_10(debug_1__EVAL_10),
    ._EVAL_11(debug_1__EVAL_11),
    ._EVAL_12(debug_1__EVAL_12),
    ._EVAL_13(debug_1__EVAL_13),
    ._EVAL_14(debug_1__EVAL_14),
    ._EVAL_15(debug_1__EVAL_15),
    ._EVAL_16(debug_1__EVAL_16),
    ._EVAL_17(debug_1__EVAL_17),
    ._EVAL_18(debug_1__EVAL_18),
    ._EVAL_19(debug_1__EVAL_19),
    ._EVAL_20(debug_1__EVAL_20),
    ._EVAL_21(debug_1__EVAL_21),
    ._EVAL_22(debug_1__EVAL_22),
    ._EVAL_23(debug_1__EVAL_23),
    ._EVAL_24(debug_1__EVAL_24),
    ._EVAL_25(debug_1__EVAL_25),
    ._EVAL_26(debug_1__EVAL_26),
    ._EVAL_27(debug_1__EVAL_27),
    ._EVAL_28(debug_1__EVAL_28),
    ._EVAL_29(debug_1__EVAL_29),
    ._EVAL_30(debug_1__EVAL_30),
    ._EVAL_31(debug_1__EVAL_31),
    ._EVAL_32(debug_1__EVAL_32),
    ._EVAL_33(debug_1__EVAL_33),
    ._EVAL_34(debug_1__EVAL_34),
    ._EVAL_35(debug_1__EVAL_35),
    ._EVAL_36(debug_1__EVAL_36),
    ._EVAL_37(debug_1__EVAL_37),
    ._EVAL_38(debug_1__EVAL_38),
    ._EVAL_39(debug_1__EVAL_39),
    ._EVAL_40(debug_1__EVAL_40),
    ._EVAL_41(debug_1__EVAL_41),
    ._EVAL_42(debug_1__EVAL_42),
    ._EVAL_43(debug_1__EVAL_43),
    ._EVAL_44(debug_1__EVAL_44),
    ._EVAL_45(debug_1__EVAL_45)
  );
  _EVAL_193 intsink_1 (
    ._EVAL(intsink_1__EVAL),
    ._EVAL_0(intsink_1__EVAL_0)
  );
  _EVAL_22 subsystem_sbus (
    ._EVAL(subsystem_sbus__EVAL),
    ._EVAL_0(subsystem_sbus__EVAL_0),
    ._EVAL_1(subsystem_sbus__EVAL_1),
    ._EVAL_2(subsystem_sbus__EVAL_2),
    ._EVAL_3(subsystem_sbus__EVAL_3),
    ._EVAL_4(subsystem_sbus__EVAL_4),
    ._EVAL_5(subsystem_sbus__EVAL_5),
    ._EVAL_6(subsystem_sbus__EVAL_6),
    ._EVAL_7(subsystem_sbus__EVAL_7),
    ._EVAL_8(subsystem_sbus__EVAL_8),
    ._EVAL_9(subsystem_sbus__EVAL_9),
    ._EVAL_10(subsystem_sbus__EVAL_10),
    ._EVAL_11(subsystem_sbus__EVAL_11),
    ._EVAL_12(subsystem_sbus__EVAL_12),
    ._EVAL_13(subsystem_sbus__EVAL_13),
    ._EVAL_14(subsystem_sbus__EVAL_14),
    ._EVAL_15(subsystem_sbus__EVAL_15),
    ._EVAL_16(subsystem_sbus__EVAL_16),
    ._EVAL_17(subsystem_sbus__EVAL_17),
    ._EVAL_18(subsystem_sbus__EVAL_18),
    ._EVAL_19(subsystem_sbus__EVAL_19),
    ._EVAL_20(subsystem_sbus__EVAL_20),
    ._EVAL_21(subsystem_sbus__EVAL_21),
    ._EVAL_22(subsystem_sbus__EVAL_22),
    ._EVAL_23(subsystem_sbus__EVAL_23),
    ._EVAL_24(subsystem_sbus__EVAL_24),
    ._EVAL_25(subsystem_sbus__EVAL_25),
    ._EVAL_26(subsystem_sbus__EVAL_26),
    ._EVAL_27(subsystem_sbus__EVAL_27),
    ._EVAL_28(subsystem_sbus__EVAL_28),
    ._EVAL_29(subsystem_sbus__EVAL_29),
    ._EVAL_30(subsystem_sbus__EVAL_30),
    ._EVAL_31(subsystem_sbus__EVAL_31),
    ._EVAL_32(subsystem_sbus__EVAL_32),
    ._EVAL_33(subsystem_sbus__EVAL_33),
    ._EVAL_34(subsystem_sbus__EVAL_34),
    ._EVAL_35(subsystem_sbus__EVAL_35),
    ._EVAL_36(subsystem_sbus__EVAL_36),
    ._EVAL_37(subsystem_sbus__EVAL_37),
    ._EVAL_38(subsystem_sbus__EVAL_38),
    ._EVAL_39(subsystem_sbus__EVAL_39),
    ._EVAL_40(subsystem_sbus__EVAL_40),
    ._EVAL_41(subsystem_sbus__EVAL_41),
    ._EVAL_42(subsystem_sbus__EVAL_42),
    ._EVAL_43(subsystem_sbus__EVAL_43),
    ._EVAL_44(subsystem_sbus__EVAL_44),
    ._EVAL_45(subsystem_sbus__EVAL_45),
    ._EVAL_46(subsystem_sbus__EVAL_46),
    ._EVAL_47(subsystem_sbus__EVAL_47),
    ._EVAL_48(subsystem_sbus__EVAL_48),
    ._EVAL_49(subsystem_sbus__EVAL_49),
    ._EVAL_50(subsystem_sbus__EVAL_50),
    ._EVAL_51(subsystem_sbus__EVAL_51),
    ._EVAL_52(subsystem_sbus__EVAL_52),
    ._EVAL_53(subsystem_sbus__EVAL_53),
    ._EVAL_54(subsystem_sbus__EVAL_54),
    ._EVAL_55(subsystem_sbus__EVAL_55),
    ._EVAL_56(subsystem_sbus__EVAL_56),
    ._EVAL_57(subsystem_sbus__EVAL_57),
    ._EVAL_58(subsystem_sbus__EVAL_58),
    ._EVAL_59(subsystem_sbus__EVAL_59),
    ._EVAL_60(subsystem_sbus__EVAL_60),
    ._EVAL_61(subsystem_sbus__EVAL_61),
    ._EVAL_62(subsystem_sbus__EVAL_62),
    ._EVAL_63(subsystem_sbus__EVAL_63),
    ._EVAL_64(subsystem_sbus__EVAL_64),
    ._EVAL_65(subsystem_sbus__EVAL_65),
    ._EVAL_66(subsystem_sbus__EVAL_66),
    ._EVAL_67(subsystem_sbus__EVAL_67),
    ._EVAL_68(subsystem_sbus__EVAL_68),
    ._EVAL_69(subsystem_sbus__EVAL_69),
    ._EVAL_70(subsystem_sbus__EVAL_70),
    ._EVAL_71(subsystem_sbus__EVAL_71),
    ._EVAL_72(subsystem_sbus__EVAL_72),
    ._EVAL_73(subsystem_sbus__EVAL_73),
    ._EVAL_74(subsystem_sbus__EVAL_74),
    ._EVAL_75(subsystem_sbus__EVAL_75),
    ._EVAL_76(subsystem_sbus__EVAL_76),
    ._EVAL_77(subsystem_sbus__EVAL_77),
    ._EVAL_78(subsystem_sbus__EVAL_78),
    ._EVAL_79(subsystem_sbus__EVAL_79),
    ._EVAL_80(subsystem_sbus__EVAL_80),
    ._EVAL_81(subsystem_sbus__EVAL_81),
    ._EVAL_82(subsystem_sbus__EVAL_82),
    ._EVAL_83(subsystem_sbus__EVAL_83),
    ._EVAL_84(subsystem_sbus__EVAL_84),
    ._EVAL_85(subsystem_sbus__EVAL_85),
    ._EVAL_86(subsystem_sbus__EVAL_86),
    ._EVAL_87(subsystem_sbus__EVAL_87),
    ._EVAL_88(subsystem_sbus__EVAL_88),
    ._EVAL_89(subsystem_sbus__EVAL_89),
    ._EVAL_90(subsystem_sbus__EVAL_90),
    ._EVAL_91(subsystem_sbus__EVAL_91),
    ._EVAL_92(subsystem_sbus__EVAL_92),
    ._EVAL_93(subsystem_sbus__EVAL_93),
    ._EVAL_94(subsystem_sbus__EVAL_94),
    ._EVAL_95(subsystem_sbus__EVAL_95),
    ._EVAL_96(subsystem_sbus__EVAL_96),
    ._EVAL_97(subsystem_sbus__EVAL_97),
    ._EVAL_98(subsystem_sbus__EVAL_98),
    ._EVAL_99(subsystem_sbus__EVAL_99),
    ._EVAL_100(subsystem_sbus__EVAL_100),
    ._EVAL_101(subsystem_sbus__EVAL_101),
    ._EVAL_102(subsystem_sbus__EVAL_102),
    ._EVAL_103(subsystem_sbus__EVAL_103),
    ._EVAL_104(subsystem_sbus__EVAL_104),
    ._EVAL_105(subsystem_sbus__EVAL_105),
    ._EVAL_106(subsystem_sbus__EVAL_106),
    ._EVAL_107(subsystem_sbus__EVAL_107),
    ._EVAL_108(subsystem_sbus__EVAL_108),
    ._EVAL_109(subsystem_sbus__EVAL_109),
    ._EVAL_110(subsystem_sbus__EVAL_110),
    ._EVAL_111(subsystem_sbus__EVAL_111),
    ._EVAL_112(subsystem_sbus__EVAL_112),
    ._EVAL_113(subsystem_sbus__EVAL_113),
    ._EVAL_114(subsystem_sbus__EVAL_114),
    ._EVAL_115(subsystem_sbus__EVAL_115),
    ._EVAL_116(subsystem_sbus__EVAL_116),
    ._EVAL_117(subsystem_sbus__EVAL_117),
    ._EVAL_118(subsystem_sbus__EVAL_118)
  );
  _EVAL_186 xbar_2 (
    ._EVAL(xbar_2__EVAL),
    ._EVAL_0(xbar_2__EVAL_0)
  );
  _EVAL_204 dtm (
    ._EVAL(dtm__EVAL),
    ._EVAL_0(dtm__EVAL_0),
    ._EVAL_1(dtm__EVAL_1),
    ._EVAL_2(dtm__EVAL_2),
    ._EVAL_3(dtm__EVAL_3),
    ._EVAL_4(dtm__EVAL_4),
    ._EVAL_5(dtm__EVAL_5),
    ._EVAL_6(dtm__EVAL_6),
    ._EVAL_7(dtm__EVAL_7),
    ._EVAL_8(dtm__EVAL_8),
    ._EVAL_9(dtm__EVAL_9),
    ._EVAL_10(dtm__EVAL_10),
    ._EVAL_11(dtm__EVAL_11),
    ._EVAL_12(dtm__EVAL_12),
    ._EVAL_13(dtm__EVAL_13),
    ._EVAL_14(dtm__EVAL_14),
    ._EVAL_15(dtm__EVAL_15),
    ._EVAL_16(dtm__EVAL_16)
  );
  SiFive_TLTestIndicator testIndicator (
    .auto_control_xing_in_a_ready(testIndicator_auto_control_xing_in_a_ready),
    .auto_control_xing_in_a_valid(testIndicator_auto_control_xing_in_a_valid),
    .auto_control_xing_in_a_bits_opcode(testIndicator_auto_control_xing_in_a_bits_opcode),
    .auto_control_xing_in_a_bits_param(testIndicator_auto_control_xing_in_a_bits_param),
    .auto_control_xing_in_a_bits_size(testIndicator_auto_control_xing_in_a_bits_size),
    .auto_control_xing_in_a_bits_source(testIndicator_auto_control_xing_in_a_bits_source),
    .auto_control_xing_in_a_bits_address(testIndicator_auto_control_xing_in_a_bits_address),
    .auto_control_xing_in_a_bits_mask(testIndicator_auto_control_xing_in_a_bits_mask),
    .auto_control_xing_in_a_bits_data(testIndicator_auto_control_xing_in_a_bits_data),
    .auto_control_xing_in_a_bits_corrupt(testIndicator_auto_control_xing_in_a_bits_corrupt),
    .auto_control_xing_in_d_ready(testIndicator_auto_control_xing_in_d_ready),
    .auto_control_xing_in_d_valid(testIndicator_auto_control_xing_in_d_valid),
    .auto_control_xing_in_d_bits_opcode(testIndicator_auto_control_xing_in_d_bits_opcode),
    .auto_control_xing_in_d_bits_size(testIndicator_auto_control_xing_in_d_bits_size),
    .auto_control_xing_in_d_bits_source(testIndicator_auto_control_xing_in_d_bits_source),
    .auto_control_xing_in_d_bits_data(testIndicator_auto_control_xing_in_d_bits_data),
    .clock(testIndicator_clock),
    .reset(testIndicator_reset)
  );
  _EVAL_186 xbar_3 (
    ._EVAL(xbar_3__EVAL),
    ._EVAL_0(xbar_3__EVAL_0)
  );
  _EVAL_151 clint (
    ._EVAL(clint__EVAL),
    ._EVAL_0(clint__EVAL_0),
    ._EVAL_1(clint__EVAL_1),
    ._EVAL_2(clint__EVAL_2),
    ._EVAL_3(clint__EVAL_3),
    ._EVAL_4(clint__EVAL_4),
    ._EVAL_5(clint__EVAL_5),
    ._EVAL_6(clint__EVAL_6),
    ._EVAL_7(clint__EVAL_7),
    ._EVAL_8(clint__EVAL_8),
    ._EVAL_9(clint__EVAL_9),
    ._EVAL_10(clint__EVAL_10),
    ._EVAL_11(clint__EVAL_11),
    ._EVAL_12(clint__EVAL_12),
    ._EVAL_13(clint__EVAL_13),
    ._EVAL_14(clint__EVAL_14),
    ._EVAL_15(clint__EVAL_15),
    ._EVAL_16(clint__EVAL_16),
    ._EVAL_17(clint__EVAL_17),
    ._EVAL_18(clint__EVAL_18),
    ._EVAL_19(clint__EVAL_19)
  );
  _EVAL_192 intsource_2 (
    ._EVAL(intsource_2__EVAL),
    ._EVAL_0(intsource_2__EVAL_0),
    ._EVAL_1(intsource_2__EVAL_1),
    ._EVAL_2(intsource_2__EVAL_2),
    ._EVAL_3(intsource_2__EVAL_3),
    ._EVAL_4(intsource_2__EVAL_4),
    ._EVAL_5(intsource_2__EVAL_5),
    ._EVAL_6(intsource_2__EVAL_6),
    ._EVAL_7(intsource_2__EVAL_7),
    ._EVAL_8(intsource_2__EVAL_8),
    ._EVAL_9(intsource_2__EVAL_9),
    ._EVAL_10(intsource_2__EVAL_10),
    ._EVAL_11(intsource_2__EVAL_11),
    ._EVAL_12(intsource_2__EVAL_12),
    ._EVAL_13(intsource_2__EVAL_13),
    ._EVAL_14(intsource_2__EVAL_14),
    ._EVAL_15(intsource_2__EVAL_15),
    ._EVAL_16(intsource_2__EVAL_16),
    ._EVAL_17(intsource_2__EVAL_17),
    ._EVAL_18(intsource_2__EVAL_18),
    ._EVAL_19(intsource_2__EVAL_19),
    ._EVAL_20(intsource_2__EVAL_20),
    ._EVAL_21(intsource_2__EVAL_21),
    ._EVAL_22(intsource_2__EVAL_22),
    ._EVAL_23(intsource_2__EVAL_23),
    ._EVAL_24(intsource_2__EVAL_24),
    ._EVAL_25(intsource_2__EVAL_25),
    ._EVAL_26(intsource_2__EVAL_26),
    ._EVAL_27(intsource_2__EVAL_27),
    ._EVAL_28(intsource_2__EVAL_28),
    ._EVAL_29(intsource_2__EVAL_29),
    ._EVAL_30(intsource_2__EVAL_30)
  );
  _EVAL_193 intsink_4 (
    ._EVAL(intsink_4__EVAL),
    ._EVAL_0(intsink_4__EVAL_0)
  );
  assign plicDomainWrapper__EVAL_24 = _EVAL_437;
  assign ibus_int_bus__EVAL_111 = _EVAL_81;
  assign _EVAL_329 = ibus_int_bus__EVAL_80;
  assign debug_1__EVAL_23 = subsystem_cbus__EVAL;
  assign _EVAL_485 = _EVAL_419;
  assign _EVAL_352 = ibus_int_bus__EVAL_101;
  assign tile_prci_domain__EVAL_6 = intsource_2__EVAL_22;
  assign plicDomainWrapper__EVAL_98 = _EVAL_151;
  assign _EVAL_472 = ibus_int_bus__EVAL_251;
  assign _EVAL_344 = ibus_int_bus__EVAL_48;
  assign ibus_int_bus__EVAL_41 = _EVAL_236;
  assign _EVAL_502 = global_interrupts[41];
  assign _EVAL_386 = _EVAL_421;
  assign tile_prci_domain__EVAL_87 = subsystem_cbus__EVAL_1;
  assign _EVAL_129 = ibus_int_bus__EVAL_240;
  assign _EVAL_68 = _EVAL_85;
  assign intsource__EVAL_4 = clint__EVAL_10;
  assign _EVAL_442 = _EVAL_304;
  assign _EVAL_214 = _EVAL_377;
  assign plicDomainWrapper__EVAL_79 = _EVAL_274;
  assign _EVAL_375 = ibus_int_bus__EVAL_159;
  assign _EVAL_250 = _EVAL_511;
  assign _EVAL_467 = global_interrupts[126];
  assign _EVAL_466 = global_interrupts[16];
  assign plicDomainWrapper__EVAL_34 = _EVAL_227;
  assign _EVAL_349 = subsystem_sbus__EVAL_5;
  assign _EVAL_2 = subsystem_sbus__EVAL_71;
  assign plicDomainWrapper__EVAL_106 = _EVAL_128;
  assign _EVAL_49 = _EVAL_255;
  assign plicDomainWrapper__EVAL_113 = _EVAL_136;
  assign _EVAL_421 = _EVAL_214;
  assign subsystem_cbus__EVAL_107 = tile_prci_domain__EVAL_92;
  assign _EVAL_356 = _EVAL_456;
  assign subsystem_cbus__EVAL_49 = _EVAL_179;
  assign tile_prci_domain__EVAL_55 = subsystem_sbus__EVAL_11;
  assign plicDomainWrapper__EVAL_28 = _EVAL_303;
  assign subsystem_sbus__EVAL_111 = subsystem_fbus__EVAL_18;
  assign _EVAL_347 = global_interrupts[28];
  assign _EVAL_110 = global_interrupts[18];
  assign subsystem_cbus__EVAL_85 = _EVAL_68;
  assign _EVAL_20 = ibus_int_bus__EVAL_128;
  assign subsystem_sbus__EVAL_61 = _EVAL_250;
  assign ibus_int_bus__EVAL_22 = _EVAL_399;
  assign intsource_2__EVAL_11 = local_interrupts_0[12];
  assign _EVAL_35 = _EVAL_359;
  assign subsystem_sbus__EVAL_79 = tile_prci_domain__EVAL_27;
  assign ibus_int_bus__EVAL_92 = _EVAL_116;
  assign _EVAL_243 = ibus_int_bus__EVAL_235;
  assign _EVAL_274 = ibus_int_bus__EVAL_156;
  assign _EVAL_39 = _EVAL_349;
  assign _EVAL_16 = global_interrupts[80];
  assign _EVAL_219 = global_interrupts[86];
  assign _EVAL_300 = ibus_int_bus__EVAL_168;
  assign _EVAL_476 = global_interrupts[40];
  assign _EVAL_42 = ibus_int_bus__EVAL_57;
  assign plicDomainWrapper__EVAL_72 = _EVAL_135;
  assign subsystem_sbus__EVAL_60 = tile_prci_domain__EVAL_38;
  assign plicDomainWrapper__EVAL_104 = _EVAL_412;
  assign _EVAL_60 = ibus_int_bus__EVAL_9;
  assign _EVAL_412 = ibus_int_bus__EVAL_97;
  assign plicDomainWrapper__EVAL_101 = _EVAL_115;
  assign _EVAL_174 = _EVAL_489;
  assign _EVAL_486 = ibus_int_bus__EVAL_228;
  assign _EVAL_202 = _EVAL_326;
  assign tile_prci_domain__EVAL_41 = subsystem_cbus__EVAL_69;
  assign debug_1__EVAL_11 = subsystem_cbus__EVAL_132;
  assign debug_1__EVAL_18 = resetctrl_hartIsInReset_0;
  assign _EVAL_493 = global_interrupts[29];
  assign _EVAL_366 = _EVAL_385;
  assign _EVAL_145 = _EVAL_210;
  assign testIndicator_auto_control_xing_in_a_bits_data = subsystem_cbus__EVAL_0;
  assign subsystem_cbus__EVAL_114 = testIndicator_auto_control_xing_in_d_bits_opcode;
  assign subsystem_cbus__EVAL_119 = testIndicator_auto_control_xing_in_d_bits_data;
  assign _EVAL_396 = _EVAL_429;
  assign subsystem_cbus__EVAL_9 = plicDomainWrapper__EVAL_128;
  assign _EVAL_363 = subsystem_sbus__EVAL_21;
  assign _EVAL_376 = global_interrupts[19];
  assign ibus_int_bus__EVAL_14 = _EVAL_431;
  assign plicDomainWrapper__EVAL_116 = _EVAL_100;
  assign ibus_int_bus__EVAL_211 = _EVAL_36;
  assign tile_prci_domain__EVAL_89 = subsystem_sbus__EVAL_36;
  assign tile_prci_domain__EVAL_93 = intsource_2__EVAL_26;
  assign ibus_int_bus__EVAL_149 = _EVAL_7;
  assign _EVAL_183 = global_interrupts[65];
  assign _EVAL_84 = _EVAL_442;
  assign _EVAL_403 = global_interrupts[11];
  assign tile_prci_domain__EVAL_32 = intsource_2__EVAL_16;
  assign debug_1__EVAL_7 = subsystem_cbus__EVAL_39;
  assign ibus_int_bus__EVAL_230 = _EVAL_401;
  assign tile_prci_domain__EVAL_25 = subsystem_cbus__EVAL_73;
  assign _EVAL_47 = global_interrupts[20];
  assign plicDomainWrapper__EVAL_141 = subsystem_cbus__EVAL_7;
  assign subsystem_cbus__EVAL_23 = tile_prci_domain__EVAL_82;
  assign debug_1__EVAL_9 = subsystem_fbus__EVAL_8;
  assign _EVAL_444 = global_interrupts[21];
  assign _EVAL_345 = global_interrupts[100];
  assign _EVAL_132 = global_interrupts[8];
  assign ibus_int_bus__EVAL_45 = _EVAL_269;
  assign _EVAL_140 = ibus_int_bus__EVAL_208;
  assign plicDomainWrapper__EVAL_7 = _EVAL_140;
  assign tile_prci_domain__EVAL_23 = subsystem_cbus__EVAL_2;
  assign clint__EVAL_5 = subsystem_cbus__EVAL_13;
  assign tile_prci_domain__EVAL_29 = tileHartIdNexusNode__EVAL;
  assign subsystem_fbus__EVAL_43 = front_port_ahb_0_hsel;
  assign tile_prci_domain__EVAL_9 = reset_vector_0;
  assign rtc_sync_chain__EVAL_0 = reset;
  assign subsystem_sbus__EVAL_70 = subsystem_fbus__EVAL_26;
  assign _EVAL_477 = global_interrupts[7];
  assign _EVAL_69 = _EVAL_111;
  assign _EVAL_10 = _EVAL_32;
  assign _EVAL_98 = _EVAL_340;
  assign plicDomainWrapper__EVAL_102 = subsystem_cbus__EVAL_54;
  assign _EVAL_462 = _EVAL_424;
  assign _EVAL_107 = global_interrupts[10];
  assign subsystem_cbus__EVAL_80 = _EVAL_479;
  assign _EVAL_28 = ibus_int_bus__EVAL_115;
  assign _EVAL_113 = subsystem_cbus__EVAL_65;
  assign debug_1__EVAL_38 = subsystem_cbus__EVAL_116;
  assign plicDomainWrapper__EVAL_86 = _EVAL_212;
  assign _EVAL_122 = _EVAL_331;
  assign ibus_int_bus__EVAL_180 = _EVAL_258;
  assign _EVAL_463 = _EVAL_172;
  assign _EVAL_4 = global_interrupts[38];
  assign _EVAL_311 = global_interrupts[102];
  assign _EVAL_302 = _EVAL_402;
  assign tile_prci_domain__EVAL_69 = subsystem_sbus__EVAL_17;
  assign plicDomainWrapper__EVAL_50 = _EVAL_222;
  assign plicDomainWrapper__EVAL_10 = _EVAL_268;
  assign plicDomainWrapper__EVAL_120 = _EVAL_17;
  assign _EVAL_256 = global_interrupts[75];
  assign _EVAL_33 = ibus_int_bus__EVAL_229;
  assign _EVAL_195 = _EVAL_279;
  assign _EVAL_266 = _EVAL_415;
  assign _EVAL_260 = ibus_int_bus__EVAL_25;
  assign tile_prci_domain__EVAL_37 = intsource_2__EVAL_20;
  assign subsystem_cbus__EVAL_56 = _EVAL_474;
  assign plicDomainWrapper__EVAL_135 = _EVAL_77;
  assign plicDomainWrapper__EVAL_127 = _EVAL_123;
  assign _EVAL_380 = _EVAL_361;
  assign _EVAL_215 = subsystem_sbus__EVAL_84;
  assign sys_port_ahb_0_haddr = subsystem_sbus__EVAL_16;
  assign ibus_int_bus__EVAL_127 = _EVAL_381;
  assign ibus_int_bus__EVAL_175 = _EVAL_335;
  assign _EVAL_286 = global_interrupts[120];
  assign _EVAL_101 = subsystem_sbus__EVAL_85;
  assign _EVAL_511 = _EVAL_266;
  assign _EVAL_308 = _EVAL_430;
  assign _EVAL_82 = _EVAL_204;
  assign dtm__EVAL_15 = debug_systemjtag_part_number;
  assign subsystem_sbus__EVAL_7 = tile_prci_domain__EVAL_47;
  assign _EVAL_426 = ibus_int_bus__EVAL_135;
  assign _EVAL_448 = ibus_int_bus__EVAL_17;
  assign _EVAL_369 = _EVAL_478;
  assign _EVAL_437 = ibus_int_bus__EVAL_43;
  assign periph_port_ahb_0_hsize = subsystem_cbus__EVAL_29;
  assign plicDomainWrapper__EVAL_80 = subsystem_cbus__EVAL_88;
  assign _EVAL_207 = ibus_int_bus__EVAL_122;
  assign _EVAL_395 = ibus_int_bus__EVAL_243;
  assign _EVAL_494 = ibus_int_bus__EVAL_35;
  assign _EVAL_201 = ibus_int_bus__EVAL_166;
  assign _EVAL_272 = _EVAL_58;
  assign _EVAL_346 = global_interrupts[53];
  assign plicDomainWrapper__EVAL_107 = _EVAL_353;
  assign _EVAL_206 = ibus_int_bus__EVAL_184;
  assign _EVAL_382 = _EVAL_165;
  assign subsystem_cbus__EVAL_4 = clint__EVAL_16;
  assign subsystem_cbus__EVAL_82 = periph_port_ahb_0_hready;
  assign ibus_int_bus__EVAL_19 = _EVAL_193;
  assign _EVAL_163 = subsystem_cbus__EVAL_43;
  assign dtm__EVAL_2 = debug_systemjtag_reset;
  assign _EVAL_359 = subsystem_cbus__EVAL_84;
  assign plicDomainWrapper__EVAL_38 = subsystem_cbus__EVAL_46;
  assign tile_prci_domain__EVAL_95 = subsystem_sbus__EVAL_43;
  assign tile_prci_domain__EVAL_52 = intsource_2__EVAL_2;
  assign subsystem_cbus__EVAL_15 = periph_port_ahb_0_hresp;
  assign plicDomainWrapper__EVAL_109 = _EVAL_217;
  assign subsystem_fbus__EVAL_25 = subsystem_sbus__EVAL_95;
  assign ibus_int_bus__EVAL_21 = _EVAL_372;
  assign ibus_int_bus__EVAL_107 = _EVAL_124;
  assign _EVAL_150 = ibus_int_bus__EVAL_133;
  assign subsystem_sbus__EVAL_19 = tile_prci_domain__EVAL_42;
  assign _EVAL_425 = ibus_int_bus__EVAL_171;
  assign plicDomainWrapper__EVAL_17 = _EVAL_384;
  assign _EVAL_85 = _EVAL_200;
  assign plicDomainWrapper__EVAL_65 = _EVAL_31;
  assign tile_prci_domain__EVAL_39 = intsource_2__EVAL_17;
  assign _EVAL_387 = _EVAL_510;
  assign _EVAL_373 = global_interrupts[72];
  assign subsystem_cbus__EVAL_34 = tile_prci_domain__EVAL;
  assign clint__EVAL_6 = subsystem_cbus__EVAL_129;
  assign subsystem_sbus__EVAL_18 = _EVAL_397;
  assign _EVAL_301 = global_interrupts[82];
  assign tile_prci_domain__EVAL_7 = subsystem_cbus__EVAL_87;
  assign _EVAL_506 = _EVAL_35;
  assign _EVAL_355 = ~_EVAL_209;
  assign plicDomainWrapper__EVAL_29 = _EVAL_262;
  assign _EVAL_217 = ibus_int_bus__EVAL_141;
  assign _EVAL_351 = _EVAL_153;
  assign subsystem_sbus__EVAL_76 = subsystem_fbus__EVAL_6;
  assign intsource_1__EVAL_2 = plicDomainWrapper__EVAL_126;
  assign _EVAL_310 = subsystem_sbus__EVAL_100;
  assign plicDomainWrapper__EVAL_121 = subsystem_cbus__EVAL_125;
  assign subsystem_cbus__EVAL_60 = testIndicator_auto_control_xing_in_d_bits_size;
  assign plicDomainWrapper__EVAL_73 = _EVAL_168;
  assign plicDomainWrapper__EVAL_66 = _EVAL_471;
  assign _EVAL_504 = global_interrupts[58];
  assign ibus_int_bus__EVAL_250 = _EVAL_114;
  assign ibus_int_bus__EVAL_32 = _EVAL_208;
  assign _EVAL_415 = _EVAL_122;
  assign _EVAL_51 = global_interrupts[68];
  assign _EVAL_294 = _EVAL_451;
  assign plicDomainWrapper__EVAL_76 = _EVAL_395;
  assign _EVAL_56 = ibus_int_bus__EVAL_219;
  assign subsystem_sbus__EVAL_102 = tile_prci_domain__EVAL_45;
  assign _EVAL_389 = ibus_int_bus__EVAL_205;
  assign subsystem_cbus__EVAL_18 = testIndicator_auto_control_xing_in_a_ready;
  assign tile_prci_domain__EVAL_40 = subsystem_cbus__EVAL_97;
  assign _EVAL_26 = _EVAL_453;
  assign _EVAL_8 = _EVAL_410;
  assign plicDomainWrapper__EVAL_6 = _EVAL_189;
  assign ibus_int_bus__EVAL_103 = _EVAL_233;
  assign rtc_sync_chain__EVAL_1 = clock;
  assign subsystem_sbus__EVAL_91 = reset;
  assign periph_port_ahb_0_hwdata = subsystem_cbus__EVAL_14;
  assign _EVAL_185 = ibus_int_bus__EVAL_252;
  assign subsystem_sbus__EVAL_82 = tile_prci_domain__EVAL_97;
  assign subsystem_fbus__EVAL_38 = front_port_ahb_0_htrans;
  assign _EVAL_119 = _EVAL_302;
  assign intsource_2__EVAL_24 = local_interrupts_0[9];
  assign _EVAL_152 = _EVAL_405;
  assign _EVAL_401 = global_interrupts[88];
  assign plicDomainWrapper__EVAL_32 = _EVAL_185;
  assign rtc_sync_chain__EVAL = rtc_toggle;
  assign _EVAL_171 = global_interrupts[26];
  assign _EVAL_166 = _EVAL_95;
  assign plicDomainWrapper__EVAL_103 = _EVAL_391;
  assign plicDomainWrapper__EVAL_33 = _EVAL_327;
  assign _EVAL_508 = subsystem_cbus__EVAL_72;
  assign subsystem_fbus__EVAL_29 = subsystem_sbus__EVAL_30;
  assign subsystem_sbus__EVAL_4 = subsystem_fbus__EVAL_41;
  assign _EVAL_118 = global_interrupts[6];
  assign _EVAL_407 = _EVAL_294;
  assign _EVAL_461 = _EVAL_112;
  assign _EVAL_408 = _EVAL_63;
  assign plicDomainWrapper__EVAL_78 = _EVAL_13;
  assign _EVAL_372 = global_interrupts[30];
  assign sys_port_ahb_0_hwdata = subsystem_sbus__EVAL_86;
  assign intsource_2__EVAL_1 = local_interrupts_0[6];
  assign ibus_int_bus__EVAL_191 = _EVAL_441;
  assign _EVAL_22 = _EVAL_407;
  assign plicDomainWrapper__EVAL_77 = _EVAL_496;
  assign _EVAL_350 = _EVAL_492;
  assign _EVAL_247 = ibus_int_bus__EVAL_124;
  assign tile_prci_domain__EVAL_77 = intsource_1__EVAL;
  assign _EVAL_53 = ibus_int_bus__EVAL_49;
  assign ibus_int_bus__EVAL_202 = _EVAL_155;
  assign plicDomainWrapper__EVAL_3 = subsystem_cbus__EVAL_117;
  assign plicDomainWrapper__EVAL_2 = _EVAL_464;
  assign _EVAL_62 = _EVAL_507;
  assign subsystem_fbus__EVAL_11 = debug_1__EVAL_27;
  assign tile_prci_domain__EVAL_57 = subsystem_sbus__EVAL_40;
  assign plicDomainWrapper__EVAL_57 = _EVAL_436;
  assign subsystem_cbus__EVAL_51 = testIndicator_auto_control_xing_in_d_bits_source;
  assign testIndicator_reset = subsystem_cbus__EVAL_17;
  assign ibus_int_bus__EVAL_198 = _EVAL_183;
  assign _EVAL_40 = global_interrupts[1];
  assign ibus_int_bus__EVAL_93 = _EVAL_458;
  assign _EVAL_488 = _EVAL_121;
  assign ibus_int_bus__EVAL_247 = _EVAL_130;
  assign _EVAL_368 = ibus_int_bus__EVAL_52;
  assign _EVAL_164 = _EVAL_83;
  assign ibus_int_bus__EVAL_126 = _EVAL_16;
  assign plicDomainWrapper__EVAL_54 = _EVAL_88;
  assign _EVAL_96 = _EVAL_174;
  assign subsystem_cbus__EVAL_122 = _EVAL_338;
  assign ibus_int_bus__EVAL_94 = _EVAL_299;
  assign plicDomainWrapper__EVAL_43 = subsystem_cbus__EVAL_81;
  assign _EVAL_322 = global_interrupts[108];
  assign plicDomainWrapper__EVAL_124 = _EVAL_404;
  assign plicDomainWrapper__EVAL_59 = subsystem_cbus__EVAL_66;
  assign dtm__EVAL = debug_1__EVAL_17;
  assign _EVAL_125 = ibus_int_bus__EVAL_36;
  assign _EVAL_189 = ibus_int_bus__EVAL_82;
  assign _EVAL_441 = global_interrupts[104];
  assign _EVAL_204 = _EVAL_94;
  assign clint__EVAL_1 = subsystem_cbus__EVAL_90;
  assign _EVAL_38 = global_interrupts[43];
  assign ibus_int_bus__EVAL_231 = _EVAL_337;
  assign _EVAL_452 = global_interrupts[84];
  assign _EVAL_227 = ibus_int_bus__EVAL_74;
  assign debug_1__EVAL_32 = debug_clock;
  assign ibus_int_bus__EVAL_95 = _EVAL_443;
  assign clint__EVAL_11 = subsystem_cbus__EVAL_77;
  assign ibus_int_bus__EVAL_200 = _EVAL_205;
  assign ibus_int_bus__EVAL_129 = _EVAL_231;
  assign ibus_int_bus__EVAL_227 = _EVAL_169;
  assign dtm__EVAL_11 = debug_systemjtag_jtag_TDI;
  assign _EVAL_27 = _EVAL_14;
  assign subsystem_fbus__EVAL_14 = subsystem_sbus__EVAL_72;
  assign _EVAL_505 = ibus_int_bus__EVAL_70;
  assign _EVAL_19 = _EVAL_319;
  assign ibus_int_bus__EVAL_8 = _EVAL_277;
  assign plicDomainWrapper__EVAL_0 = _EVAL_154;
  assign _EVAL_117 = global_interrupts[56];
  assign ibus_int_bus__EVAL_158 = _EVAL_45;
  assign plicDomainWrapper__EVAL_70 = _EVAL_92;
  assign _EVAL_158 = ibus_int_bus__EVAL_216;
  assign subsystem_sbus__EVAL_63 = tile_prci_domain__EVAL_12;
  assign subsystem_fbus__EVAL_17 = front_port_ahb_0_hburst;
  assign clint__EVAL_12 = _EVAL_161;
  assign _EVAL_283 = ibus_int_bus__EVAL_245;
  assign debug_1__EVAL_1 = debug_systemjtag_jtag_TCK;
  assign subsystem_cbus__EVAL_11 = clint__EVAL_17;
  assign xbar__EVAL_0 = intsink_1__EVAL;
  assign plicDomainWrapper__EVAL_115 = _EVAL_352;
  assign debug_ndreset = debug_1__EVAL_26;
  assign subsystem_fbus__EVAL_36 = subsystem_sbus__EVAL_20;
  assign tile_prci_domain__EVAL_78 = subsystem_sbus__EVAL;
  assign _EVAL_220 = ibus_int_bus__EVAL_177;
  assign _EVAL_509 = global_interrupts[121];
  assign _EVAL_489 = _EVAL_446;
  assign _EVAL_154 = ibus_int_bus__EVAL_96;
  assign _EVAL_46 = _EVAL_485;
  assign dtm__EVAL_6 = debug_systemjtag_jtag_TMS;
  assign _EVAL_88 = ibus_int_bus__EVAL_204;
  assign _EVAL_239 = _EVAL_396;
  assign _EVAL_106 = ibus_int_bus__EVAL_220;
  assign _EVAL_383 = _EVAL_159;
  assign _EVAL_233 = global_interrupts[92];
  assign plicDomainWrapper__EVAL = _EVAL_23;
  assign subsystem_fbus__EVAL_24 = debug_1__EVAL_39;
  assign _EVAL_232 = _EVAL_182;
  assign ibus_int_bus__EVAL_142 = _EVAL_477;
  assign _EVAL_324 = _EVAL_215;
  assign periph_port_ahb_0_hmastlock = 1'h0;
  assign _EVAL_58 = _EVAL_22;
  assign _EVAL_263 = global_interrupts[2];
  assign ibus_int_bus__EVAL_118 = _EVAL_341;
  assign plicDomainWrapper__EVAL_64 = _EVAL_448;
  assign tile_prci_domain__EVAL_102 = subsystem_sbus__EVAL_97;
  assign tile_prci_domain__EVAL_65 = subsystem_sbus__EVAL_74;
  assign _EVAL_399 = global_interrupts[5];
  assign ibus_int_bus__EVAL_234 = _EVAL_93;
  assign tile_prci_domain__EVAL_106 = subsystem_cbus__EVAL_100;
  assign periph_port_ahb_0_htrans = subsystem_cbus__EVAL_106;
  assign _EVAL_456 = _EVAL_152;
  assign tile_prci_domain__EVAL_66 = subsystem_cbus__EVAL_31;
  assign _EVAL_358 = global_interrupts[83];
  assign plicDomainWrapper__EVAL_42 = _EVAL_484;
  assign subsystem_sbus__EVAL_47 = subsystem_fbus__EVAL_46;
  assign _EVAL_258 = global_interrupts[101];
  assign _EVAL_281 = global_interrupts[51];
  assign _EVAL_13 = ibus_int_bus__EVAL_85;
  assign ibus_int_bus__EVAL_174 = _EVAL_330;
  assign ibus_int_bus__EVAL_54 = _EVAL_293;
  assign ibus_int_bus__EVAL_153 = _EVAL_281;
  assign _EVAL_334 = _EVAL_369;
  assign plicDomainWrapper__EVAL_52 = _EVAL_240;
  assign _EVAL_479 = _EVAL_3;
  assign _EVAL_111 = _EVAL_19;
  assign plicDomainWrapper__EVAL_142 = _EVAL_425;
  assign subsystem_fbus__EVAL_20 = debug_1__EVAL_10;
  assign ibus_int_bus__EVAL_0 = _EVAL_379;
  assign _EVAL_155 = global_interrupts[27];
  assign _EVAL_208 = global_interrupts[96];
  assign tile_prci_domain__EVAL_72 = subsystem_sbus__EVAL_94;
  assign subsystem_cbus__EVAL_123 = plicDomainWrapper__EVAL_44;
  assign _EVAL_397 = _EVAL_378;
  assign subsystem_sbus__EVAL_44 = tile_prci_domain__EVAL_56;
  assign _EVAL_178 = _EVAL_414;
  assign plicDomainWrapper__EVAL_63 = _EVAL_15;
  assign _EVAL_438 = global_interrupts[9];
  assign _EVAL_475 = global_interrupts[33];
  assign tile_prci_domain__EVAL_21 = subsystem_sbus__EVAL_1;
  assign clint__EVAL_7 = subsystem_cbus__EVAL_124;
  assign ibus_int_bus__EVAL_23 = _EVAL_134;
  assign _EVAL_31 = ibus_int_bus__EVAL_218;
  assign _EVAL_134 = global_interrupts[95];
  assign debug_systemjtag_jtag_TDO_data = dtm__EVAL_7;
  assign debug_1__EVAL_28 = dtm__EVAL_9;
  assign plicDomainWrapper__EVAL_99 = _EVAL_426;
  assign _EVAL_314 = ibus_int_bus__EVAL_162;
  assign _EVAL_282 = ibus_int_bus__EVAL_31;
  assign _EVAL_416 = global_interrupts[74];
  assign _EVAL_507 = _EVAL_272;
  assign _EVAL_440 = _EVAL_196;
  assign debug_systemjtag_jtag_TDO_driven = dtm__EVAL_3;
  assign ibus_int_bus__EVAL_2 = _EVAL_423;
  assign _EVAL_141 = ibus_int_bus__EVAL_1;
  assign tile_prci_domain__EVAL_64 = intsource_2__EVAL_21;
  assign tile_prci_domain__EVAL_75 = subsystem_sbus__EVAL_83;
  assign plicDomainWrapper__EVAL_14 = _EVAL_317;
  assign tile_prci_domain__EVAL_18 = nmi_0_rnmi_interrupt_vector;
  assign _EVAL_431 = global_interrupts[67];
  assign tile_prci_domain__EVAL_53 = intsource_2__EVAL_23;
  assign _EVAL_337 = global_interrupts[32];
  assign ibus_int_bus__EVAL_114 = _EVAL_191;
  assign _EVAL_254 = ibus_int_bus__EVAL_181;
  assign _EVAL_269 = global_interrupts[81];
  assign ibus_int_bus__EVAL_51 = _EVAL_256;
  assign ibus_int_bus__EVAL_88 = _EVAL_38;
  assign ibus_int_bus__EVAL_113 = _EVAL_286;
  assign _EVAL_251 = ibus_int_bus__EVAL_150;
  assign plicDomainWrapper__EVAL_110 = _EVAL_486;
  assign tile_prci_domain__EVAL_73 = intsource__EVAL;
  assign _EVAL_48 = global_interrupts[61];
  assign ibus_int_bus__EVAL_61 = _EVAL_364;
  assign ibus_int_bus__EVAL_222 = _EVAL_238;
  assign plicDomainWrapper__EVAL_130 = _EVAL_158;
  assign _EVAL_126 = ibus_int_bus__EVAL_117;
  assign subsystem_cbus__EVAL_26 = _EVAL_27;
  assign dtm__EVAL_12 = debug_1__EVAL_6;
  assign _EVAL_480 = ibus_int_bus__EVAL_108;
  assign _EVAL_304 = _EVAL_357;
  assign ibus_int_bus__EVAL_75 = _EVAL_117;
  assign _EVAL_74 = _EVAL_24;
  assign _EVAL_0 = global_interrupts[103];
  assign intsource_2__EVAL_6 = local_interrupts_0[5];
  assign testIndicator_auto_control_xing_in_a_bits_opcode = subsystem_cbus__EVAL_131;
  assign _EVAL_279 = _EVAL_508;
  assign _EVAL_318 = ibus_int_bus__EVAL_242;
  assign _EVAL_285 = ibus_int_bus__EVAL_29;
  assign _EVAL_381 = global_interrupts[0];
  assign dtm__EVAL_14 = debug_systemjtag_version;
  assign subsystem_sbus__EVAL_58 = tile_prci_domain__EVAL_79;
  assign ibus_int_bus__EVAL_157 = _EVAL_34;
  assign ibus_int_bus__EVAL_11 = _EVAL_110;
  assign subsystem_sbus__EVAL_96 = clock;
  assign _EVAL_411 = subsystem_sbus__EVAL_99;
  assign subsystem_sbus__EVAL_73 = subsystem_fbus__EVAL_19;
  assign intsource_2__EVAL_7 = local_interrupts_0[4];
  assign subsystem_sbus__EVAL_55 = tile_prci_domain__EVAL_98;
  assign subsystem_fbus__EVAL_45 = front_port_ahb_0_hwrite;
  assign _EVAL_127 = ibus_int_bus__EVAL_110;
  assign testIndicator_auto_control_xing_in_a_bits_size = subsystem_cbus__EVAL_10;
  assign _EVAL_265 = ibus_int_bus__EVAL_3;
  assign tile_prci_domain__EVAL_8 = subsystem_sbus__EVAL_117;
  assign _EVAL_131 = global_interrupts[89];
  assign clint__EVAL_4 = subsystem_cbus__EVAL_92;
  assign _EVAL_365 = rtc_sync_chain__EVAL_2;
  assign plicDomainWrapper__EVAL_71 = _EVAL_78;
  assign dtm__EVAL_1 = debug_1__EVAL_4;
  assign tile_prci_domain__EVAL_90 = subsystem_sbus__EVAL_33;
  assign ibus_int_bus__EVAL_161 = _EVAL_211;
  assign ibus_int_bus__EVAL_102 = _EVAL_476;
  assign intsource_2__EVAL_14 = local_interrupts_0[14];
  assign _EVAL_325 = global_interrupts[24];
  assign plicDomainWrapper__EVAL_61 = _EVAL_499;
  assign subsystem_cbus__EVAL_133 = _EVAL_186;
  assign _EVAL_228 = _EVAL_113;
  assign _EVAL_212 = ibus_int_bus__EVAL_5;
  assign subsystem_sbus__EVAL_49 = tile_prci_domain__EVAL_88;
  assign _EVAL_32 = subsystem_sbus__EVAL_115;
  assign sys_port_ahb_0_hwrite = subsystem_sbus__EVAL_57;
  assign _EVAL_162 = global_interrupts[99];
  assign subsystem_fbus__EVAL_1 = front_port_ahb_0_hready;
  assign subsystem_sbus__EVAL_3 = subsystem_fbus__EVAL_10;
  assign subsystem_fbus__EVAL_28 = subsystem_sbus__EVAL_46;
  assign ibus_int_bus__EVAL_140 = _EVAL_358;
  assign intsink_4__EVAL_0 = tile_prci_domain__EVAL_28;
  assign _EVAL_11 = global_interrupts[122];
  assign _EVAL_410 = subsystem_cbus__EVAL_115;
  assign intsource_2__EVAL_28 = local_interrupts_0[7];
  assign _EVAL_3 = _EVAL_445;
  assign clint__EVAL_14 = subsystem_cbus__EVAL_41;
  assign tile_prci_domain__EVAL_63 = subsystem_cbus__EVAL_130;
  assign _EVAL_328 = ibus_int_bus__EVAL_71;
  assign _EVAL_391 = ibus_int_bus__EVAL_214;
  assign _EVAL_169 = global_interrupts[111];
  assign intsource_1__EVAL_1 = reset;
  assign _EVAL_65 = ibus_int_bus__EVAL_112;
  assign _EVAL_156 = _EVAL_166;
  assign _EVAL_120 = subsystem_cbus__EVAL_3;
  assign intsource_2__EVAL_25 = local_interrupts_0[0];
  assign _EVAL_191 = global_interrupts[13];
  assign subsystem_sbus__EVAL_109 = tile_prci_domain__EVAL_51;
  assign _EVAL_418 = _EVAL_354;
  assign testIndicator_clock = subsystem_cbus__EVAL_102;
  assign _EVAL_205 = global_interrupts[94];
  assign ibus_int_bus__EVAL_232 = _EVAL_503;
  assign _EVAL_320 = global_interrupts[119];
  assign _EVAL_226 = global_interrupts[70];
  assign ibus_int_bus__EVAL_33 = _EVAL_454;
  assign ibus_int_bus__EVAL_119 = _EVAL_0;
  assign subsystem_cbus__EVAL_24 = tile_prci_domain__EVAL_81;
  assign testIndicator_auto_control_xing_in_a_bits_source = subsystem_cbus__EVAL_21;
  assign subsystem_cbus__EVAL_113 = _EVAL_119;
  assign subsystem_sbus__EVAL_116 = reset;
  assign _EVAL_327 = ibus_int_bus__EVAL_236;
  assign plicDomainWrapper__EVAL_69 = _EVAL_146;
  assign _EVAL_354 = subsystem_cbus__EVAL_38;
  assign plicDomainWrapper__EVAL_49 = _EVAL_127;
  assign _EVAL_89 = ibus_int_bus__EVAL_183;
  assign ibus_int_bus__EVAL_99 = _EVAL_497;
  assign _EVAL_276 = _EVAL_432;
  assign _EVAL_221 = ibus_int_bus__EVAL_6;
  assign ibus_int_bus__EVAL_72 = _EVAL_107;
  assign subsystem_cbus__EVAL_94 = tile_prci_domain__EVAL_15;
  assign subsystem_sbus__EVAL_101 = _EVAL_84;
  assign _EVAL_445 = _EVAL_197;
  assign _EVAL_75 = ibus_int_bus__EVAL_195;
  assign clint__EVAL_13 = subsystem_cbus__EVAL_102;
  assign ibus_int_bus__EVAL_16 = _EVAL_362;
  assign _EVAL_378 = _EVAL_422;
  assign subsystem_cbus__EVAL_83 = tile_prci_domain__EVAL_34;
  assign _EVAL_57 = ibus_int_bus__EVAL_189;
  assign plicDomainWrapper__EVAL_22 = _EVAL_220;
  assign tile_prci_domain__EVAL_4 = intsource_2__EVAL_8;
  assign _EVAL_455 = ibus_int_bus__EVAL_246;
  assign _EVAL_180 = ibus_int_bus__EVAL_221;
  assign subsystem_cbus__EVAL_63 = tile_prci_domain__EVAL_71;
  assign debug_1__EVAL_33 = debug_reset;
  assign _EVAL_138 = ibus_int_bus__EVAL_167;
  assign _EVAL_343 = _EVAL_137;
  assign plicDomainWrapper__EVAL_5 = subsystem_cbus__EVAL_86;
  assign subsystem_fbus__EVAL_3 = subsystem_sbus__EVAL_106;
  assign _EVAL_474 = _EVAL_468;
  assign subsystem_sbus__EVAL_92 = _EVAL_270;
  assign front_port_ahb_0_hreadyout = subsystem_fbus__EVAL_34;
  assign _EVAL_335 = global_interrupts[115];
  assign ibus_int_bus__EVAL_20 = _EVAL_263;
  assign ibus_int_bus__EVAL_77 = _EVAL_444;
  assign _EVAL_54 = ibus_int_bus__EVAL_83;
  assign _EVAL_338 = _EVAL_276;
  assign _EVAL_432 = _EVAL_356;
  assign plicDomainWrapper__EVAL_12 = _EVAL_254;
  assign ibus_int_bus__EVAL_64 = _EVAL_483;
  assign plicDomainWrapper__EVAL_75 = _EVAL_321;
  assign plicDomainWrapper__EVAL_35 = _EVAL_318;
  assign _EVAL_70 = ibus_int_bus__EVAL_55;
  assign subsystem_sbus__EVAL_66 = tile_prci_domain__EVAL_84;
  assign plicDomainWrapper__EVAL_13 = _EVAL_392;
  assign _EVAL_172 = _EVAL_288;
  assign ibus_int_bus__EVAL_210 = _EVAL_490;
  assign tile_prci_domain__EVAL_2 = subsystem_cbus__EVAL_110;
  assign subsystem_sbus__EVAL_78 = tile_prci_domain__EVAL_26;
  assign ibus_int_bus__EVAL_123 = _EVAL_409;
  assign _EVAL_176 = global_interrupts[87];
  assign _EVAL_124 = global_interrupts[37];
  assign subsystem_fbus__EVAL_42 = front_port_ahb_0_hsize;
  assign _EVAL_135 = ibus_int_bus__EVAL_165;
  assign _EVAL_478 = subsystem_sbus__EVAL_89;
  assign debug_1__EVAL_44 = subsystem_cbus__EVAL_33;
  assign testIndicator_auto_control_xing_in_a_bits_mask = subsystem_cbus__EVAL_12;
  assign subsystem_sbus__EVAL_6 = tile_prci_domain__EVAL_35;
  assign subsystem_fbus__EVAL_30 = debug_1__EVAL_21;
  assign testIndicator_auto_control_xing_in_a_bits_param = subsystem_cbus__EVAL_111;
  assign tile_prci_domain__EVAL_61 = intsource__EVAL_2;
  assign dtm__EVAL_10 = debug_1__EVAL_19;
  assign subsystem_sbus__EVAL_81 = tile_prci_domain__EVAL_108;
  assign _EVAL_170 = _EVAL_386;
  assign _EVAL_44 = _EVAL_26;
  assign tile_prci_domain__EVAL_100 = psd_test_clock_enable;
  assign _EVAL_498 = global_interrupts[116];
  assign _EVAL_182 = _EVAL_195;
  assign plicDomainWrapper__EVAL_46 = _EVAL_141;
  assign _EVAL_231 = global_interrupts[85];
  assign ibus_int_bus__EVAL_249 = _EVAL_416;
  assign _EVAL_316 = _EVAL_413;
  assign _EVAL_321 = ibus_int_bus__EVAL_248;
  assign _EVAL_370 = _EVAL_1;
  assign _EVAL_496 = ibus_int_bus__EVAL_226;
  assign subsystem_sbus__EVAL_108 = tile_prci_domain__EVAL_60;
  assign intsource_2__EVAL_5 = local_interrupts_0[11];
  assign subsystem_sbus__EVAL_22 = reset;
  assign _EVAL_295 = ibus_int_bus__EVAL_65;
  assign _EVAL_18 = global_interrupts[93];
  assign ibus_int_bus__EVAL_164 = _EVAL_504;
  assign _EVAL_481 = _EVAL_108;
  assign _EVAL_224 = _EVAL_133;
  assign sys_port_ahb_0_hsize = subsystem_sbus__EVAL_59;
  assign plicDomainWrapper__EVAL_23 = _EVAL_57;
  assign plicDomainWrapper__EVAL_36 = _EVAL_201;
  assign _EVAL_179 = _EVAL_316;
  assign ibus_int_bus__EVAL_116 = _EVAL_132;
  assign _EVAL_249 = _EVAL_367;
  assign _EVAL_108 = _EVAL_178;
  assign _EVAL_240 = ibus_int_bus__EVAL_172;
  assign subsystem_sbus__EVAL_14 = subsystem_fbus__EVAL_35;
  assign _EVAL_78 = ibus_int_bus__EVAL_151;
  assign _EVAL_464 = ibus_int_bus__EVAL_212;
  assign _EVAL_198 = global_interrupts[25];
  assign subsystem_sbus__EVAL_90 = tile_prci_domain__EVAL_17;
  assign _EVAL_353 = ibus_int_bus__EVAL_76;
  assign _EVAL_268 = ibus_int_bus__EVAL_125;
  assign plicDomainWrapper__EVAL_85 = _EVAL_328;
  assign _EVAL_165 = _EVAL_342;
  assign _EVAL_377 = subsystem_sbus__EVAL_62;
  assign _EVAL_398 = _EVAL_82;
  assign subsystem_fbus__EVAL_31 = subsystem_sbus__EVAL_75;
  assign _EVAL_116 = global_interrupts[45];
  assign ibus_int_bus__EVAL_225 = _EVAL_291;
  assign _EVAL_262 = ibus_int_bus__EVAL_138;
  assign _EVAL_271 = global_interrupts[14];
  assign debug_1__EVAL_34 = subsystem_fbus__EVAL_15;
  assign _EVAL_392 = ibus_int_bus__EVAL_136;
  assign _EVAL_261 = global_interrupts[123];
  assign _EVAL_97 = global_interrupts[46];
  assign ibus_int_bus__EVAL_86 = _EVAL_403;
  assign plicDomainWrapper__EVAL_8 = _EVAL_54;
  assign _EVAL_61 = _EVAL_160;
  assign debug_1__EVAL = subsystem_fbus__EVAL_9;
  assign ibus_int_bus__EVAL_144 = _EVAL_90;
  assign _EVAL_288 = _EVAL_8;
  assign _EVAL_55 = ibus_int_bus__EVAL_237;
  assign _EVAL_400 = global_interrupts[117];
  assign subsystem_fbus__EVAL_33 = subsystem_sbus__EVAL_118;
  assign plicDomainWrapper__EVAL_111 = _EVAL_28;
  assign _EVAL_137 = _EVAL_374;
  assign subsystem_fbus__EVAL_32 = front_port_ahb_0_hwdata;
  assign subsystem_cbus__EVAL_16 = clint__EVAL_15;
  assign subsystem_sbus__EVAL_87 = _EVAL_290;
  assign plicDomainWrapper__EVAL_53 = _EVAL_344;
  assign _EVAL_259 = global_interrupts[113];
  assign _EVAL_86 = _EVAL_350;
  assign _EVAL_147 = ibus_int_bus__EVAL_91;
  assign testIndicator_auto_control_xing_in_a_bits_corrupt = subsystem_cbus__EVAL_112;
  assign _EVAL_29 = _EVAL_163;
  assign tile_prci_domain__EVAL_3 = intsource_2__EVAL_12;
  assign subsystem_sbus__EVAL_107 = clock;
  assign _EVAL_148 = _EVAL_324;
  assign _EVAL_453 = subsystem_cbus__EVAL_89;
  assign _EVAL_112 = _EVAL_388;
  assign subsystem_cbus__EVAL_68 = periph_port_ahb_0_hrdata;
  assign _EVAL_446 = _EVAL_99;
  assign sys_port_ahb_0_hburst = subsystem_sbus__EVAL_41;
  assign plicDomainWrapper__EVAL_39 = _EVAL_206;
  assign ibus_int_bus__EVAL_12 = _EVAL_371;
  assign ibus_int_bus__EVAL_209 = _EVAL_400;
  assign subsystem_cbus__EVAL_28 = tile_prci_domain__EVAL_5;
  assign sys_port_ahb_0_hmastlock = 1'h0;
  assign ibus_int_bus__EVAL_7 = _EVAL_105;
  assign dtm__EVAL_8 = debug_systemjtag_mfr_id;
  assign _EVAL_203 = _EVAL_30;
  assign tile_prci_domain__EVAL_59 = subsystem_sbus__EVAL_42;
  assign intsource__EVAL_0 = clint__EVAL_9;
  assign plicDomainWrapper__EVAL_100 = _EVAL_180;
  assign front_port_ahb_0_hresp = subsystem_fbus__EVAL_2;
  assign subsystem_cbus__EVAL_42 = _EVAL_62;
  assign _EVAL_487 = ibus_int_bus__EVAL_176;
  assign _EVAL_142 = ibus_int_bus__EVAL_215;
  assign subsystem_cbus__EVAL_50 = _EVAL_79;
  assign debug_1__EVAL_36 = debug_systemjtag_reset;
  assign plicDomainWrapper__EVAL_137 = _EVAL_143;
  assign _EVAL_420 = global_interrupts[59];
  assign tile_prci_domain__EVAL_67 = subsystem_cbus__EVAL_52;
  assign plicDomainWrapper__EVAL_84 = _EVAL_375;
  assign subsystem_sbus__EVAL_45 = external_source_for_core_0_clock;
  assign _EVAL_197 = _EVAL_273;
  assign _EVAL_413 = _EVAL_461;
  assign subsystem_sbus__EVAL_26 = subsystem_fbus__EVAL_12;
  assign ibus_int_bus__EVAL_66 = _EVAL_103;
  assign _EVAL_319 = _EVAL_29;
  assign plicDomainWrapper__EVAL_96 = _EVAL_285;
  assign tile_prci_domain__EVAL_0 = subsystem_sbus__EVAL_110;
  assign sys_port_ahb_0_htrans = subsystem_sbus__EVAL_38;
  assign _EVAL_153 = _EVAL_380;
  assign _EVAL_471 = ibus_int_bus__EVAL_78;
  assign _EVAL_99 = _EVAL_449;
  assign debug_1__EVAL_40 = subsystem_cbus__EVAL_6;
  assign plicDomainWrapper__EVAL_25 = _EVAL_505;
  assign plicDomainWrapper__EVAL_31 = subsystem_cbus__EVAL_103;
  assign periph_port_ahb_0_haddr = subsystem_cbus__EVAL_105;
  assign subsystem_fbus__EVAL_23 = subsystem_sbus__EVAL_53;
  assign _EVAL_385 = _EVAL_39;
  assign _EVAL_490 = global_interrupts[49];
  assign plicDomainWrapper__EVAL_90 = _EVAL_314;
  assign clint__EVAL_19 = subsystem_cbus__EVAL_71;
  assign tile_prci_domain__EVAL_14 = subsystem_cbus__EVAL_121;
  assign _EVAL_168 = ibus_int_bus__EVAL_44;
  assign plicDomainWrapper__EVAL_56 = _EVAL_225;
  assign ibus_int_bus__EVAL_233 = _EVAL_376;
  assign _EVAL_43 = ibus_int_bus__EVAL_47;
  assign _EVAL_419 = subsystem_sbus__EVAL_56;
  assign _EVAL_307 = _EVAL_418;
  assign tile_prci_domain__EVAL_91 = nmi_0_rnmi_exception_vector;
  assign _EVAL_429 = _EVAL_440;
  assign _EVAL_291 = global_interrupts[76];
  assign _EVAL_121 = subsystem_sbus__EVAL_35;
  assign plicDomainWrapper__EVAL_117 = subsystem_cbus__EVAL_53;
  assign plicDomainWrapper__EVAL_45 = _EVAL_282;
  assign _EVAL_450 = _EVAL_164;
  assign _EVAL_100 = ibus_int_bus__EVAL_244;
  assign _EVAL_298 = _EVAL_382;
  assign subsystem_cbus__EVAL_118 = debug_1__EVAL_16;
  assign clint__EVAL_0 = subsystem_cbus__EVAL_20;
  assign testIndicator_auto_control_xing_in_a_bits_address = subsystem_cbus__EVAL_45;
  assign subsystem_cbus__EVAL_30 = plicDomainWrapper__EVAL_11;
  assign plicDomainWrapper__EVAL_83 = _EVAL_472;
  assign _EVAL_104 = global_interrupts[106];
  assign _EVAL_299 = global_interrupts[34];
  assign _EVAL_167 = _EVAL_120;
  assign ibus_int_bus__EVAL_90 = _EVAL_305;
  assign subsystem_cbus__EVAL_27 = tile_prci_domain__EVAL_19;
  assign subsystem_sbus__EVAL_31 = tile_prci_domain__EVAL_70;
  assign debug_1__EVAL_20 = subsystem_cbus__EVAL_95;
  assign ibus_int_bus__EVAL_28 = _EVAL_176;
  assign _EVAL_253 = _EVAL_46;
  assign _EVAL_128 = ibus_int_bus__EVAL_173;
  assign plicDomainWrapper__EVAL_114 = _EVAL_106;
  assign plicDomainWrapper__EVAL_105 = _EVAL_500;
  assign subsystem_fbus__EVAL_40 = front_port_ahb_0_haddr;
  assign _EVAL_394 = ibus_int_bus__EVAL_178;
  assign tile_prci_domain__EVAL_68 = subsystem_sbus__EVAL_67;
  assign plicDomainWrapper__EVAL_30 = _EVAL_199;
  assign _EVAL_357 = _EVAL_25;
  assign _EVAL_374 = _EVAL_91;
  assign plicDomainWrapper__EVAL_139 = _EVAL_394;
  assign _EVAL_41 = _EVAL_253;
  assign _EVAL_379 = global_interrupts[97];
  assign ibus_int_bus__EVAL_26 = _EVAL_373;
  assign _EVAL_177 = ibus_int_bus__EVAL_143;
  assign plicDomainWrapper__EVAL_51 = _EVAL_221;
  assign subsystem_cbus__EVAL_128 = debug_1__EVAL_3;
  assign plicDomainWrapper__EVAL_112 = _EVAL_129;
  assign xbar_3__EVAL_0 = intsink_4__EVAL;
  assign _EVAL_83 = _EVAL_2;
  assign subsystem_sbus__EVAL_69 = tile_prci_domain__EVAL_16;
  assign intsink_3__EVAL_0 = tile_prci_domain__EVAL_96;
  assign ibus_int_bus__EVAL_146 = _EVAL_406;
  assign _EVAL_303 = ibus_int_bus__EVAL_73;
  assign _EVAL_34 = global_interrupts[22];
  assign plicDomainWrapper__EVAL_60 = _EVAL_284;
  assign _EVAL_184 = global_interrupts[39];
  assign _EVAL_289 = ibus_int_bus__EVAL_84;
  assign intsource__EVAL_3 = clock;
  assign debug_1__EVAL_5 = subsystem_cbus__EVAL_93;
  assign plicDomainWrapper__EVAL_87 = _EVAL_243;
  assign ibus_int_bus__EVAL_155 = _EVAL;
  assign _EVAL_361 = _EVAL_44;
  assign _EVAL_63 = _EVAL_506;
  assign _EVAL_278 = global_interrupts[17];
  assign _EVAL_484 = ibus_int_bus__EVAL_147;
  assign tile_prci_domain__EVAL_36 = nmi_0_rnmi;
  assign tile_prci_domain__EVAL_13 = subsystem_cbus__EVAL_48;
  assign subsystem_sbus__EVAL_52 = tile_prci_domain__EVAL_99;
  assign clint__EVAL = subsystem_cbus__EVAL_22;
  assign intsource_1__EVAL_0 = clock;
  assign ibus_int_bus__EVAL_196 = _EVAL_97;
  assign _EVAL_230 = subsystem_sbus__EVAL_25;
  assign plicDomainWrapper__EVAL_82 = _EVAL_473;
  assign plicDomainWrapper__EVAL_81 = _EVAL_53;
  assign _EVAL_238 = global_interrupts[23];
  assign ibus_int_bus__EVAL_79 = _EVAL_438;
  assign _EVAL_7 = global_interrupts[12];
  assign subsystem_sbus__EVAL_64 = tile_prci_domain__EVAL_20;
  assign _EVAL_500 = ibus_int_bus__EVAL_4;
  assign debug_1__EVAL_42 = debug_dmactiveAck;
  assign tile_prci_domain__EVAL_30 = subsystem_cbus__EVAL_37;
  assign wfi_from_tile_0 = xbar_1__EVAL;
  assign plicDomainWrapper__EVAL_132 = _EVAL_455;
  assign _EVAL_211 = global_interrupts[54];
  assign _EVAL_497 = global_interrupts[78];
  assign plicDomainWrapper__EVAL_125 = _EVAL_247;
  assign plicDomainWrapper__EVAL_133 = _EVAL_60;
  assign _EVAL_297 = global_interrupts[31];
  assign intsource_2__EVAL_19 = local_interrupts_0[2];
  assign ibus_int_bus__EVAL_190 = _EVAL_509;
  assign subsystem_fbus__EVAL_7 = subsystem_sbus__EVAL_114;
  assign subsystem_sbus__EVAL_29 = tile_prci_domain__EVAL_11;
  assign subsystem_sbus__EVAL_93 = subsystem_fbus__EVAL_37;
  assign tile_prci_domain__EVAL_10 = subsystem_sbus__EVAL_32;
  assign tile_prci_domain__EVAL_74 = intsource_2__EVAL;
  assign tile_prci_domain__EVAL_86 = subsystem_cbus__EVAL_101;
  assign plicDomainWrapper__EVAL_122 = _EVAL_332;
  assign _EVAL_234 = global_interrupts[69];
  assign subsystem_cbus__EVAL_76 = _EVAL_202;
  assign plicDomainWrapper__EVAL_58 = _EVAL_300;
  assign _EVAL_451 = subsystem_sbus__EVAL_50;
  assign ibus_int_bus__EVAL_154 = _EVAL_420;
  assign plicDomainWrapper__EVAL_93 = _EVAL_177;
  assign _EVAL_503 = global_interrupts[62];
  assign tile_prci_domain__EVAL_101 = subsystem_cbus__EVAL_79;
  assign subsystem_sbus__EVAL_68 = _EVAL_249;
  assign _EVAL_236 = global_interrupts[109];
  assign ibus_int_bus__EVAL_130 = _EVAL_40;
  assign _EVAL_436 = ibus_int_bus__EVAL_194;
  assign subsystem_cbus__EVAL_104 = debug_1__EVAL_29;
  assign _EVAL_309 = _EVAL_167;
  assign dtm__EVAL_4 = debug_systemjtag_jtag_TCK;
  assign _EVAL_499 = ibus_int_bus__EVAL_13;
  assign subsystem_sbus__EVAL_8 = subsystem_fbus__EVAL_44;
  assign periph_port_ahb_0_hprot = subsystem_cbus__EVAL_127;
  assign subsystem_sbus__EVAL_88 = subsystem_fbus__EVAL_16;
  assign _EVAL_468 = _EVAL_387;
  assign _EVAL_341 = global_interrupts[42];
  assign _EVAL_196 = subsystem_cbus__EVAL_44;
  assign _EVAL_67 = ibus_int_bus__EVAL;
  assign _EVAL_296 = _EVAL_41;
  assign _EVAL_460 = ibus_int_bus__EVAL_239;
  assign subsystem_cbus__EVAL_40 = debug_1__EVAL_14;
  assign _EVAL_284 = ibus_int_bus__EVAL_134;
  assign _EVAL_492 = _EVAL_398;
  assign _EVAL_199 = ibus_int_bus__EVAL_217;
  assign plicDomainWrapper__EVAL_129 = _EVAL_70;
  assign _EVAL_92 = ibus_int_bus__EVAL_27;
  assign _EVAL_81 = global_interrupts[63];
  assign ibus_int_bus__EVAL_187 = _EVAL_475;
  assign cease_from_tile_0 = xbar_2__EVAL;
  assign _EVAL_326 = _EVAL_296;
  assign _EVAL_79 = _EVAL_148;
  assign tile_prci_domain__EVAL_58 = subsystem_cbus__EVAL_108;
  assign plicDomainWrapper__EVAL_20 = _EVAL_71;
  assign intsource_2__EVAL_29 = local_interrupts_0[15];
  assign ibus_int_bus__EVAL_213 = _EVAL_278;
  assign _EVAL_94 = _EVAL_230;
  assign tile_prci_domain__EVAL_104 = subsystem_sbus__EVAL_48;
  assign debug_1__EVAL_0 = dtm__EVAL_0;
  assign plicDomainWrapper__EVAL_62 = _EVAL_245;
  assign _EVAL_193 = global_interrupts[124];
  assign tile_prci_domain__EVAL_24 = intsource_2__EVAL_9;
  assign plicDomainWrapper__EVAL_131 = _EVAL_147;
  assign subsystem_cbus__EVAL_35 = _EVAL_96;
  assign _EVAL_430 = _EVAL_203;
  assign ibus_int_bus__EVAL_163 = _EVAL_311;
  assign _EVAL_30 = _EVAL_194;
  assign subsystem_cbus__EVAL_74 = clint__EVAL_2;
  assign subsystem_cbus__EVAL_5 = tile_prci_domain__EVAL_105;
  assign front_port_ahb_0_hrdata = subsystem_fbus__EVAL_39;
  assign ibus_int_bus__EVAL_185 = _EVAL_322;
  assign plicDomainWrapper__EVAL_68 = _EVAL_138;
  assign ibus_int_bus__EVAL_15 = _EVAL_184;
  assign testIndicator_auto_control_xing_in_a_valid = subsystem_cbus__EVAL_64;
  assign plicDomainWrapper__EVAL_37 = subsystem_cbus__EVAL_91;
  assign debug_dmactive = debug_1__EVAL_43;
  assign debug_1__EVAL_25 = dtm__EVAL_5;
  assign ibus_int_bus__EVAL_50 = _EVAL_248;
  assign _EVAL_280 = _EVAL_309;
  assign _EVAL_105 = global_interrupts[107];
  assign ibus_int_bus__EVAL_87 = _EVAL_297;
  assign _EVAL_146 = ibus_int_bus__EVAL_46;
  assign _EVAL_225 = ibus_int_bus__EVAL_132;
  assign plicDomainWrapper__EVAL_89 = _EVAL_190;
  assign _EVAL_491 = _EVAL_101;
  assign _EVAL_36 = global_interrupts[60];
  assign plicDomainWrapper__EVAL_21 = _EVAL_283;
  assign ibus_int_bus__EVAL_106 = _EVAL_234;
  assign plicDomainWrapper__EVAL_144 = _EVAL_42;
  assign _EVAL_449 = _EVAL_488;
  assign periph_port_ahb_0_hwrite = subsystem_cbus__EVAL_58;
  assign _EVAL_330 = global_interrupts[64];
  assign subsystem_sbus__EVAL_54 = _EVAL_64;
  assign _EVAL_109 = _EVAL_482;
  assign subsystem_sbus__EVAL_37 = sys_port_ahb_0_hrdata;
  assign ibus_int_bus__EVAL_182 = _EVAL_47;
  assign _EVAL_115 = ibus_int_bus__EVAL_68;
  assign tile_prci_domain__EVAL_94 = subsystem_sbus__EVAL_105;
  assign intsink_2__EVAL_0 = tile_prci_domain__EVAL_80;
  assign ibus_int_bus__EVAL_131 = _EVAL_467;
  assign ibus_int_bus__EVAL_63 = _EVAL_144;
  assign _EVAL_424 = _EVAL_12;
  assign _EVAL_264 = global_interrupts[44];
  assign tile_prci_domain__EVAL_44 = intsource_2__EVAL_0;
  assign _EVAL_371 = global_interrupts[79];
  assign plicDomainWrapper__EVAL_97 = _EVAL_75;
  assign _EVAL_332 = ibus_int_bus__EVAL_193;
  assign _EVAL_14 = _EVAL_481;
  assign _EVAL_342 = _EVAL_280;
  assign ibus_int_bus__EVAL_170 = _EVAL_271;
  assign plicDomainWrapper__EVAL_55 = _EVAL_295;
  assign subsystem_sbus__EVAL_24 = clock;
  assign plicDomainWrapper__EVAL_67 = _EVAL_267;
  assign _EVAL_181 = global_interrupts[90];
  assign ibus_int_bus__EVAL_186 = _EVAL_48;
  assign tile_prci_domain__EVAL_49 = subsystem_cbus__EVAL_57;
  assign tile_prci_domain__EVAL_43 = intsource_2__EVAL_10;
  assign ibus_int_bus__EVAL_160 = _EVAL_118;
  assign ibus_int_bus__EVAL_37 = _EVAL_320;
  assign tile_prci_domain__EVAL_48 = subsystem_sbus__EVAL_80;
  assign subsystem_cbus__EVAL_96 = tile_prci_domain__EVAL_22;
  assign plicDomainWrapper__EVAL_47 = _EVAL_265;
  assign _EVAL_248 = global_interrupts[125];
  assign xbar_1__EVAL_0 = intsink_2__EVAL;
  assign plicDomainWrapper__EVAL_138 = _EVAL_65;
  assign _EVAL_290 = _EVAL_351;
  assign _EVAL_384 = ibus_int_bus__EVAL_206;
  assign _EVAL_186 = _EVAL_334;
  assign subsystem_fbus__EVAL_21 = front_port_ahb_0_hprot;
  assign intsink_1__EVAL_0 = tile_prci_domain__EVAL_46;
  assign plicDomainWrapper__EVAL_95 = _EVAL_55;
  assign _EVAL_469 = _EVAL_365 & _EVAL_355;
  assign ibus_int_bus__EVAL_89 = _EVAL_261;
  assign _EVAL_133 = _EVAL_308;
  assign subsystem_sbus__EVAL_103 = sys_port_ahb_0_hresp;
  assign ibus_int_bus__EVAL_120 = _EVAL_4;
  assign tile_prci_domain__EVAL_83 = subsystem_sbus__EVAL_2;
  assign _EVAL = global_interrupts[15];
  assign _EVAL_510 = _EVAL_156;
  assign subsystem_sbus__EVAL_9 = _EVAL_145;
  assign subsystem_cbus__EVAL_62 = clint__EVAL_3;
  assign ibus_int_bus__EVAL_100 = _EVAL_466;
  assign sys_port_ahb_0_hprot = subsystem_sbus__EVAL_28;
  assign subsystem_cbus__EVAL_120 = testIndicator_auto_control_xing_in_d_valid;
  assign tile_prci_domain__EVAL_85 = intsource_2__EVAL_13;
  assign subsystem_sbus__EVAL_104 = tile_prci_domain__EVAL_50;
  assign _EVAL_364 = global_interrupts[52];
  assign subsystem_cbus__EVAL_75 = _EVAL_465;
  assign debug_1__EVAL_15 = subsystem_cbus__EVAL_25;
  assign intsource_2__EVAL_4 = local_interrupts_0[8];
  assign ibus_int_bus__EVAL_34 = _EVAL_452;
  assign plicDomainWrapper__EVAL_74 = _EVAL_56;
  assign ibus_int_bus__EVAL_152 = _EVAL_313;
  assign _EVAL_130 = global_interrupts[73];
  assign intsource_2__EVAL_27 = local_interrupts_0[13];
  assign debug_1__EVAL_2 = subsystem_cbus__EVAL_78;
  assign _EVAL_144 = global_interrupts[77];
  assign _EVAL_458 = global_interrupts[98];
  assign _EVAL_443 = global_interrupts[110];
  assign _EVAL_305 = global_interrupts[3];
  assign _EVAL_95 = _EVAL_310;
  assign xbar_2__EVAL_0 = intsink_3__EVAL;
  assign _EVAL_362 = global_interrupts[48];
  assign _EVAL_313 = global_interrupts[114];
  assign _EVAL_473 = ibus_int_bus__EVAL_24;
  assign subsystem_fbus__EVAL_13 = subsystem_sbus__EVAL_39;
  assign _EVAL_245 = ibus_int_bus__EVAL_60;
  assign plicDomainWrapper__EVAL_15 = _EVAL_43;
  assign subsystem_fbus__EVAL_5 = subsystem_sbus__EVAL_65;
  assign _EVAL_423 = global_interrupts[91];
  assign _EVAL_160 = _EVAL_408;
  assign tile_prci_domain__EVAL_103 = subsystem_sbus__EVAL_77;
  assign plicDomainWrapper__EVAL_1 = _EVAL_260;
  assign ibus_int_bus__EVAL_69 = _EVAL_259;
  assign _EVAL_123 = ibus_int_bus__EVAL_10;
  assign subsystem_sbus__EVAL_51 = tile_prci_domain__EVAL_54;
  assign subsystem_sbus__EVAL_23 = tile_prci_domain__EVAL_76;
  assign ibus_int_bus__EVAL_201 = _EVAL_325;
  assign subsystem_sbus__EVAL_10 = _EVAL_298;
  assign debug_1__EVAL_35 = subsystem_cbus__EVAL_8;
  assign intsource_2__EVAL_3 = local_interrupts_0[10];
  assign subsystem_cbus__EVAL_126 = clint__EVAL_8;
  assign _EVAL_23 = ibus_int_bus__EVAL_109;
  assign plicDomainWrapper__EVAL_88 = _EVAL_150;
  assign _EVAL_194 = subsystem_cbus__EVAL_109;
  assign _EVAL_159 = subsystem_sbus__EVAL_34;
  assign _EVAL_465 = _EVAL_393;
  assign intsource_2__EVAL_18 = local_interrupts_0[1];
  assign periph_port_ahb_0_hburst = 3'h0;
  assign _EVAL_200 = _EVAL_188;
  assign plicDomainWrapper__EVAL_27 = _EVAL_251;
  assign clint__EVAL_18 = subsystem_cbus__EVAL_17;
  assign _EVAL_270 = _EVAL_61;
  assign ibus_int_bus__EVAL_137 = _EVAL_502;
  assign _EVAL_406 = global_interrupts[105];
  assign subsystem_sbus__EVAL_13 = external_source_for_core_0_reset;
  assign subsystem_cbus__EVAL_32 = plicDomainWrapper__EVAL_140;
  assign intsource_2__EVAL_30 = local_interrupts_0[3];
  assign ibus_int_bus__EVAL_42 = _EVAL_162;
  assign testIndicator_auto_control_xing_in_d_ready = subsystem_cbus__EVAL_47;
  assign ibus_int_bus__EVAL_104 = _EVAL_493;
  assign _EVAL_188 = _EVAL_98;
  assign subsystem_cbus__EVAL_70 = plicDomainWrapper__EVAL_108;
  assign _EVAL_277 = global_interrupts[57];
  assign subsystem_sbus__EVAL_12 = subsystem_fbus__EVAL_22;
  assign _EVAL_222 = ibus_int_bus__EVAL_148;
  assign _EVAL_15 = ibus_int_bus__EVAL_145;
  assign _EVAL_90 = global_interrupts[4];
  assign _EVAL_388 = _EVAL_287;
  assign plicDomainWrapper__EVAL_16 = _EVAL_33;
  assign ibus_int_bus__EVAL_241 = _EVAL_219;
  assign _EVAL_273 = _EVAL_434;
  assign ibus_int_bus__EVAL_67 = _EVAL_181;
  assign subsystem_sbus__EVAL_27 = subsystem_fbus__EVAL_47;
  assign _EVAL_17 = ibus_int_bus__EVAL_53;
  assign _EVAL_405 = _EVAL_363;
  assign _EVAL_434 = _EVAL_491;
  assign _EVAL_422 = _EVAL_463;
  assign subsystem_cbus__EVAL_67 = debug_1__EVAL_24;
  assign plicDomainWrapper__EVAL_118 = _EVAL_207;
  assign subsystem_sbus__EVAL_0 = _EVAL_462;
  assign ibus_int_bus__EVAL_39 = _EVAL_131;
  assign plicDomainWrapper__EVAL_92 = _EVAL_480;
  assign plicDomainWrapper__EVAL_40 = _EVAL_218;
  assign ibus_int_bus__EVAL_223 = _EVAL_198;
  assign _EVAL_91 = _EVAL_383;
  assign _EVAL_12 = _EVAL_232;
  assign _EVAL_143 = ibus_int_bus__EVAL_105;
  assign _EVAL_103 = global_interrupts[35];
  assign ibus_int_bus__EVAL_18 = _EVAL_347;
  assign _EVAL_1 = _EVAL_366;
  assign ibus_int_bus__EVAL_38 = _EVAL_104;
  assign ibus_int_bus__EVAL_238 = _EVAL_226;
  assign _EVAL_483 = global_interrupts[55];
  assign ibus_int_bus__EVAL_81 = _EVAL_345;
  assign debug_1__EVAL_41 = dtm__EVAL_16;
  assign tile_prci_domain__EVAL_107 = intsource_2__EVAL_15;
  assign subsystem_sbus__EVAL_98 = tile_prci_domain__EVAL_31;
  assign plicDomainWrapper__EVAL_26 = _EVAL_126;
  assign tile_prci_domain__EVAL_1 = debug_1__EVAL_30;
  assign _EVAL_255 = _EVAL_170;
  assign _EVAL_190 = ibus_int_bus__EVAL_62;
  assign _EVAL_151 = ibus_int_bus__EVAL_207;
  assign _EVAL_59 = _EVAL_450;
  assign _EVAL_367 = _EVAL_192;
  assign subsystem_cbus__EVAL_36 = _EVAL_86;
  assign _EVAL_331 = _EVAL_228;
  assign _EVAL_45 = global_interrupts[47];
  assign _EVAL_77 = ibus_int_bus__EVAL_203;
  assign ibus_int_bus__EVAL_199 = _EVAL_498;
  assign subsystem_sbus__EVAL_15 = tile_prci_domain__EVAL_33;
  assign subsystem_cbus__EVAL_98 = tile_prci_domain__EVAL_62;
  assign _EVAL_5 = global_interrupts[36];
  assign plicDomainWrapper__EVAL_119 = _EVAL_20;
  assign _EVAL_267 = ibus_int_bus__EVAL_179;
  assign plicDomainWrapper__EVAL_91 = _EVAL_368;
  assign intsource__EVAL_1 = reset;
  assign _EVAL_52 = _EVAL_49;
  assign _EVAL_340 = _EVAL_10;
  assign plicDomainWrapper__EVAL_4 = _EVAL_389;
  assign _EVAL_25 = _EVAL_307;
  assign _EVAL_409 = global_interrupts[71];
  assign plicDomainWrapper__EVAL_136 = _EVAL_142;
  assign _EVAL_454 = global_interrupts[50];
  assign ibus_int_bus__EVAL_56 = _EVAL_11;
  assign plicDomainWrapper__EVAL_41 = _EVAL_494;
  assign _EVAL_71 = ibus_int_bus__EVAL_169;
  assign plicDomainWrapper__EVAL_134 = _EVAL_460;
  assign subsystem_sbus__EVAL_113 = sys_port_ahb_0_hready;
  assign _EVAL_393 = _EVAL_370;
  assign subsystem_fbus__EVAL_4 = debug_1__EVAL_13;
  assign subsystem_cbus__EVAL_19 = debug_1__EVAL_31;
  assign debug_1__EVAL_12 = subsystem_fbus__EVAL;
  assign _EVAL_192 = _EVAL_239;
  assign plicDomainWrapper__EVAL_123 = _EVAL_329;
  assign plicDomainWrapper__EVAL_9 = _EVAL_67;
  assign ibus_int_bus__EVAL_30 = _EVAL_301;
  assign _EVAL_404 = ibus_int_bus__EVAL_139;
  assign plicDomainWrapper__EVAL_94 = _EVAL_89;
  assign _EVAL_218 = ibus_int_bus__EVAL_188;
  assign ibus_int_bus__EVAL_40 = _EVAL_264;
  assign ibus_int_bus__EVAL_121 = _EVAL_5;
  assign subsystem_fbus__EVAL_27 = debug_1__EVAL_8;
  assign _EVAL_136 = ibus_int_bus__EVAL_224;
  assign ibus_int_bus__EVAL_197 = _EVAL_51;
  assign plicDomainWrapper__EVAL_18 = _EVAL_289;
  assign debug_from_tile_0 = xbar_3__EVAL;
  assign _EVAL_317 = ibus_int_bus__EVAL_192;
  assign subsystem_cbus__EVAL_55 = _EVAL_74;
  assign _EVAL_114 = global_interrupts[118];
  assign debug_1__EVAL_45 = dtm__EVAL_13;
  assign ibus_int_bus__EVAL_59 = _EVAL_346;
  assign debug_1__EVAL_37 = subsystem_cbus__EVAL_99;
  assign _EVAL_293 = global_interrupts[66];
  assign _EVAL_414 = _EVAL_109;
  assign _EVAL_64 = _EVAL_224;
  assign _EVAL_93 = global_interrupts[112];
  assign ibus_int_bus__EVAL_98 = _EVAL_171;
  assign _EVAL_24 = _EVAL_343;
  assign halt_from_tile_0 = xbar__EVAL;
  assign _EVAL_210 = _EVAL_69;
  assign plicDomainWrapper__EVAL_48 = _EVAL_487;
  assign _EVAL_287 = _EVAL_411;
  assign ibus_int_bus__EVAL_58 = _EVAL_18;
  assign plicDomainWrapper__EVAL_143 = _EVAL_125;
  assign _EVAL_402 = _EVAL_59;
  assign _EVAL_482 = subsystem_sbus__EVAL_112;
  assign debug_1__EVAL_22 = subsystem_fbus__EVAL_0;
  assign subsystem_cbus__EVAL_61 = _EVAL_52;
  assign subsystem_cbus__EVAL_59 = plicDomainWrapper__EVAL_19;
  always @(posedge clock) begin
    if (reset) begin
      _EVAL_161 <= 1'h0;
    end else begin
      _EVAL_161 <= _EVAL_469;
    end
    if (reset) begin
      _EVAL_209 <= 1'h0;
    end else begin
      _EVAL_209 <= _EVAL_365;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_161 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_209 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
