//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_127(
  output        _EVAL,
  output [1:0]  _EVAL_0,
  output [31:0] _EVAL_1,
  output        _EVAL_2,
  output        _EVAL_3,
  output [31:0] _EVAL_4,
  input         _EVAL_5,
  output        _EVAL_6,
  output        _EVAL_7,
  output        _EVAL_8,
  output        _EVAL_9,
  input         _EVAL_10,
  output        _EVAL_11,
  output        _EVAL_12,
  output [1:0]  _EVAL_13,
  output [1:0]  _EVAL_14,
  output [31:0] _EVAL_15,
  output        _EVAL_16,
  output        _EVAL_17,
  input         _EVAL_18,
  output        _EVAL_19,
  input         _EVAL_20,
  input         _EVAL_21,
  output        _EVAL_22,
  input         _EVAL_23,
  output [1:0]  _EVAL_24,
  output        _EVAL_25,
  output [1:0]  _EVAL_26,
  input  [31:0] _EVAL_27,
  input  [31:0] _EVAL_28,
  output        _EVAL_29,
  output        _EVAL_30,
  output [1:0]  _EVAL_31,
  output        _EVAL_32,
  output        _EVAL_33,
  output [31:0] _EVAL_34,
  output        _EVAL_35,
  output        _EVAL_36,
  output        _EVAL_37,
  output        _EVAL_38,
  output        _EVAL_39,
  output [29:0] _EVAL_40,
  input         _EVAL_41,
  output [29:0] _EVAL_42,
  output [1:0]  _EVAL_43,
  output [31:0] _EVAL_44,
  input         _EVAL_45,
  output [31:0] _EVAL_46,
  output        _EVAL_47,
  output        _EVAL_48,
  input         _EVAL_49,
  input  [31:0] _EVAL_50,
  input         _EVAL_51,
  output [31:0] _EVAL_52,
  output        _EVAL_53,
  output        _EVAL_54,
  output        _EVAL_55,
  output [31:0] _EVAL_56,
  input         _EVAL_57,
  output        _EVAL_58,
  output        _EVAL_59,
  output [1:0]  _EVAL_60,
  output        _EVAL_61,
  input         _EVAL_62,
  input         _EVAL_63,
  output [31:0] _EVAL_64,
  output        _EVAL_65,
  input         _EVAL_66,
  output [1:0]  _EVAL_67,
  output        _EVAL_68,
  output        _EVAL_69,
  output [31:0] _EVAL_70,
  output [31:0] _EVAL_71,
  output        _EVAL_72,
  input  [31:0] _EVAL_73,
  output        _EVAL_74,
  output        _EVAL_75,
  output        _EVAL_76,
  output        _EVAL_77,
  output        _EVAL_78,
  output        _EVAL_79,
  output        _EVAL_80,
  output        _EVAL_81,
  output [7:0]  _EVAL_82,
  input         _EVAL_83,
  input         _EVAL_84,
  input         _EVAL_85,
  input         _EVAL_86,
  output [29:0] _EVAL_87,
  input         _EVAL_88,
  output [1:0]  _EVAL_89,
  input         _EVAL_90,
  output        _EVAL_91,
  output [1:0]  _EVAL_92,
  output        _EVAL_93,
  output [31:0] _EVAL_94,
  output        _EVAL_95,
  output        _EVAL_96,
  output [31:0] _EVAL_97,
  output        _EVAL_98,
  output        _EVAL_99,
  output [1:0]  _EVAL_100,
  input  [31:0] _EVAL_101,
  input         _EVAL_102,
  output [31:0] _EVAL_103,
  output [31:0] _EVAL_104,
  output [29:0] _EVAL_105,
  output        _EVAL_106,
  output        _EVAL_107,
  output [2:0]  _EVAL_108,
  output        _EVAL_109,
  output        _EVAL_110,
  output        _EVAL_111,
  output        _EVAL_112,
  input  [11:0] _EVAL_113,
  output        _EVAL_114,
  output        _EVAL_115,
  output [31:0] _EVAL_116,
  output        _EVAL_117,
  output [31:0] _EVAL_118,
  output        _EVAL_119,
  input         _EVAL_120,
  input         _EVAL_121,
  output [26:0] _EVAL_122,
  output [1:0]  _EVAL_123,
  output [31:0] _EVAL_124,
  output [1:0]  _EVAL_125,
  input         _EVAL_126,
  output        _EVAL_127,
  output        _EVAL_128,
  output        _EVAL_129,
  input  [31:0] _EVAL_130,
  output        _EVAL_131,
  output        _EVAL_132,
  input  [31:0] _EVAL_133,
  input  [2:0]  _EVAL_134,
  input         _EVAL_135,
  output        _EVAL_136,
  output        _EVAL_137,
  output        _EVAL_138,
  output [1:0]  _EVAL_139,
  output [31:0] _EVAL_140,
  input         _EVAL_141,
  output        _EVAL_142,
  output [1:0]  _EVAL_143,
  output [29:0] _EVAL_144,
  output [31:0] _EVAL_145,
  output        _EVAL_146,
  output        _EVAL_147,
  output [29:0] _EVAL_148,
  output        _EVAL_149,
  output        _EVAL_150,
  input  [11:0] _EVAL_151,
  output        _EVAL_152,
  input         _EVAL_153,
  output        _EVAL_154,
  output        _EVAL_155,
  output        _EVAL_156,
  output        _EVAL_157,
  output [31:0] _EVAL_158,
  output        _EVAL_159,
  output [29:0] _EVAL_160,
  output [31:0] _EVAL_161,
  output [1:0]  _EVAL_162,
  output [29:0] _EVAL_163,
  output        _EVAL_164,
  output [31:0] _EVAL_165,
  input         _EVAL_166,
  input         _EVAL_167,
  output        _EVAL_168,
  output [31:0] _EVAL_169,
  output        _EVAL_170,
  output [1:0]  _EVAL_171,
  output        _EVAL_172,
  output        _EVAL_173,
  output        _EVAL_174,
  output        _EVAL_175,
  output [1:0]  _EVAL_176,
  output [1:0]  _EVAL_177,
  output        _EVAL_178,
  output        _EVAL_179,
  output        _EVAL_180,
  output        _EVAL_181,
  output        _EVAL_182,
  output        _EVAL_183,
  output        _EVAL_184,
  output        _EVAL_185,
  output        _EVAL_186
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [63:0] _RAND_163;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_194;
  wire [33:0] _EVAL_195;
  wire  _EVAL_196;
  wire [31:0] _EVAL_197;
  wire [102:0] _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_204;
  wire [31:0] _EVAL_205;
  wire [32:0] _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire [102:0] _EVAL_210;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire [4:0] _EVAL_216;
  wire [102:0] _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_221;
  wire [30:0] _EVAL_222;
  wire [31:0] _EVAL_223;
  wire  _EVAL_225;
  reg [29:0] _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_230;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire [6:0] _EVAL_234;
  wire [31:0] _EVAL_235;
  wire  _EVAL_236;
  reg [1:0] _EVAL_237;
  wire [7:0] _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_242;
  wire [30:0] _EVAL_243;
  wire  _EVAL_244;
  reg  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_248;
  wire [31:0] _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire [4:0] _EVAL_253;
  wire [31:0] _EVAL_254;
  wire [39:0] _EVAL_256;
  wire  _EVAL_258;
  wire  _EVAL_260;
  wire [31:0] _EVAL_262;
  wire [102:0] _EVAL_265;
  wire  _EVAL_267;
  wire [31:0] _EVAL_268;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_277;
  wire  _EVAL_279;
  reg [31:0] _EVAL_280;
  wire  _EVAL_281;
  reg  _EVAL_282;
  wire [4:0] _EVAL_283;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire [39:0] _EVAL_289;
  wire  _EVAL_291;
  wire [31:0] _EVAL_293;
  wire  _EVAL_295;
  wire  _EVAL_297;
  wire [31:0] _EVAL_298;
  wire  _EVAL_299;
  wire [6:0] _EVAL_300;
  wire [63:0] _EVAL_302;
  wire  _EVAL_304;
  wire [31:0] _EVAL_305;
  wire [1:0] _EVAL_306;
  wire [4:0] _EVAL_307;
  wire [7:0] _EVAL_308;
  wire  _EVAL_311;
  reg [1:0] _EVAL_312;
  reg  _EVAL_313;
  wire  _EVAL_314;
  wire [31:0] _EVAL_315;
  wire  _EVAL_316;
  wire [102:0] _EVAL_317;
  wire [102:0] _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_320;
  wire [1:0] _EVAL_321;
  wire [102:0] _EVAL_322;
  wire  _EVAL_323;
  wire  _EVAL_324;
  wire [31:0] _EVAL_325;
  wire  _EVAL_326;
  wire  _EVAL_327;
  wire [1:0] _EVAL_329;
  wire [31:0] _EVAL_330;
  wire  _EVAL_332;
  wire  _EVAL_333;
  wire  _EVAL_334;
  wire [4:0] _EVAL_336;
  wire  _EVAL_337;
  wire  _EVAL_342;
  wire  _EVAL_343;
  wire  _EVAL_345;
  wire  _EVAL_346;
  wire  _EVAL_348;
  wire  _EVAL_349;
  wire  _EVAL_350;
  wire  _EVAL_351;
  wire  _EVAL_353;
  wire  _EVAL_354;
  wire  _EVAL_355;
  wire  _EVAL_356;
  wire  _EVAL_357;
  wire  _EVAL_358;
  reg [29:0] _EVAL_359;
  wire  _EVAL_360;
  wire  _EVAL_361;
  wire [6:0] _EVAL_362;
  wire [31:0] _EVAL_363;
  wire [31:0] _EVAL_364;
  reg [1:0] _EVAL_365;
  reg  _EVAL_366;
  wire [102:0] _EVAL_367;
  wire  _EVAL_368;
  wire  _EVAL_369;
  reg  _EVAL_370;
  wire  _EVAL_372;
  wire  _EVAL_373;
  wire [31:0] _EVAL_375;
  wire [31:0] _EVAL_377;
  wire [4:0] _EVAL_378;
  wire [2:0] _EVAL_379;
  wire  _EVAL_380;
  wire [31:0] _EVAL_381;
  wire  _EVAL_382;
  wire [30:0] _EVAL_384;
  reg [31:0] _EVAL_385;
  wire  _EVAL_386;
  reg [31:0] _EVAL_387;
  wire  _EVAL_388;
  wire  _EVAL_389;
  wire  _EVAL_390;
  wire [1:0] _EVAL_391;
  wire [1:0] _EVAL_392;
  wire  _EVAL_394;
  reg [1:0] _EVAL_395;
  wire  _EVAL_397;
  wire  _EVAL_398;
  wire [1:0] _EVAL_400;
  wire [29:0] _EVAL_401;
  wire [31:0] _EVAL_402;
  wire [29:0] _EVAL_403;
  wire  _EVAL_404;
  wire [30:0] _EVAL_405;
  wire  _EVAL_407;
  wire [30:0] _EVAL_408;
  wire  _EVAL_410;
  wire  _EVAL_412;
  wire [31:0] _EVAL_413;
  wire  _EVAL_414;
  reg  _EVAL_417;
  wire [57:0] _EVAL_418;
  wire  _EVAL_419;
  wire  _EVAL_420;
  wire  _EVAL_424;
  wire  _EVAL_426;
  wire [1:0] _EVAL_427;
  wire  _EVAL_428;
  wire [31:0] _EVAL_429;
  wire [30:0] _EVAL_430;
  wire  _EVAL_431;
  wire  _EVAL_432;
  wire  _EVAL_434;
  wire  _EVAL_436;
  wire [57:0] _EVAL_437;
  wire [30:0] _EVAL_438;
  wire [31:0] _EVAL_439;
  wire [31:0] _EVAL_440;
  wire [31:0] _EVAL_441;
  wire [15:0] _EVAL_443;
  wire  _EVAL_444;
  wire  _EVAL_445;
  wire  _EVAL_446;
  wire [4:0] _EVAL_447;
  wire  _EVAL_448;
  wire  _EVAL_450;
  wire [31:0] _EVAL_451;
  wire  _EVAL_452;
  reg  _EVAL_454;
  wire  _EVAL_456;
  wire  _EVAL_459;
  reg  _EVAL_460;
  reg [1:0] _EVAL_461;
  wire  _EVAL_465;
  wire [31:0] _EVAL_466;
  wire [4:0] _EVAL_469;
  wire  _EVAL_470;
  wire  _EVAL_471;
  wire [102:0] _EVAL_472;
  wire [102:0] _EVAL_473;
  wire  _EVAL_474;
  wire  _EVAL_476;
  wire  _EVAL_477;
  wire [102:0] _EVAL_480;
  wire  _EVAL_481;
  wire [31:0] _EVAL_482;
  wire [31:0] _EVAL_483;
  wire  _EVAL_484;
  wire  _EVAL_485;
  wire  _EVAL_486;
  wire [5:0] _EVAL_488;
  wire [31:0] _EVAL_490;
  wire  _EVAL_491;
  wire  _EVAL_492;
  wire  _EVAL_493;
  wire  _EVAL_494;
  wire [4:0] _EVAL_495;
  wire  _EVAL_497;
  reg [5:0] _EVAL_498;
  wire  _EVAL_499;
  reg  _EVAL_500;
  wire  _EVAL_501;
  wire [31:0] _EVAL_502;
  wire  _EVAL_503;
  wire [31:0] _EVAL_504;
  wire [31:0] _EVAL_505;
  wire  _EVAL_506;
  wire [1:0] _EVAL_507;
  wire [1:0] _EVAL_509;
  wire  _EVAL_511;
  wire  _EVAL_512;
  wire  _EVAL_513;
  wire [31:0] _EVAL_514;
  wire  _EVAL_515;
  wire  _EVAL_516;
  wire  _EVAL_517;
  wire  _EVAL_519;
  wire [7:0] _EVAL_521;
  wire  _EVAL_523;
  wire [4:0] _EVAL_524;
  wire  _EVAL_525;
  wire  _EVAL_527;
  wire [39:0] _EVAL_528;
  wire  _EVAL_530;
  wire [31:0] _EVAL_531;
  wire [102:0] _EVAL_532;
  wire  _EVAL_533;
  wire  _EVAL_535;
  wire [31:0] _EVAL_536;
  wire  _EVAL_537;
  wire  _EVAL_539;
  reg [29:0] _EVAL_540;
  wire  _EVAL_541;
  wire  _EVAL_542;
  wire  _EVAL_543;
  wire [31:0] _EVAL_545;
  wire  _EVAL_546;
  wire [4:0] _EVAL_547;
  wire  _EVAL_548;
  wire  _EVAL_549;
  wire  _EVAL_550;
  wire [102:0] _EVAL_552;
  wire  _EVAL_553;
  wire  _EVAL_554;
  wire [4:0] _EVAL_555;
  wire  _EVAL_556;
  wire  _EVAL_558;
  wire [34:0] _EVAL_560;
  wire  _EVAL_563;
  wire [7:0] _EVAL_564;
  wire  _EVAL_565;
  wire  _EVAL_566;
  wire [1:0] _EVAL_567;
  wire  _EVAL_568;
  wire  _EVAL_569;
  wire  _EVAL_571;
  wire [57:0] _EVAL_572;
  wire  _EVAL_573;
  wire [5:0] _EVAL_575;
  wire  _EVAL_576;
  wire [102:0] _EVAL_577;
  wire  _EVAL_579;
  wire  _EVAL_580;
  wire  _EVAL_582;
  wire  _EVAL_584;
  wire  _EVAL_585;
  wire  _EVAL_587;
  wire [33:0] _EVAL_589;
  wire  _EVAL_590;
  wire  _EVAL_591;
  wire [31:0] _EVAL_592;
  wire  _EVAL_593;
  wire [31:0] _EVAL_594;
  wire  _EVAL_595;
  wire [4:0] _EVAL_596;
  wire [31:0] _EVAL_597;
  wire  _EVAL_598;
  wire [31:0] _EVAL_599;
  wire [4:0] _EVAL_602;
  wire [63:0] _EVAL_604;
  wire [31:0] _EVAL_607;
  wire [102:0] _EVAL_608;
  wire  _EVAL_610;
  reg  _EVAL_611;
  wire  _EVAL_612;
  wire [31:0] _EVAL_614;
  wire [102:0] _EVAL_616;
  reg  _EVAL_617;
  wire [31:0] _EVAL_618;
  wire [102:0] _EVAL_619;
  wire  _EVAL_620;
  wire  _EVAL_621;
  wire [31:0] _EVAL_622;
  wire  _EVAL_624;
  wire  _EVAL_625;
  wire [4:0] _EVAL_626;
  wire  _EVAL_627;
  wire  _EVAL_628;
  wire [31:0] _EVAL_629;
  reg  _EVAL_630;
  wire  _EVAL_631;
  wire  _EVAL_632;
  wire  _EVAL_634;
  wire [3:0] _EVAL_635;
  wire  _EVAL_637;
  wire  _EVAL_638;
  wire [31:0] _EVAL_639;
  wire [31:0] _EVAL_640;
  wire  _EVAL_642;
  wire  _EVAL_646;
  reg [31:0] _EVAL_647;
  wire  _EVAL_650;
  wire  _EVAL_651;
  wire  _EVAL_652;
  wire  _EVAL_653;
  wire  _EVAL_654;
  wire [29:0] _EVAL_655;
  wire  _EVAL_657;
  wire  _EVAL_658;
  wire [1:0] _EVAL_659;
  wire [4:0] _EVAL_661;
  wire  _EVAL_662;
  wire  _EVAL_663;
  reg  _EVAL_665;
  wire  _EVAL_666;
  reg  _EVAL_668;
  wire  _EVAL_670;
  wire  _EVAL_671;
  wire  _EVAL_672;
  wire  _EVAL_673;
  wire  _EVAL_674;
  wire [30:0] _EVAL_675;
  wire [31:0] _EVAL_676;
  reg [1:0] _EVAL_679;
  wire  _EVAL_681;
  wire [57:0] _EVAL_682;
  wire  _EVAL_683;
  wire  _EVAL_684;
  wire [31:0] _EVAL_685;
  wire  _EVAL_687;
  wire  _EVAL_688;
  reg [11:0] _EVAL_689;
  wire  _EVAL_691;
  wire  _EVAL_692;
  wire  _EVAL_694;
  wire [31:0] _EVAL_695;
  wire [31:0] _EVAL_696;
  wire  _EVAL_697;
  wire  _EVAL_699;
  wire  _EVAL_700;
  wire  _EVAL_701;
  wire  _EVAL_702;
  wire  _EVAL_704;
  wire [31:0] _EVAL_705;
  wire  _EVAL_706;
  wire  _EVAL_707;
  wire  _EVAL_708;
  wire  _EVAL_710;
  wire  _EVAL_711;
  wire  _EVAL_712;
  wire  _EVAL_713;
  wire  _EVAL_714;
  wire  _EVAL_715;
  wire  _EVAL_717;
  wire [31:0] _EVAL_720;
  wire  _EVAL_721;
  reg [7:0] _EVAL_722;
  wire  _EVAL_723;
  wire  _EVAL_724;
  wire [4:0] _EVAL_725;
  wire  _EVAL_726;
  wire [1:0] _EVAL_727;
  wire  _EVAL_728;
  wire  _EVAL_730;
  wire [31:0] _EVAL_732;
  wire  _EVAL_734;
  wire [7:0] _EVAL_735;
  wire  _EVAL_736;
  wire [31:0] _EVAL_737;
  wire [30:0] _EVAL_739;
  reg [2:0] _EVAL_740;
  reg  _EVAL_741;
  reg  _EVAL_743;
  wire  _EVAL_744;
  wire  _EVAL_747;
  wire  _EVAL_748;
  wire  _EVAL_753;
  wire [31:0] _EVAL_754;
  wire [1:0] _EVAL_755;
  wire  _EVAL_757;
  wire  _EVAL_759;
  wire  _EVAL_760;
  wire  _EVAL_763;
  wire [31:0] _EVAL_765;
  reg  _EVAL_767;
  wire  _EVAL_768;
  wire  _EVAL_769;
  wire [102:0] _EVAL_770;
  wire [102:0] _EVAL_771;
  wire  _EVAL_773;
  wire  _EVAL_775;
  wire  _EVAL_776;
  wire  _EVAL_778;
  wire  _EVAL_779;
  wire [3:0] _EVAL_780;
  wire  _EVAL_781;
  wire  _EVAL_782;
  wire [30:0] _EVAL_783;
  wire  _EVAL_784;
  wire  _EVAL_787;
  wire  _EVAL_791;
  wire  _EVAL_792;
  reg  _EVAL_793;
  reg  _EVAL_795;
  wire  _EVAL_796;
  wire [102:0] _EVAL_797;
  wire [31:0] _EVAL_798;
  reg  _EVAL_799;
  wire  _EVAL_800;
  wire  _EVAL_801;
  wire  _EVAL_802;
  wire  _EVAL_803;
  reg  _EVAL_804;
  wire  _EVAL_807;
  wire  _EVAL_809;
  wire [31:0] _EVAL_810;
  wire [30:0] _EVAL_811;
  wire  _EVAL_815;
  wire  _EVAL_817;
  wire [31:0] _EVAL_818;
  wire [7:0] _EVAL_819;
  reg  _EVAL_820;
  wire  _EVAL_821;
  wire  _EVAL_823;
  wire [31:0] _EVAL_824;
  wire  _EVAL_825;
  wire  _EVAL_828;
  wire  _EVAL_830;
  wire  _EVAL_831;
  wire [31:0] _EVAL_832;
  wire  _EVAL_833;
  reg  _EVAL_834;
  wire  _EVAL_835;
  wire  _EVAL_836;
  wire [31:0] _EVAL_837;
  wire  _EVAL_843;
  wire  _EVAL_844;
  wire [39:0] _EVAL_845;
  wire  _EVAL_847;
  wire [31:0] _EVAL_849;
  wire [102:0] _EVAL_850;
  wire  _EVAL_851;
  wire  _EVAL_852;
  wire [1:0] _EVAL_853;
  reg [31:0] _EVAL_855;
  wire [1:0] _EVAL_856;
  wire [102:0] _EVAL_857;
  wire  _EVAL_858;
  wire [29:0] _EVAL_860;
  wire  _EVAL_861;
  wire  _EVAL_862;
  wire  _EVAL_863;
  wire [102:0] _EVAL_865;
  wire  _EVAL_866;
  wire  _EVAL_867;
  wire [31:0] _EVAL_870;
  wire [4:0] _EVAL_871;
  reg  _EVAL_872;
  wire [1:0] _EVAL_873;
  wire  _EVAL_874;
  wire [63:0] _EVAL_875;
  wire  _EVAL_876;
  reg [1:0] _EVAL_877;
  wire  _EVAL_878;
  wire [30:0] _EVAL_879;
  wire  _EVAL_880;
  wire  _EVAL_881;
  wire  _EVAL_882;
  wire  _EVAL_883;
  wire  _EVAL_885;
  wire  _EVAL_888;
  wire [4:0] _EVAL_889;
  reg [1:0] _EVAL_890;
  reg  _EVAL_891;
  wire  _EVAL_892;
  wire [1:0] _EVAL_893;
  wire  _EVAL_895;
  wire [31:0] _EVAL_896;
  wire  _EVAL_897;
  wire [31:0] _EVAL_898;
  wire  _EVAL_899;
  wire  _EVAL_902;
  wire [31:0] _EVAL_904;
  reg  _EVAL_905;
  wire  _EVAL_906;
  wire  _EVAL_907;
  wire  _EVAL_909;
  wire [102:0] _EVAL_910;
  wire [7:0] _EVAL_911;
  wire  _EVAL_912;
  wire  _EVAL_913;
  wire  _EVAL_914;
  wire [4:0] _EVAL_915;
  wire [31:0] _EVAL_916;
  wire  _EVAL_917;
  wire [30:0] _EVAL_918;
  wire [31:0] _EVAL_919;
  wire [6:0] _EVAL_920;
  wire  _EVAL_921;
  wire  _EVAL_924;
  wire [1:0] _EVAL_926;
  wire  _EVAL_928;
  wire [31:0] _EVAL_929;
  wire [4:0] _EVAL_930;
  wire [6:0] _EVAL_931;
  wire  _EVAL_932;
  wire  _EVAL_933;
  wire  _EVAL_934;
  wire [31:0] _EVAL_935;
  wire  _EVAL_936;
  reg  _EVAL_937;
  wire  _EVAL_938;
  wire [33:0] _EVAL_939;
  wire [31:0] _EVAL_942;
  wire [31:0] _EVAL_943;
  wire  _EVAL_945;
  wire  _EVAL_947;
  reg  _EVAL_949;
  wire [102:0] _EVAL_951;
  wire  _EVAL_952;
  wire  _EVAL_954;
  wire [102:0] _EVAL_955;
  wire [31:0] _EVAL_956;
  wire  _EVAL_957;
  wire  _EVAL_958;
  wire [31:0] _EVAL_959;
  reg  _EVAL_962;
  wire [7:0] _EVAL_963;
  wire [31:0] _EVAL_964;
  reg [1:0] _EVAL_965;
  wire [18:0] _EVAL_966;
  wire [4:0] _EVAL_967;
  wire [4:0] _EVAL_968;
  wire  _EVAL_972;
  wire  _EVAL_973;
  wire  _EVAL_974;
  wire [7:0] _EVAL_975;
  wire  _EVAL_980;
  wire  _EVAL_981;
  wire  _EVAL_983;
  reg  _EVAL_985;
  wire  _EVAL_989;
  wire  _EVAL_990;
  wire [32:0] _EVAL_991;
  wire  _EVAL_995;
  wire  _EVAL_997;
  wire  _EVAL_999;
  reg [1:0] _EVAL_1001;
  wire  _EVAL_1002;
  wire  _EVAL_1003;
  wire  _EVAL_1005;
  wire [102:0] _EVAL_1006;
  wire [1:0] _EVAL_1007;
  wire  _EVAL_1009;
  wire  _EVAL_1010;
  wire  _EVAL_1012;
  wire [4:0] _EVAL_1013;
  wire  _EVAL_1014;
  wire [31:0] _EVAL_1015;
  wire  _EVAL_1016;
  reg  _EVAL_1017;
  wire  _EVAL_1018;
  wire  _EVAL_1019;
  wire  _EVAL_1022;
  wire  _EVAL_1023;
  wire  _EVAL_1024;
  wire [1:0] _EVAL_1025;
  reg  _EVAL_1027;
  wire  _EVAL_1028;
  wire [63:0] _EVAL_1029;
  wire [4:0] _EVAL_1030;
  wire  _EVAL_1031;
  reg  _EVAL_1032;
  wire  _EVAL_1034;
  wire  _EVAL_1035;
  wire  _EVAL_1036;
  wire [102:0] _EVAL_1037;
  wire [6:0] _EVAL_1038;
  wire  _EVAL_1039;
  wire [3:0] _EVAL_1040;
  wire  _EVAL_1041;
  wire  _EVAL_1042;
  wire [31:0] _EVAL_1043;
  wire [29:0] _EVAL_1046;
  wire [1:0] _EVAL_1047;
  wire  _EVAL_1048;
  wire [32:0] _EVAL_1049;
  wire  _EVAL_1050;
  wire [31:0] _EVAL_1051;
  wire  _EVAL_1052;
  wire  _EVAL_1056;
  wire  _EVAL_1057;
  wire  _EVAL_1058;
  reg [1:0] _EVAL_1059;
  wire [4:0] _EVAL_1060;
  reg [57:0] _EVAL_1062;
  wire  _EVAL_1063;
  wire [7:0] _EVAL_1064;
  wire  _EVAL_1065;
  wire  _EVAL_1066;
  wire [34:0] _EVAL_1068;
  wire  _EVAL_1069;
  reg [31:0] _EVAL_1070;
  wire  _EVAL_1072;
  wire [4:0] _EVAL_1073;
  reg  _EVAL_1075;
  wire  _EVAL_1076;
  wire  _EVAL_1080;
  wire  _EVAL_1081;
  wire  _EVAL_1082;
  wire [63:0] _EVAL_1083;
  wire  _EVAL_1084;
  wire [11:0] _EVAL_1085;
  wire [24:0] _EVAL_1086;
  wire  _EVAL_1088;
  wire  _EVAL_1090;
  wire  _EVAL_1091;
  wire  _EVAL_1092;
  wire  _EVAL_1094;
  wire [29:0] _EVAL_1095;
  wire  _EVAL_1096;
  wire  _EVAL_1097;
  wire  _EVAL_1099;
  wire [31:0] _EVAL_1100;
  wire  _EVAL_1102;
  wire  _EVAL_1103;
  wire [39:0] _EVAL_1105;
  wire [1:0] _EVAL_1107;
  wire [31:0] _EVAL_1109;
  wire  _EVAL_1110;
  wire  _EVAL_1111;
  wire  _EVAL_1112;
  reg [1:0] _EVAL_1113;
  wire [31:0] _EVAL_1114;
  wire [31:0] _EVAL_1116;
  wire  _EVAL_1118;
  wire  _EVAL_1119;
  reg  _EVAL_1120;
  wire  _EVAL_1121;
  wire [102:0] _EVAL_1122;
  wire [4:0] _EVAL_1123;
  wire [63:0] _EVAL_1124;
  wire  _EVAL_1125;
  wire [33:0] _EVAL_1126;
  wire [31:0] _EVAL_1129;
  wire  _EVAL_1130;
  wire  _EVAL_1131;
  wire [31:0] _EVAL_1132;
  wire  _EVAL_1133;
  wire  _EVAL_1136;
  wire [5:0] _EVAL_1137;
  wire [31:0] _EVAL_1140;
  wire  _EVAL_1141;
  wire  _EVAL_1142;
  wire  _EVAL_1143;
  wire  _EVAL_1144;
  wire [11:0] _EVAL_1145;
  wire  _EVAL_1146;
  wire  _EVAL_1147;
  wire  _EVAL_1150;
  wire  _EVAL_1151;
  wire [102:0] _EVAL_1153;
  reg [29:0] _EVAL_1155;
  wire  _EVAL_1157;
  reg [31:0] _EVAL_1159;
  wire [102:0] _EVAL_1160;
  reg  _EVAL_1161;
  wire  _EVAL_1164;
  wire [31:0] _EVAL_1168;
  wire [31:0] _EVAL_1169;
  wire [4:0] _EVAL_1170;
  wire  _EVAL_1172;
  wire [1:0] _EVAL_1174;
  wire  _EVAL_1175;
  wire  _EVAL_1177;
  wire  _EVAL_1178;
  wire [31:0] _EVAL_1179;
  wire  _EVAL_1180;
  wire [31:0] _EVAL_1181;
  wire  _EVAL_1182;
  wire [102:0] _EVAL_1183;
  wire [31:0] _EVAL_1186;
  reg [31:0] _EVAL_1187;
  wire  _EVAL_1189;
  wire [31:0] _EVAL_1190;
  wire  _EVAL_1191;
  wire  _EVAL_1192;
  wire  _EVAL_1194;
  wire  _EVAL_1198;
  wire [4:0] _EVAL_1200;
  wire  _EVAL_1201;
  wire  _EVAL_1202;
  wire  _EVAL_1203;
  wire  _EVAL_1204;
  reg  _EVAL_1206;
  wire  _EVAL_1208;
  wire [31:0] _EVAL_1209;
  wire  _EVAL_1210;
  wire [31:0] _EVAL_1211;
  reg [1:0] _EVAL_1212;
  reg [26:0] _EVAL_1213;
  wire  _EVAL_1214;
  wire  _EVAL_1215;
  reg [31:0] _EVAL_1217;
  wire  _EVAL_1218;
  wire [31:0] _EVAL_1219;
  wire  _EVAL_1220;
  wire [3:0] _EVAL_1221;
  wire  _EVAL_1222;
  reg  _EVAL_1227;
  wire  _EVAL_1228;
  reg  _EVAL_1229;
  wire  _EVAL_1230;
  reg  _EVAL_1231;
  wire [102:0] _EVAL_1233;
  wire [31:0] _EVAL_1235;
  wire [7:0] _EVAL_1239;
  wire  _EVAL_1240;
  wire [102:0] _EVAL_1244;
  wire  _EVAL_1245;
  wire  _EVAL_1246;
  wire  _EVAL_1248;
  wire  _EVAL_1249;
  wire  _EVAL_1250;
  wire  _EVAL_1251;
  wire  _EVAL_1254;
  wire  _EVAL_1255;
  wire  _EVAL_1256;
  wire [4:0] _EVAL_1259;
  wire [31:0] _EVAL_1260;
  wire [31:0] _EVAL_1261;
  wire  _EVAL_1262;
  wire [4:0] _EVAL_1264;
  wire [31:0] _EVAL_1265;
  wire  _EVAL_1266;
  wire  _EVAL_1270;
  wire [4:0] _EVAL_1273;
  wire [31:0] _EVAL_1274;
  wire  _EVAL_1275;
  wire [63:0] _EVAL_1279;
  reg  _EVAL_1280;
  wire [4:0] _EVAL_1283;
  wire  _EVAL_1284;
  wire  _EVAL_1285;
  wire  _EVAL_1286;
  wire  _EVAL_1287;
  wire  _EVAL_1288;
  wire  _EVAL_1289;
  wire  _EVAL_1290;
  wire  _EVAL_1291;
  wire [31:0] _EVAL_1293;
  wire [31:0] _EVAL_1297;
  wire  _EVAL_1298;
  reg  _EVAL_1300;
  wire  _EVAL_1301;
  reg [31:0] _EVAL_1302;
  wire  _EVAL_1303;
  wire [63:0] _EVAL_1304;
  reg  _EVAL_1306;
  wire  _EVAL_1308;
  wire [4:0] _EVAL_1309;
  wire  _EVAL_1310;
  wire  _EVAL_1311;
  wire  _EVAL_1312;
  wire [1:0] _EVAL_1313;
  wire  _EVAL_1315;
  wire  _EVAL_1316;
  wire  _EVAL_1318;
  wire  _EVAL_1319;
  wire  _EVAL_1321;
  wire  _EVAL_1322;
  wire  _EVAL_1323;
  wire  _EVAL_1324;
  reg  _EVAL_1326;
  wire [102:0] _EVAL_1327;
  wire  _EVAL_1328;
  wire  _EVAL_1329;
  wire  _EVAL_1330;
  wire [31:0] _EVAL_1332;
  reg [31:0] _EVAL_1334;
  wire  _EVAL_1335;
  wire  _EVAL_1336;
  wire  _EVAL_1339;
  wire [102:0] _EVAL_1340;
  wire [4:0] _EVAL_1341;
  wire  _EVAL_1342;
  reg  _EVAL_1344;
  wire  _EVAL_1345;
  wire  _EVAL_1346;
  wire  _EVAL_1347;
  wire [31:0] _EVAL_1348;
  wire  _EVAL_1349;
  wire  _EVAL_1350;
  wire  _EVAL_1351;
  wire  _EVAL_1354;
  wire [31:0] _EVAL_1355;
  reg [31:0] _EVAL_1357;
  wire  _EVAL_1358;
  wire [4:0] _EVAL_1359;
  wire  _EVAL_1360;
  wire  _EVAL_1363;
  wire  _EVAL_1364;
  wire [4:0] _EVAL_1366;
  wire  _EVAL_1367;
  wire [33:0] _EVAL_1369;
  wire  _EVAL_1371;
  wire [102:0] _EVAL_1373;
  wire  _EVAL_1374;
  wire [102:0] _EVAL_1378;
  wire [102:0] _EVAL_1379;
  wire  _EVAL_1380;
  wire  _EVAL_1381;
  reg  _EVAL_1383;
  wire [102:0] _EVAL_1384;
  wire  _EVAL_1385;
  wire  _EVAL_1386;
  wire  _EVAL_1388;
  wire [31:0] _EVAL_1389;
  wire  _EVAL_1391;
  wire [31:0] _EVAL_1392;
  wire  _EVAL_1393;
  wire  _EVAL_1395;
  wire [4:0] _EVAL_1396;
  wire  _EVAL_1398;
  reg  _EVAL_1399;
  wire  _EVAL_1401;
  wire [31:0] _EVAL_1402;
  wire  _EVAL_1404;
  wire [31:0] _EVAL_1405;
  wire  _EVAL_1406;
  wire [31:0] _EVAL_1407;
  wire  _EVAL_1410;
  wire [31:0] _EVAL_1411;
  wire  _EVAL_1413;
  wire  _EVAL_1415;
  wire [63:0] _EVAL_1416;
  wire  _EVAL_1417;
  wire  _EVAL_1418;
  wire  _EVAL_1421;
  wire  _EVAL_1422;
  wire  _EVAL_1423;
  wire  _EVAL_1424;
  wire  _EVAL_1425;
  wire  _EVAL_1427;
  wire  _EVAL_1429;
  wire  _EVAL_1430;
  wire  _EVAL_1431;
  wire [4:0] _EVAL_1436;
  wire  _EVAL_1438;
  reg [33:0] _EVAL_1439;
  wire  _EVAL_1440;
  wire [39:0] _EVAL_1441;
  wire  _EVAL_1442;
  wire  _EVAL_1444;
  wire [30:0] _EVAL_1445;
  wire [102:0] _EVAL_1447;
  wire  _EVAL_1448;
  wire [30:0] _EVAL_1450;
  wire [1:0] _EVAL_1451;
  wire  _EVAL_1452;
  wire [30:0] _EVAL_1454;
  wire [31:0] _EVAL_1455;
  wire [31:0] _EVAL_1456;
  wire  _EVAL_1457;
  wire  _EVAL_1458;
  wire  _EVAL_1460;
  wire  _EVAL_1461;
  reg  _EVAL_1463;
  wire  _EVAL_1465;
  wire  _EVAL_1468;
  wire  _EVAL_1470;
  wire  _EVAL_1471;
  wire  _EVAL_1472;
  wire  _EVAL_1476;
  reg  _EVAL_1478;
  wire [102:0] _EVAL_1479;
  wire  _EVAL_1480;
  wire [31:0] _EVAL_1481;
  wire  _EVAL_1482;
  wire [3:0] _EVAL_1483;
  wire [7:0] _EVAL_1484;
  wire  _EVAL_1485;
  wire  _EVAL_1487;
  wire  _EVAL_1489;
  wire [31:0] _EVAL_1490;
  wire [31:0] _EVAL_1492;
  wire  _EVAL_1493;
  wire  _EVAL_1495;
  reg  _EVAL_1496;
  wire [4:0] _EVAL_1497;
  wire [1:0] _EVAL_1498;
  wire  _EVAL_1500;
  wire  _EVAL_1501;
  wire  _EVAL_1502;
  wire  _EVAL_1503;
  reg  _EVAL_1504;
  reg [5:0] _EVAL_1505;
  wire  _EVAL_1509;
  wire [102:0] _EVAL_1510;
  reg [1:0] _EVAL_1511;
  wire [4:0] _EVAL_1512;
  wire [11:0] _EVAL_1514;
  wire  _EVAL_1515;
  wire [31:0] _EVAL_1516;
  wire  _EVAL_1517;
  wire  _EVAL_1518;
  wire  _EVAL_1519;
  wire  _EVAL_1520;
  wire [4:0] _EVAL_1524;
  reg [1:0] _EVAL_1525;
  wire  _EVAL_1526;
  wire  _EVAL_1527;
  wire  _EVAL_1528;
  wire  _EVAL_1529;
  wire  _EVAL_1531;
  wire  _EVAL_1532;
  wire [30:0] _EVAL_1533;
  reg  _EVAL_1534;
  wire  _EVAL_1535;
  wire [32:0] _EVAL_1536;
  wire  _EVAL_1537;
  wire  _EVAL_1539;
  wire [102:0] _EVAL_1540;
  reg [1:0] _EVAL_1541;
  wire  _EVAL_1544;
  reg  _EVAL_1545;
  wire [3:0] _EVAL_1546;
  wire  _EVAL_1549;
  wire  _EVAL_1550;
  wire [31:0] _EVAL_1551;
  wire  _EVAL_1553;
  wire [31:0] _EVAL_1554;
  wire [32:0] _EVAL_1556;
  reg  _EVAL_1557;
  wire [1:0] _EVAL_1558;
  wire  _EVAL_1560;
  wire  _EVAL_1561;
  wire [13:0] _EVAL_1562;
  wire [5:0] _EVAL_1563;
  wire  _EVAL_1564;
  wire [31:0] _EVAL_1565;
  wire [31:0] _EVAL_1566;
  wire  _EVAL_1567;
  wire  _EVAL_1568;
  wire  _EVAL_1569;
  wire [102:0] _EVAL_1571;
  wire  _EVAL_1573;
  wire [23:0] _EVAL_1574;
  wire  _EVAL_1575;
  wire [31:0] _EVAL_1580;
  wire  _EVAL_1581;
  wire [4:0] _EVAL_1583;
  wire  _EVAL_1584;
  wire  _EVAL_1586;
  wire  _EVAL_1588;
  wire [4:0] _EVAL_1589;
  wire [31:0] _EVAL_1592;
  wire [15:0] _EVAL_1593;
  wire [31:0] _EVAL_1594;
  reg  _EVAL_1595;
  wire  _EVAL_1597;
  wire  _EVAL_1598;
  wire [3:0] _EVAL_1599;
  wire  _EVAL_1600;
  wire  _EVAL_1601;
  wire  _EVAL_1602;
  wire  _EVAL_1604;
  wire  _EVAL_1607;
  wire [4:0] _EVAL_1609;
  wire [31:0] _EVAL_1612;
  wire  _EVAL_1613;
  wire [31:0] _EVAL_1616;
  reg  _EVAL_1618;
  wire  _EVAL_1619;
  reg  _EVAL_1620;
  wire [31:0] _EVAL_1621;
  wire  _EVAL_1623;
  wire  _EVAL_1625;
  wire  _EVAL_1627;
  wire [31:0] _EVAL_1628;
  wire [31:0] _EVAL_1629;
  wire  _EVAL_1630;
  wire  _EVAL_1631;
  reg [1:0] _EVAL_1633;
  wire  _EVAL_1634;
  wire  _EVAL_1635;
  wire [31:0] _EVAL_1636;
  wire  _EVAL_1637;
  wire [4:0] _EVAL_1639;
  wire [31:0] _EVAL_1640;
  wire [31:0] _EVAL_1642;
  wire  _EVAL_1643;
  wire  _EVAL_1644;
  wire  _EVAL_1645;
  wire  _EVAL_1647;
  wire [102:0] _EVAL_1648;
  wire [31:0] _EVAL_1651;
  wire [102:0] _EVAL_1652;
  wire  _EVAL_1654;
  reg  _EVAL_1657;
  wire  _EVAL_1658;
  wire  _EVAL_1659;
  wire [30:0] _EVAL_1660;
  wire [31:0] _EVAL_1661;
  wire  _EVAL_1662;
  wire  _EVAL_1663;
  wire [58:0] _EVAL_1664;
  wire  _EVAL_1665;
  wire  _EVAL_1667;
  wire [31:0] _EVAL_1668;
  wire [102:0] _EVAL_1669;
  wire [63:0] _EVAL_1670;
  reg  _EVAL_1672;
  wire [31:0] _EVAL_1677;
  wire  _EVAL_1678;
  wire  _EVAL_1679;
  wire [39:0] _EVAL_1681;
  wire  _EVAL_1682;
  wire  _EVAL_1683;
  wire [3:0] _EVAL_1684;
  wire  _EVAL_1686;
  wire  _EVAL_1687;
  wire [102:0] _EVAL_1688;
  wire  _EVAL_1689;
  wire  _EVAL_1690;
  wire  _EVAL_1691;
  wire [57:0] _EVAL_1692;
  wire  _EVAL_1693;
  reg  _EVAL_1694;
  wire  _EVAL_1695;
  reg [1:0] _EVAL_1696;
  wire [4:0] _EVAL_1697;
  wire  _EVAL_1698;
  wire  _EVAL_1699;
  wire [32:0] _EVAL_1700;
  wire  _EVAL_1701;
  wire  _EVAL_1702;
  wire  _EVAL_1705;
  wire [31:0] _EVAL_1706;
  wire [30:0] _EVAL_1707;
  wire  _EVAL_1708;
  wire  _EVAL_1709;
  wire  _EVAL_1710;
  wire  _EVAL_1712;
  wire  _EVAL_1714;
  wire  _EVAL_1715;
  wire [1:0] _EVAL_1716;
  wire  _EVAL_1717;
  wire  _EVAL_1718;
  wire  _EVAL_1719;
  wire  _EVAL_1720;
  wire  _EVAL_1721;
  wire  _EVAL_1722;
  wire  _EVAL_1723;
  wire  _EVAL_1724;
  wire [6:0] _EVAL_1725;
  wire [4:0] _EVAL_1729;
  wire [2:0] _EVAL_1730;
  wire  _EVAL_1731;
  wire  _EVAL_1732;
  reg [4:0] _EVAL_1733;
  wire [32:0] _EVAL_1734;
  wire  _EVAL_1735;
  wire  _EVAL_1736;
  wire  _EVAL_1737;
  reg [1:0] _EVAL_1738;
  wire  _EVAL_1739;
  wire [4:0] _EVAL_1740;
  wire [63:0] _EVAL_1741;
  wire  _EVAL_1742;
  wire [31:0] _EVAL_1744;
  wire  _EVAL_1745;
  wire [102:0] _EVAL_1748;
  wire  _EVAL_1749;
  wire  _EVAL_1750;
  wire  _EVAL_1752;
  wire  _EVAL_1753;
  wire [6:0] _EVAL_1755;
  wire [30:0] _EVAL_1756;
  reg  _EVAL_1757;
  wire  _EVAL_1758;
  wire  _EVAL_1759;
  wire  _EVAL_1760;
  reg  _EVAL_1761;
  wire [31:0] _EVAL_1762;
  wire [4:0] _EVAL_1764;
  wire [31:0] _EVAL_1765;
  wire [31:0] _EVAL_1766;
  wire  _EVAL_1767;
  wire  _EVAL_1768;
  wire [4:0] _EVAL_1770;
  wire  _EVAL_1771;
  wire [102:0] _EVAL_1773;
  wire  _EVAL_1775;
  wire [4:0] _EVAL_1776;
  wire [31:0] _EVAL_1777;
  wire  _EVAL_1778;
  wire  _EVAL_1779;
  wire [29:0] _EVAL_1782;
  wire [6:0] _EVAL_1783;
  wire  _EVAL_1785;
  wire [7:0] _EVAL_1787;
  reg  _EVAL_1788;
  wire  _EVAL_1789;
  wire  _EVAL_1790;
  wire [4:0] _EVAL_1792;
  wire  _EVAL_1793;
  wire  _EVAL_1794;
  wire  _EVAL_1795;
  reg  _EVAL_1796;
  wire  _EVAL_1797;
  wire [57:0] _EVAL_1798;
  wire  _EVAL_1800;
  wire  _EVAL_1801;
  wire  _EVAL_1802;
  wire  _EVAL_1803;
  wire  _EVAL_1804;
  wire  _EVAL_1806;
  wire [1:0] _EVAL_1807;
  wire  _EVAL_1808;
  wire  _EVAL_1809;
  wire [7:0] _EVAL_1810;
  wire [7:0] _EVAL_1812;
  reg [29:0] _EVAL_1813;
  wire  _EVAL_1816;
  reg [33:0] _EVAL_1817;
  wire  _EVAL_1818;
  wire  _EVAL_1819;
  wire  _EVAL_1820;
  wire  _EVAL_1821;
  wire [102:0] _EVAL_1822;
  wire [31:0] _EVAL_1823;
  wire  _EVAL_1824;
  wire [1:0] _EVAL_1825;
  wire [102:0] _EVAL_1826;
  wire [31:0] _EVAL_1827;
  reg [1:0] _EVAL_1828;
  wire  _EVAL_1829;
  wire  _EVAL_1830;
  wire [102:0] _EVAL_1832;
  wire [57:0] _EVAL_1833;
  wire [33:0] _EVAL_1834;
  wire [1:0] _EVAL_1835;
  wire  _EVAL_1836;
  wire  _EVAL_1838;
  wire  _EVAL_1839;
  wire  _EVAL_1841;
  wire  _EVAL_1845;
  reg [31:0] _EVAL_1847;
  wire  _EVAL_1848;
  reg  _EVAL_1849;
  wire  _EVAL_1850;
  wire  _EVAL_1851;
  wire  _EVAL_1852;
  wire  _EVAL_1854;
  wire [4:0] _EVAL_1855;
  wire  _EVAL_1856;
  wire [30:0] _EVAL_1857;
  reg [1:0] _EVAL_1858;
  wire [31:0] _EVAL_1859;
  wire  _EVAL_1860;
  wire  _EVAL_1861;
  wire  _EVAL_1862;
  wire [102:0] _EVAL_1863;
  wire  _EVAL_1866;
  reg  _EVAL_1867;
  wire  _EVAL_1869;
  reg [31:0] _EVAL_1870;
  wire  _EVAL_1872;
  wire  _EVAL_1873;
  wire [6:0] _EVAL_1874;
  wire [29:0] _EVAL_1876;
  wire  _EVAL_1877;
  reg  _EVAL_1878;
  wire  _EVAL_1879;
  wire  _EVAL_1880;
  wire  _EVAL_1881;
  wire [31:0] _EVAL_1882;
  wire [7:0] _EVAL_1883;
  wire  _EVAL_1884;
  wire  _EVAL_1885;
  wire  _EVAL_1886;
  wire [7:0] _EVAL_1887;
  wire [15:0] _EVAL_1888;
  wire [31:0] _EVAL_1890;
  wire  _EVAL_1891;
  wire  _EVAL_1892;
  wire  _EVAL_1893;
  wire [39:0] _EVAL_1894;
  wire  _EVAL_1896;
  wire  _EVAL_1897;
  wire  _EVAL_1898;
  wire  _EVAL_1901;
  wire  _EVAL_1903;
  wire [1:0] _EVAL_1904;
  wire  _EVAL_1905;
  wire  _EVAL_1906;
  wire  _EVAL_1907;
  wire [32:0] _EVAL_1909;
  reg [29:0] _EVAL_1910;
  wire  _EVAL_1911;
  wire  _EVAL_1912;
  wire [3:0] _EVAL_1913;
  wire [31:0] _EVAL_1914;
  wire  _EVAL_1915;
  wire  _EVAL_1916;
  reg  _EVAL_1918;
  wire  _EVAL_1919;
  reg  _EVAL_1920;
  wire  _EVAL_1921;
  wire [31:0] _EVAL_1922;
  wire  _EVAL_1923;
  wire  _EVAL_1924;
  wire [31:0] _EVAL_1925;
  wire  _EVAL_1926;
  wire  _EVAL_1927;
  wire  _EVAL_1928;
  wire  _EVAL_1929;
  wire  _EVAL_1930;
  wire  _EVAL_1931;
  wire [4:0] _EVAL_1933;
  wire [4:0] _EVAL_1934;
  reg  _EVAL_1935;
  wire  _EVAL_1936;
  wire  _EVAL_1938;
  wire  _EVAL_1939;
  wire [6:0] _EVAL_1940;
  wire [102:0] _EVAL_1941;
  wire [102:0] _EVAL_1942;
  wire [6:0] _EVAL_1944;
  wire  _EVAL_1945;
  wire [1:0] _EVAL_1946;
  reg  _EVAL_1947;
  wire  _EVAL_1948;
  wire [30:0] _EVAL_1949;
  wire [30:0] _EVAL_1950;
  wire  _EVAL_1952;
  wire  _EVAL_1953;
  wire [4:0] _EVAL_1954;
  reg  _EVAL_1955;
  wire  _EVAL_1956;
  wire  _EVAL_1957;
  wire  _EVAL_1958;
  reg [31:0] _EVAL_1959;
  wire [31:0] _EVAL_1961;
  wire  _EVAL_1962;
  wire  _EVAL_1963;
  wire  _EVAL_1964;
  reg  _EVAL_1967;
  wire [6:0] _EVAL_1968;
  wire [31:0] _EVAL_1969;
  wire [39:0] _EVAL_1970;
  wire  _EVAL_1971;
  wire [1:0] _EVAL_1976;
  wire  _EVAL_1977;
  reg [31:0] _EVAL_1978;
  wire  _EVAL_1981;
  wire  _EVAL_1983;
  wire  _EVAL_1984;
  wire [30:0] _EVAL_1985;
  wire  _EVAL_1987;
  wire  _EVAL_1988;
  wire [1:0] _EVAL_1989;
  wire  _EVAL_1990;
  wire [31:0] _EVAL_1991;
  wire [39:0] _EVAL_1992;
  wire [31:0] _EVAL_1993;
  wire  _EVAL_1994;
  wire  _EVAL_1995;
  wire  _EVAL_1997;
  wire [32:0] _EVAL_1998;
  wire [31:0] _EVAL_1999;
  wire  _EVAL_2000;
  wire [1:0] _EVAL_2003;
  wire  _EVAL_2004;
  wire  _EVAL_2006;
  wire  _EVAL_2007;
  wire  _EVAL_2009;
  wire [11:0] _EVAL_2011;
  wire [31:0] _EVAL_2013;
  wire  _EVAL_2014;
  wire [102:0] _EVAL_2015;
  wire [31:0] _EVAL_2016;
  wire  _EVAL_2017;
  wire  _EVAL_2018;
  wire  _EVAL_2020;
  wire  _EVAL_2021;
  wire [4:0] _EVAL_2022;
  wire  _EVAL_2024;
  wire [31:0] _EVAL_2025;
  wire  _EVAL_2026;
  wire  _EVAL_2027;
  wire [63:0] _EVAL_2028;
  wire [31:0] _EVAL_2029;
  wire  _EVAL_2030;
  wire [3:0] _EVAL_2031;
  wire [102:0] _EVAL_2032;
  wire  _EVAL_2033;
  wire  _EVAL_2034;
  wire [1:0] _EVAL_2035;
  wire  _EVAL_2036;
  wire  _EVAL_2037;
  wire [102:0] _EVAL_2039;
  wire  _EVAL_2041;
  reg [31:0] _EVAL_2042;
  wire [4:0] _EVAL_2043;
  wire  _EVAL_2044;
  wire [4:0] _EVAL_2045;
  wire [31:0] _EVAL_2046;
  wire  _EVAL_2047;
  wire [30:0] _EVAL_2048;
  wire [31:0] _EVAL_2049;
  wire  _EVAL_2052;
  wire  _EVAL_2053;
  wire [30:0] _EVAL_2054;
  wire  _EVAL_2055;
  wire [31:0] _EVAL_2056;
  wire  _EVAL_2057;
  wire [31:0] _EVAL_2058;
  wire [102:0] _EVAL_2059;
  wire  _EVAL_2060;
  wire  _EVAL_2061;
  wire  _EVAL_2062;
  wire  _EVAL_2063;
  wire  _EVAL_2064;
  wire  _EVAL_2065;
  wire  _EVAL_2066;
  wire  _EVAL_2067;
  reg  _EVAL_2069;
  wire  _EVAL_2071;
  wire  _EVAL_2072;
  wire  _EVAL_2073;
  wire  _EVAL_2074;
  reg  _EVAL_2075;
  wire [3:0] _EVAL_2077;
  wire [31:0] _EVAL_2078;
  wire  _EVAL_2079;
  wire  _EVAL_2080;
  reg [1:0] _EVAL_2082;
  wire [31:0] _EVAL_2084;
  wire [31:0] _EVAL_2085;
  wire  _EVAL_2086;
  wire  _EVAL_2087;
  wire  _EVAL_2088;
  wire [1:0] _EVAL_2089;
  wire [4:0] _EVAL_2091;
  wire  _EVAL_2092;
  wire  _EVAL_2093;
  wire [1:0] _EVAL_2096;
  wire  _EVAL_2098;
  reg [31:0] _EVAL_2099;
  wire  _EVAL_2102;
  wire  _EVAL_2103;
  wire  _EVAL_2104;
  wire [3:0] _EVAL_2105;
  wire  _EVAL_2107;
  wire  _EVAL_2108;
  wire  _EVAL_2109;
  wire  _EVAL_2110;
  wire  _EVAL_2112;
  wire [29:0] _EVAL_2113;
  wire [4:0] _EVAL_2114;
  wire [31:0] _EVAL_2117;
  wire  _EVAL_2119;
  wire  _EVAL_2120;
  wire  _EVAL_2121;
  wire  _EVAL_2122;
  wire [63:0] _EVAL_2124;
  wire [3:0] _EVAL_2126;
  wire  _EVAL_2127;
  reg [31:0] _EVAL_2128;
  wire  _EVAL_2129;
  wire  _EVAL_2130;
  wire  _EVAL_2131;
  wire  _EVAL_2132;
  wire [33:0] _EVAL_2133;
  wire [4:0] _EVAL_2134;
  wire [31:0] _EVAL_2135;
  wire [1:0] _EVAL_2137;
  wire [31:0] _EVAL_2138;
  wire  _EVAL_2140;
  wire  _EVAL_2142;
  wire  _EVAL_2143;
  wire [3:0] _EVAL_2144;
  wire  _EVAL_2145;
  wire  _EVAL_2146;
  wire  _EVAL_2147;
  wire [31:0] _EVAL_2148;
  reg  _EVAL_2149;
  wire [4:0] _EVAL_2150;
  wire  _EVAL_2151;
  wire  _EVAL_2153;
  wire [102:0] _EVAL_2154;
  reg  _EVAL_2159;
  wire [31:0] _EVAL_2160;
  wire  _EVAL_2162;
  reg [1:0] _EVAL_2163;
  wire [39:0] _EVAL_2164;
  wire  _EVAL_2165;
  wire [31:0] _EVAL_2166;
  wire [57:0] _EVAL_2168;
  wire  _EVAL_2169;
  wire [4:0] _EVAL_2170;
  wire  _EVAL_2171;
  wire [31:0] _EVAL_2172;
  wire [32:0] _EVAL_2173;
  reg  _EVAL_2174;
  wire [63:0] _EVAL_2175;
  wire  _EVAL_2177;
  wire  _EVAL_2178;
  wire  _EVAL_2179;
  wire [39:0] _EVAL_2180;
  wire  _EVAL_2181;
  reg [1:0] _EVAL_2182;
  wire [31:0] _EVAL_2183;
  wire  _EVAL_2184;
  reg  _EVAL_2185;
  wire  _EVAL_2188;
  wire  _EVAL_2189;
  wire  _EVAL_2190;
  wire  _EVAL_2191;
  wire  _EVAL_2192;
  wire  _EVAL_2193;
  wire [102:0] _EVAL_2195;
  wire  _EVAL_2196;
  wire [102:0] _EVAL_2197;
  wire [4:0] _EVAL_2198;
  wire  _EVAL_2199;
  wire  _EVAL_2200;
  wire  _EVAL_2202;
  wire  _EVAL_2206;
  wire [4:0] _EVAL_2208;
  wire [31:0] _EVAL_2209;
  wire  _EVAL_2210;
  wire  _EVAL_2211;
  wire  _EVAL_2212;
  wire  _EVAL_2214;
  wire  _EVAL_2217;
  wire  _EVAL_2218;
  wire  _EVAL_2219;
  wire  _EVAL_2221;
  wire [102:0] _EVAL_2223;
  wire  _EVAL_2225;
  wire  _EVAL_2226;
  wire  _EVAL_2232;
  wire [31:0] _EVAL_2234;
  wire  _EVAL_2239;
  wire  _EVAL_2241;
  wire [102:0] _EVAL_2242;
  wire [39:0] _EVAL_2243;
  wire  _EVAL_2244;
  reg [31:0] _EVAL_2245;
  wire  _EVAL_2246;
  wire  _EVAL_2247;
  reg [5:0] _EVAL_2248;
  wire  _EVAL_2249;
  wire  _EVAL_2250;
  wire  _EVAL_2251;
  wire  _EVAL_2253;
  wire [102:0] _EVAL_2255;
  wire  _EVAL_2256;
  wire  _EVAL_2257;
  wire  _EVAL_2258;
  wire  _EVAL_2260;
  reg [29:0] _EVAL_2262;
  wire [31:0] _EVAL_2263;
  wire  _EVAL_2265;
  wire [31:0] _EVAL_2266;
  wire  _EVAL_2267;
  wire  _EVAL_2268;
  wire  _EVAL_2269;
  wire  _EVAL_2270;
  wire  _EVAL_2271;
  reg  _EVAL_2272;
  wire  _EVAL_2274;
  wire  _EVAL_2276;
  wire  _EVAL_2277;
  wire  _EVAL_2278;
  wire  _EVAL_2279;
  wire [7:0] _EVAL_2280;
  wire [30:0] _EVAL_2282;
  wire  _EVAL_2283;
  wire  _EVAL_2284;
  wire [30:0] _EVAL_2285;
  wire  _EVAL_2291;
  wire  _EVAL_2292;
  wire  _EVAL_2294;
  wire  _EVAL_2295;
  wire  _EVAL_2296;
  reg [1:0] _EVAL_2297;
  reg  _EVAL_2301;
  wire [31:0] _EVAL_2303;
  wire [31:0] _EVAL_2304;
  wire [31:0] _EVAL_2305;
  wire  _EVAL_2306;
  wire  _EVAL_2307;
  wire  _EVAL_2309;
  wire  _EVAL_2310;
  wire [102:0] _EVAL_2313;
  wire [31:0] _EVAL_2314;
  reg [31:0] _EVAL_2315;
  wire  _EVAL_2316;
  wire [102:0] _EVAL_2318;
  wire [63:0] _EVAL_2319;
  wire  _EVAL_2320;
  wire [4:0] _EVAL_2321;
  wire  _EVAL_2322;
  wire  _EVAL_2323;
  wire  _EVAL_2325;
  wire  _EVAL_2326;
  wire [30:0] _EVAL_2327;
  wire [39:0] _EVAL_2328;
  reg [31:0] _EVAL_2329;
  wire  _EVAL_2330;
  reg  _EVAL_2331;
  wire [31:0] _EVAL_2333;
  wire [33:0] _EVAL_2334;
  wire [30:0] _EVAL_2335;
  wire [31:0] _EVAL_2336;
  wire  _EVAL_2338;
  wire  _EVAL_2339;
  wire [1:0] _EVAL_2340;
  reg [5:0] _EVAL_2342;
  wire  _EVAL_2343;
  wire  _EVAL_2344;
  wire [39:0] _EVAL_2345;
  wire  _EVAL_2346;
  wire [1:0] _EVAL_2347;
  wire  _EVAL_2349;
  wire  _EVAL_2350;
  reg [2:0] _EVAL_2352;
  wire  _EVAL_2357;
  wire  _EVAL_2358;
  wire  _EVAL_2359;
  wire  _EVAL_2361;
  wire [31:0] _EVAL_2363;
  wire  _EVAL_2365;
  reg  _EVAL_2366;
  wire [31:0] _EVAL_2367;
  wire  _EVAL_2368;
  wire  _EVAL_2369;
  wire  _EVAL_2371;
  wire  _EVAL_2372;
  wire [31:0] _EVAL_2374;
  wire  _EVAL_2376;
  wire  _EVAL_2377;
  wire  _EVAL_2378;
  wire [16:0] _EVAL_2379;
  wire [31:0] _EVAL_2382;
  wire [2:0] _EVAL_2385;
  wire  _EVAL_2386;
  wire  _EVAL_2387;
  wire  _EVAL_2389;
  wire [39:0] _EVAL_2390;
  reg  _EVAL_2391;
  wire [31:0] _EVAL_2392;
  wire  _EVAL_2393;
  wire [30:0] _EVAL_2394;
  wire  _EVAL_2396;
  wire  _EVAL_2397;
  wire  _EVAL_2398;
  wire [31:0] _EVAL_2399;
  wire  _EVAL_2400;
  wire  _EVAL_2401;
  wire [1:0] _EVAL_2402;
  wire  _EVAL_2404;
  wire [6:0] _EVAL_2405;
  wire  _EVAL_2409;
  wire  _EVAL_2410;
  wire  _EVAL_2411;
  wire [4:0] _EVAL_2412;
  wire [102:0] _EVAL_2413;
  wire [15:0] _EVAL_2414;
  wire [31:0] _EVAL_2415;
  wire  _EVAL_2416;
  wire  _EVAL_2417;
  reg [29:0] _EVAL_2418;
  reg  _EVAL_2420;
  wire  _EVAL_2421;
  reg  _EVAL_2422;
  wire  _EVAL_2423;
  reg  _EVAL_2425;
  reg  _EVAL_2426;
  wire [31:0] _EVAL_2427;
  wire  _EVAL_2428;
  wire [6:0] _EVAL_2429;
  wire  _EVAL_2430;
  wire  _EVAL_2432;
  wire  _EVAL_2433;
  wire [1:0] _EVAL_2434;
  wire [30:0] _EVAL_2435;
  wire  _EVAL_2436;
  wire [31:0] _EVAL_2437;
  wire  _EVAL_2439;
  wire  _EVAL_2440;
  wire [31:0] _EVAL_2441;
  wire [30:0] _EVAL_2442;
  wire [31:0] _EVAL_2444;
  wire [63:0] _EVAL_2445;
  wire [31:0] _EVAL_2446;
  wire  _EVAL_2447;
  wire [31:0] _EVAL_2448;
  wire [102:0] _EVAL_2449;
  reg  _EVAL_2451;
  wire  _EVAL_2452;
  wire  _EVAL_2454;
  wire  _EVAL_2456;
  wire  _EVAL_2457;
  wire [102:0] _EVAL_2460;
  reg  _EVAL_2461;
  wire  _EVAL_2462;
  wire [102:0] _EVAL_2463;
  reg  _EVAL_2465;
  wire  _EVAL_2466;
  wire  _EVAL_2467;
  wire  _EVAL_2468;
  wire [4:0] _EVAL_2469;
  wire [102:0] _EVAL_2471;
  wire  _EVAL_2473;
  wire  _EVAL_2474;
  wire  _EVAL_2475;
  wire [102:0] _EVAL_2476;
  wire [4:0] _EVAL_2477;
  wire [31:0] _EVAL_2478;
  wire  _EVAL_2479;
  wire [30:0] _EVAL_2480;
  reg [1:0] _EVAL_2481;
  wire [31:0] _EVAL_2482;
  wire  _EVAL_2484;
  wire  _EVAL_2485;
  wire [31:0] _EVAL_2486;
  wire [31:0] _EVAL_2487;
  wire  _EVAL_2488;
  wire  _EVAL_2489;
  wire [31:0] _EVAL_2490;
  wire  _EVAL_2491;
  reg [31:0] _EVAL_2492;
  wire  _EVAL_2493;
  wire  _EVAL_2494;
  wire  _EVAL_2495;
  wire  _EVAL_2496;
  wire [102:0] _EVAL_2497;
  wire [31:0] _EVAL_2498;
  wire  _EVAL_2500;
  wire  _EVAL_2501;
  wire [3:0] _EVAL_2502;
  wire  _EVAL_2503;
  wire  _EVAL_2504;
  wire  _EVAL_2505;
  wire  _EVAL_2508;
  wire [58:0] _EVAL_2510;
  wire [31:0] _EVAL_2511;
  wire [31:0] _EVAL_2512;
  wire  _EVAL_2513;
  wire  _EVAL_2514;
  wire  _EVAL_2516;
  wire  _EVAL_2517;
  wire  _EVAL_2518;
  wire [7:0] _EVAL_2519;
  wire  _EVAL_2520;
  reg  _EVAL_2521;
  wire [31:0] _EVAL_2522;
  wire  _EVAL_2524;
  wire  _EVAL_2527;
  wire  _EVAL_2528;
  wire  _EVAL_2529;
  wire  _EVAL_2530;
  reg  _EVAL_2532;
  wire [6:0] _EVAL_2534;
  wire [14:0] _EVAL_2535;
  wire  _EVAL_2536;
  wire  _EVAL_2537;
  wire  _EVAL_2538;
  wire [3:0] _EVAL_2541;
  wire [31:0] _EVAL_2542;
  wire [31:0] _EVAL_2543;
  wire  _EVAL_2544;
  wire  _EVAL_2547;
  wire  _EVAL_2548;
  wire [31:0] _EVAL_2549;
  reg [57:0] _EVAL_2550;
  wire  _EVAL_2551;
  assign _EVAL_117 = _EVAL_1399;
  assign _EVAL_1182 = _EVAL_286 | _EVAL_434;
  assign _EVAL_2387 = _EVAL_1222 & _EVAL_773;
  assign _EVAL_2078 = ~_EVAL_482;
  assign _EVAL_213 = _EVAL_610 | _EVAL_834;
  assign _EVAL_1023 = _EVAL_1551[13];
  assign _EVAL_1201 = _EVAL_332 & _EVAL_1240;
  assign _EVAL_1291 = _EVAL_113 == 12'hc8b;
  assign _EVAL_253 = _EVAL_2142 ? 5'hd : _EVAL_626;
  assign _EVAL_275 = _EVAL_862 | _EVAL_584;
  assign _EVAL_1140 = _EVAL_2064 ? _EVAL_2042 : 32'h0;
  assign _EVAL_492 = _EVAL_2225 | _EVAL_215;
  assign _EVAL_1913 = {_EVAL_1144, 3'h0};
  assign _EVAL_627 = _EVAL_711 | _EVAL_2007;
  assign _EVAL_1515 = _EVAL_1861 | _EVAL_448;
  assign _EVAL_2385 = _EVAL_2069 ? 3'h4 : {{1'd0}, _EVAL_2434};
  assign _EVAL_1584 = _EVAL_759 | _EVAL_1298;
  assign _EVAL_2071 = _EVAL_702 | _EVAL_389;
  assign _EVAL_1834 = _EVAL_1992[39:6];
  assign _EVAL_137 = _EVAL_2174;
  assign _EVAL_2129 = _EVAL_2067 | _EVAL_1722;
  assign _EVAL_1085 = _EVAL_113 & 12'hc10;
  assign _EVAL_1480 = _EVAL_151 == 12'hc02;
  assign _EVAL_1544 = _EVAL_744 | _EVAL_1489;
  assign _EVAL_1034 = _EVAL_1458 | _EVAL_582;
  assign _EVAL_1500 = _EVAL_280[2];
  assign _EVAL_2382 = _EVAL_291 ? _EVAL_2099 : _EVAL_1392;
  assign _EVAL_2473 = _EVAL_2474 | _EVAL_2069;
  assign _EVAL_1102 = _EVAL_708 | _EVAL_914;
  assign _EVAL_324 = _EVAL_1845 & _EVAL_1097;
  assign _EVAL_1451 = 2'h2 == _EVAL_1541 ? _EVAL_2082 : _EVAL_853;
  assign _EVAL_2198 = _EVAL_895 ? 5'h1 : _EVAL_1639;
  assign _EVAL_2009 = _EVAL_1598 | _EVAL_757;
  assign _EVAL_1719 = ~_EVAL_1601;
  assign _EVAL_434 = _EVAL_113 == 12'hb1f;
  assign _EVAL_700 = _EVAL_402[3];
  assign _EVAL_662 = _EVAL_621 | _EVAL_2475;
  assign _EVAL_2430 = _EVAL_66 & _EVAL_1306;
  assign _EVAL_2505 = _EVAL_151 == 12'h3b2;
  assign _EVAL_2260 = _EVAL_113 == 12'h32e;
  assign _EVAL_2543 = _EVAL_291 ? _EVAL_2315 : _EVAL_2512;
  assign _EVAL_1553 = _EVAL_113 == 12'hc14;
  assign _EVAL_1112 = _EVAL_2535[3];
  assign _EVAL_1512 = _EVAL_1143 ? 5'h15 : _EVAL_1497;
  assign _EVAL_1246 = _EVAL_591 | _EVAL_1682;
  assign _EVAL_501 = _EVAL_2490[15];
  assign _EVAL_1571 = {{39'd0}, _EVAL_1741};
  assign _EVAL_828 = _EVAL_113 == 12'hb10;
  assign _EVAL_2482 = _EVAL_2320 ? _EVAL_325 : _EVAL_1187;
  assign _EVAL_1938 = _EVAL_113 == 12'h327;
  assign _EVAL_186 = _EVAL_1657;
  assign _EVAL_2325 = _EVAL_454 & _EVAL_304;
  assign _EVAL_2441 = _EVAL_1065 ? _EVAL_1265 : {{2'd0}, _EVAL_2262};
  assign _EVAL_911 = {_EVAL_454,2'h0,_EVAL_2481,_EVAL_1231,_EVAL_370,_EVAL_2159};
  assign _EVAL_35 = _EVAL_96;
  assign _EVAL_1736 = ~_EVAL_491;
  assign _EVAL_1423 = _EVAL_1427 | _EVAL_1010;
  assign _EVAL_1150 = ~_EVAL_1539;
  assign _EVAL_1468 = _EVAL_1787[0];
  assign _EVAL_1954 = _EVAL_2475 ? 5'h0 : _EVAL_1366;
  assign _EVAL_1879 = _EVAL_2508 | _EVAL_2044;
  assign _EVAL_1575 = ~_EVAL_2211;
  assign _EVAL_2274 = _EVAL_1848 | _EVAL_1142;
  assign _EVAL_2530 = _EVAL_151 == 12'h7b1;
  assign _EVAL_2494 = _EVAL_113 == 12'hb87;
  assign _EVAL_1574 = _EVAL_2490[31:8];
  assign _EVAL_149 = _EVAL_366;
  assign _EVAL_488 = {{5'd0}, _EVAL_1679};
  assign _EVAL_1147 = _EVAL_151 == 12'h7c0;
  assign _EVAL_1076 = ~_EVAL_1306;
  assign _EVAL_70 = _EVAL_130;
  assign _EVAL_2401 = _EVAL_2371 ? _EVAL_277 : _EVAL_1534;
  assign _EVAL_1956 = _EVAL_646 | _EVAL_1885;
  assign _EVAL_2446 = _EVAL_1065 ? _EVAL_1566 : {{30'd0}, _EVAL_1541};
  assign _EVAL_730 = _EVAL_402[28];
  assign _EVAL_71 = _EVAL_28;
  assign _EVAL_242 = _EVAL_113 == 12'hc98;
  assign _EVAL_2413 = {{71'd0}, _EVAL_2336};
  assign _EVAL_432 = _EVAL_1903 | _EVAL_2000;
  assign _EVAL_93 = _EVAL_1967;
  assign _EVAL_1734 = {_EVAL_879,2'h3};
  assign _EVAL_254 = _EVAL_1065 ? _EVAL_2448 : {{2'd0}, _EVAL_227};
  assign _EVAL_1890 = _EVAL_622 & _EVAL_490;
  assign _EVAL_1441 = {_EVAL_2280,_EVAL_1481};
  assign _EVAL_628 = _EVAL_113 == 12'hb04;
  assign _EVAL_983 = _EVAL_306[0];
  assign _EVAL_2306 = _EVAL_151 == 12'h350;
  assign _EVAL_587 = _EVAL_1915 | _EVAL_1367;
  assign _EVAL_801 = _EVAL_2268 | _EVAL_2272;
  assign _EVAL_825 = _EVAL_2182 < _EVAL_1174;
  assign _EVAL_952 = _EVAL_113 == 12'hc8d;
  assign _EVAL_913 = _EVAL_151 == 12'h3b6;
  assign _EVAL_2544 = _EVAL_1551[29];
  assign _EVAL_1174 = _EVAL_113[9:8];
  assign _EVAL_2428 = _EVAL_1838 | _EVAL_1561;
  assign _EVAL_589 = _EVAL_2164[39:6];
  assign _EVAL_1180 = _EVAL_618[11];
  assign _EVAL_530 = _EVAL_113 == 12'h330;
  assign _EVAL_2517 = _EVAL_1551[31];
  assign _EVAL_1448 = _EVAL_113 == 12'h3a1;
  assign _EVAL_1770 = _EVAL_730 ? 5'h1c : _EVAL_1341;
  assign _EVAL_87 = _EVAL_359;
  assign _EVAL_2104 = _EVAL_492 | _EVAL_1249;
  assign _EVAL_1934 = _EVAL_2162 ? 5'h1b : _EVAL_1123;
  assign _EVAL_1189 = _EVAL_113 == 12'hb19;
  assign _EVAL_2108 = _EVAL_2535[14];
  assign _EVAL_608 = {{39'd0}, _EVAL_604};
  assign _EVAL_545 = ~_EVAL_1978;
  assign _EVAL_1297 = _EVAL_2371 ? _EVAL_1355 : _EVAL_1070;
  assign _EVAL_2107 = _EVAL_1983 ? _EVAL_192 : _EVAL_892;
  assign _EVAL_2309 = _EVAL_113 == 12'hc92;
  assign _EVAL_1775 = _EVAL_2182 == 2'h1;
  assign _EVAL_528 = {_EVAL_1439,_EVAL_1505};
  assign _EVAL_2175 = _EVAL_1480 ? _EVAL_1416 : 64'h0;
  assign _EVAL_681 = _EVAL_1218 | _EVAL_1250;
  assign _EVAL_550 = _EVAL_494 | _EVAL_20;
  assign _EVAL_1311 = _EVAL_151 == 12'hb83;
  assign _EVAL_67 = 2'h0;
  assign _EVAL_1065 = _EVAL_2129 | _EVAL_2087;
  assign _EVAL_517 = _EVAL_1562[7];
  assign _EVAL_1829 = _EVAL_113 == 12'h334;
  assign _EVAL_2085 = _EVAL_405 + 31'h1;
  assign _EVAL_1198 = _EVAL_240 | _EVAL_1081;
  assign _EVAL_566 = _EVAL_113 == 12'h7b2;
  assign _EVAL_1930 = _EVAL_151 == 12'hc03;
  assign _EVAL_164 = _EVAL_2420;
  assign _EVAL_15 = _EVAL_1049[31:0];
  assign _EVAL_1804 = _EVAL_1562[5];
  assign _EVAL_1642 = {_EVAL_1450, 1'h0};
  assign _EVAL_692 = _EVAL_113 == 12'hc91;
  assign _EVAL_1906 = _EVAL_113 == 12'hb95;
  assign _EVAL_1082 = _EVAL_1619 | _EVAL_2310;
  assign _EVAL_2358 = _EVAL_402[30];
  assign _EVAL_1391 = _EVAL_402[1];
  assign _EVAL_114 = _EVAL_2473 & _EVAL_2109;
  assign _EVAL_1619 = _EVAL_1544 | _EVAL_2217;
  assign _EVAL_771 = {{71'd0}, _EVAL_2314};
  assign _EVAL_192 = _EVAL_2371 ? _EVAL_2218 : _EVAL_1399;
  assign _EVAL_1729 = _EVAL_2358 ? 5'h1e : _EVAL_336;
  assign _EVAL_2151 = _EVAL_402[16];
  assign _EVAL_1476 = _EVAL_113 == 12'h7c1;
  assign _EVAL_1702 = _EVAL_151 == 12'h353;
  assign _EVAL_1519 = _EVAL_1787[1];
  assign _EVAL_107 = _EVAL_460;
  assign _EVAL_1663 = ~_EVAL_355;
  assign _EVAL_912 = _EVAL_1787[7];
  assign _EVAL_1528 = _EVAL_2256 & _EVAL_1994;
  assign _EVAL_1592 = _EVAL_291 ? _EVAL_2329 : _EVAL_1114;
  assign _EVAL_2386 = _EVAL_1551[4];
  assign _EVAL_502 = _EVAL_1124[63:32];
  assign _EVAL_2035 = _EVAL_1698 ? 2'h3 : _EVAL_2182;
  assign _EVAL_1985 = ~_EVAL_1949;
  assign _EVAL_2334 = _EVAL_1441[39:6];
  assign _EVAL_1339 = _EVAL_2291 & _EVAL_1623;
  assign _EVAL_1369 = _EVAL_560[33:0];
  assign _EVAL_493 = _EVAL_1809 | _EVAL_456;
  assign _EVAL_1514 = {_EVAL_1757,_EVAL_1545,_EVAL_611,_EVAL_740,_EVAL_2352,_EVAL_1496,_EVAL_237};
  assign _EVAL_519 = _EVAL_2415 == 32'h100000;
  assign _EVAL_491 = _EVAL_1733[2];
  assign _EVAL_1630 = _EVAL_113 == 12'hb16;
  assign _EVAL_849 = ~_EVAL_2522;
  assign _EVAL_333 = 2'h1 == _EVAL_1541 ? _EVAL_1618 : _EVAL_2331;
  assign _EVAL_427 = _EVAL_809 ? 2'h2 : 2'h1;
  assign _EVAL_148 = _EVAL_1813;
  assign _EVAL_2067 = _EVAL_134 == 3'h6;
  assign _EVAL_1797 = _EVAL_662 | _EVAL_2386;
  assign _EVAL_1876 = _EVAL_913 ? _EVAL_1910 : 30'h0;
  assign _EVAL_980 = _EVAL_1301 | _EVAL_368;
  assign _EVAL_1752 = _EVAL_113 == 12'hc10;
  assign _EVAL_1103 = _EVAL_2006 & _EVAL_2378;
  assign _EVAL_503 = _EVAL_113 == 12'h32a;
  assign _EVAL_990 = ~_EVAL_699;
  assign _EVAL_914 = _EVAL_113 == 12'h3b1;
  assign _EVAL_1455 = _EVAL_1997 ? _EVAL_2490 : {{2'd0}, _EVAL_1813};
  assign _EVAL_326 = _EVAL_1248 | _EVAL_763;
  assign _EVAL_81 = _EVAL_617;
  assign _EVAL_1284 = _EVAL_402[7];
  assign _EVAL_1003 = _EVAL_1584 | _EVAL_2265;
  assign _EVAL_748 = ~_EVAL_20;
  assign _EVAL_942 = ~_EVAL_130;
  assign _EVAL_1303 = _EVAL_1841 & _EVAL_244;
  assign _EVAL_152 = _EVAL_1075;
  assign _EVAL_2346 = _EVAL_1520 | _EVAL_1146;
  assign _EVAL_1550 = _EVAL_113 == 12'hc05;
  assign _EVAL_1714 = _EVAL_113 == 12'h340;
  assign _EVAL_1259 = _EVAL_2517 ? 5'h1f : _EVAL_1740;
  assign _EVAL_1366 = _EVAL_2386 ? 5'h4 : _EVAL_871;
  assign _EVAL_2114 = _EVAL_250 ? 5'h7 : _EVAL_1396;
  assign _EVAL_521 = _EVAL_2328[39:32];
  assign _EVAL_401 = _EVAL_1080 ? _EVAL_1155 : 30'h0;
  assign _EVAL_1105 = _EVAL_882 ? _EVAL_528 : 40'h0;
  assign _EVAL_44 = _EVAL_2173[31:0];
  assign _EVAL_2295 = _EVAL_113 == 12'hb9d;
  assign _EVAL_115 = _EVAL_834 | _EVAL_164;
  assign _EVAL_1240 = _EVAL_618[12];
  assign _EVAL_2516 = ~_EVAL_1836;
  assign _EVAL_2318 = {{71'd0}, _EVAL_696};
  assign _EVAL_452 = _EVAL_312[0];
  assign _EVAL_1963 = _EVAL_402[24];
  assign _EVAL_815 = _EVAL_1881 | _EVAL_933;
  assign _EVAL_105 = _EVAL_2262;
  assign _EVAL_16 = _EVAL_500;
  assign _EVAL_1293 = _EVAL_1465 ? _EVAL_1642 : _EVAL_1516;
  assign _EVAL_1389 = _EVAL_1065 ? _EVAL_505 : {{2'd0}, _EVAL_1155};
  assign _EVAL_2197 = _EVAL_2242 | _EVAL_1822;
  assign _EVAL_796 = _EVAL_291 ? _EVAL_974 : _EVAL_2272;
  assign _EVAL_1411 = _EVAL_1526 ? _EVAL_754 : 32'h0;
  assign _EVAL_672 = _EVAL_2490[2];
  assign _EVAL_642 = _EVAL_1035 | _EVAL_2400;
  assign _EVAL_1562 = {_EVAL_2430, 13'h0};
  assign _EVAL_1052 = _EVAL_113 == 12'h333;
  assign _EVAL_1039 = _EVAL_151 == 12'h320;
  assign _EVAL_1096 = ~_EVAL_2485;
  assign _EVAL_2322 = _EVAL_1306 & _EVAL_1717;
  assign _EVAL_398 = _EVAL_113 == 12'hc93;
  assign _EVAL_2447 = _EVAL_151 == 12'hb82;
  assign _EVAL_1644 = _EVAL_329 < 2'h3;
  assign _EVAL_1094 = ~_EVAL_1161;
  assign _EVAL_1907 = _EVAL_372 & _EVAL_1088;
  assign _EVAL_1286 = _EVAL_2320 ? _EVAL_214 : _EVAL_1306;
  assign _EVAL_2433 = _EVAL_113 == 12'h344;
  assign _EVAL_108 = {_EVAL_2272,_EVAL_2182};
  assign _EVAL_2335 = _EVAL_1677[30:0];
  assign _EVAL_1457 = _EVAL_1518 & _EVAL_204;
  assign _EVAL_755 = _EVAL_2320 ? {{1'd0}, _EVAL_1280} : _EVAL_392;
  assign _EVAL_576 = ~_EVAL_273;
  assign _EVAL_56 = _EVAL_280;
  assign _EVAL_235 = _EVAL_1043 | _EVAL_2046;
  assign _EVAL_420 = 2'h3 == _EVAL_1541 ? _EVAL_1967 : _EVAL_624;
  assign _EVAL_2440 = _EVAL_113 == 12'hc1e;
  assign _EVAL_2284 = _EVAL_2439 & _EVAL_945;
  assign _EVAL_881 = _EVAL_151 == 12'hf11;
  assign _EVAL_614 = ~_EVAL_235;
  assign _EVAL_246 = _EVAL_113 == 12'h32d;
  assign _EVAL_624 = 2'h2 == _EVAL_1541 ? _EVAL_2301 : _EVAL_866;
  assign _EVAL_931 = {_EVAL_149,_EVAL_183,_EVAL_72,_EVAL_129,_EVAL_184,_EVAL_127,_EVAL_174};
  assign _EVAL_1018 = _EVAL_819[1];
  assign _EVAL_1454 = ~_EVAL_408;
  assign _EVAL_1569 = _EVAL_113 == 12'h306;
  assign _EVAL_1520 = _EVAL_1063 | _EVAL_1042;
  assign _EVAL_1209 = _EVAL_909 ? _EVAL_280 : 32'h0;
  assign _EVAL_866 = 2'h1 == _EVAL_1541 ? _EVAL_949 : _EVAL_1075;
  assign _EVAL_2394 = ~_EVAL_1660;
  assign _EVAL_1945 = _EVAL_1444 | _EVAL_397;
  assign _EVAL_1957 = _EVAL_632 | _EVAL_348;
  assign _EVAL_1667 = &_EVAL_1716;
  assign _EVAL_24 = _EVAL_2297;
  assign _EVAL_98 = _EVAL_891;
  assign _EVAL_1825 = _EVAL_291 ? _EVAL_365 : _EVAL_507;
  assign _EVAL_158 = _EVAL_385;
  assign _EVAL_1679 = ~_EVAL_115;
  assign _EVAL_321 = _EVAL_1500 ? 2'h1 : 2'h3;
  assign _EVAL_610 = _EVAL_1303 & _EVAL_1698;
  assign _EVAL_2439 = 2'h2 == _EVAL_1541;
  assign _EVAL_2519 = _EVAL_528[39:32];
  assign _EVAL_1364 = _EVAL_1461 & _EVAL_1482;
  assign _EVAL_1740 = _EVAL_2339 ? 5'h1e : _EVAL_547;
  assign _EVAL_407 = _EVAL_1051 == 32'h10000000;
  assign _EVAL_2256 = _EVAL_861 & _EVAL_2292;
  assign _EVAL_1549 = _EVAL_113 == 12'hc90;
  assign _EVAL_2054 = {_EVAL_1910,_EVAL_835};
  assign _EVAL_451 = _EVAL_1109 | _EVAL_1706;
  assign _EVAL_2044 = _EVAL_113 == 12'hc8f;
  assign _EVAL_1998 = {_EVAL_811,2'h3};
  assign _EVAL_525 = _EVAL_2210 & _EVAL_1393;
  assign _EVAL_511 = 2'h1 == _EVAL_1541;
  assign _EVAL_441 = {_EVAL_151, 20'h0};
  assign _EVAL_176 = _EVAL_1828;
  assign _EVAL_875 = _EVAL_1041 ? _EVAL_1670 : {{57'd0}, _EVAL_1944};
  assign _EVAL_959 = _EVAL_1136 ? _EVAL_439 : 32'h0;
  assign _EVAL_1049 = {_EVAL_675,2'h3};
  assign _EVAL_2013 = _EVAL_2359 ? _EVAL_2315 : 32'h0;
  assign _EVAL_367 = _EVAL_318 | _EVAL_1379;
  assign _EVAL_369 = _EVAL_113 == 12'hf14;
  assign _EVAL_2079 = _EVAL_113 == 12'h353;
  assign _EVAL_2053 = _EVAL_1040[0];
  assign _EVAL_2162 = _EVAL_1551[27];
  assign _EVAL_1153 = {{71'd0}, _EVAL_1235};
  assign _EVAL_765 = _EVAL_2492 & 32'h1f;
  assign _EVAL_1721 = _EVAL_113 == 12'h3b2;
  assign _EVAL_1941 = {{63'd0}, _EVAL_1894};
  assign _EVAL_569 = _EVAL_113 == 12'hb8d;
  assign _EVAL_1731 = _EVAL_151 == 12'hc83;
  assign _EVAL_2105 = _EVAL_763 ? 4'hb : _EVAL_635;
  assign _EVAL_592 = {_EVAL_1032,2'h0,_EVAL_679,_EVAL_1229,_EVAL_1694,_EVAL_2521,_EVAL_911,_EVAL_2414};
  assign _EVAL_512 = _EVAL_402[0];
  assign _EVAL_89 = _EVAL_1738;
  assign _EVAL_2199 = _EVAL_1877 | _EVAL_1048;
  assign _EVAL_1949 = _EVAL_2333[30:0];
  assign _EVAL_1471 = _EVAL_113 == 12'hb05;
  assign _EVAL_2221 = _EVAL_2080 | _EVAL_637;
  assign _EVAL_1892 = _EVAL_2368 | _EVAL_828;
  assign _EVAL_1260 = _EVAL_1773[31:0];
  assign _EVAL_916 = _EVAL_1084 ? _EVAL_929 : 32'h0;
  assign _EVAL_22 = _EVAL_1463;
  assign _EVAL_1100 = {_EVAL_1086,_EVAL_920};
  assign _EVAL_612 = _EVAL_973 & _EVAL_2241;
  assign _EVAL_1554 = _EVAL_197 & _EVAL_490;
  assign _EVAL_563 = ~_EVAL_2174;
  assign _EVAL_1009 = _EVAL_1551[24];
  assign _EVAL_883 = _EVAL_113 == 12'hc11;
  assign _EVAL_2474 = _EVAL_1850 & _EVAL_244;
  assign _EVAL_2103 = _EVAL_402[26];
  assign _EVAL_430 = ~_EVAL_783;
  assign _EVAL_1288 = _EVAL_631 & _EVAL_753;
  assign _EVAL_2534 = _EVAL_1482 ? _EVAL_300 : {{1'd0}, _EVAL_1505};
  assign _EVAL_1588 = _EVAL_511 & _EVAL_2529;
  assign _EVAL_412 = _EVAL_113 == 12'h325;
  assign _EVAL_1146 = _EVAL_113 == 12'hc18;
  assign _EVAL_1417 = 2'h1 == _EVAL_1541 ? _EVAL_2465 : _EVAL_2425;
  assign _EVAL_1717 = _EVAL_1695 | _EVAL_1534;
  assign _EVAL_1143 = _EVAL_402[21];
  assign _EVAL_974 = _EVAL_1698 | _EVAL_2272;
  assign _EVAL_896 = _EVAL_1065 ? _EVAL_720 : {{27'd0}, _EVAL_1733};
  assign _EVAL_170 = _EVAL_1504;
  assign _EVAL_127 = _EVAL_2185;
  assign _EVAL_858 = _EVAL_2548 | _EVAL_1927;
  assign _EVAL_547 = _EVAL_2544 ? 5'h1d : _EVAL_967;
  assign _EVAL_1518 = ~_EVAL_861;
  assign _EVAL_2444 = _EVAL_1909[31:0];
  assign _EVAL_2263 = _EVAL_268 | _EVAL_2138;
  assign _EVAL_1346 = _EVAL_113 == 12'h329;
  assign _EVAL_2181 = _EVAL_1551[11];
  assign _EVAL_2496 = _EVAL_113 == 12'h3bf;
  assign _EVAL_2402 = _EVAL_1528 ? 2'h3 : 2'h2;
  assign _EVAL_1251 = _EVAL_2338 & _EVAL_576;
  assign _EVAL_466 = _EVAL_440 & _EVAL_2374;
  assign _EVAL_1404 = _EVAL_402[12];
  assign _EVAL_619 = _EVAL_577 | _EVAL_1669;
  assign _EVAL_2126 = {{2'd0}, _EVAL_2182};
  assign _EVAL_1479 = _EVAL_1832 | _EVAL_1648;
  assign _EVAL_920 = {_EVAL_524, 2'h0};
  assign _EVAL_92 = _EVAL_2082;
  assign _EVAL_823 = _EVAL_151[10];
  assign _EVAL_1593 = {_EVAL_2174,2'h0,_EVAL_395,_EVAL_1557,_EVAL_1227,_EVAL_313,_EVAL_238};
  assign _EVAL_1750 = _EVAL_972 | _EVAL_1604;
  assign _EVAL_1925 = _EVAL_2466 ? _EVAL_1616 : 32'h0;
  assign _EVAL_184 = _EVAL_905;
  assign _EVAL_273 = _EVAL_2391 | _EVAL_287;
  assign _EVAL_1992 = {_EVAL_2519,_EVAL_2490};
  assign _EVAL_1430 = _EVAL_113 == 12'hb90;
  assign _EVAL_917 = _EVAL_2451 & _EVAL_236;
  assign _EVAL_1753 = _EVAL_823 & _EVAL_373;
  assign _EVAL_776 = _EVAL_113 == 12'hc9b;
  assign _EVAL_168 = _EVAL_1977 | _EVAL_2279;
  assign _EVAL_2542 = _EVAL_298 | _EVAL_916;
  assign _EVAL_685 = _EVAL_2056 & 32'hffff0888;
  assign _EVAL_1929 = _EVAL_402[17];
  assign _EVAL_852 = _EVAL_681 | _EVAL_897;
  assign _EVAL_1447 = _EVAL_2059 | _EVAL_2318;
  assign _EVAL_1785 = _EVAL_2490[12];
  assign _EVAL_147 = _EVAL_1161;
  assign _EVAL_1384 = {{63'd0}, _EVAL_2243};
  assign _EVAL_1855 = _EVAL_2098 ? 5'h5 : _EVAL_1013;
  assign _EVAL_889 = _EVAL_2504 ? 5'h10 : _EVAL_1309;
  assign _EVAL_1465 = _EVAL_2320 | _EVAL_1076;
  assign _EVAL_1961 = 2'h2 == _EVAL_1541 ? _EVAL_385 : _EVAL_1405;
  assign _EVAL_1367 = _EVAL_113 == 12'hb09;
  assign _EVAL_1347 = _EVAL_113 == 12'h7a3;
  assign _EVAL_893 = _EVAL_1322 ? 2'h3 : 2'h0;
  assign _EVAL_342 = _EVAL_1988 | _EVAL_334;
  assign _EVAL_47 = _EVAL_2461;
  assign _EVAL_880 = _EVAL_113 == 12'hc80;
  assign _EVAL_2218 = _EVAL_291 ? _EVAL_1399 : _EVAL_2027;
  assign _EVAL_1460 = _EVAL_1658 | _EVAL_2276;
  assign _EVAL_975 = _EVAL_1912 ? _EVAL_521 : 8'h0;
  assign _EVAL_2165 = _EVAL_1562[3];
  assign _EVAL_1607 = _EVAL_769 & _EVAL_1698;
  assign _EVAL_778 = _EVAL_2182 > 2'h1;
  assign _EVAL_904 = _EVAL_441 & 32'h20400000;
  assign _EVAL_1718 = 2'h3 == _EVAL_1541 ? _EVAL_460 : _EVAL_1351;
  assign _EVAL_1818 = _EVAL_1034 | _EVAL_2326;
  assign _EVAL_1869 = _EVAL_721 & _EVAL_2323;
  assign _EVAL_205 = _EVAL_1306 ? _EVAL_2549 : _EVAL_1070;
  assign _EVAL_1429 = _EVAL_113 == 12'hb83;
  assign _EVAL_428 = _EVAL_2535[0];
  assign _EVAL_104 = _EVAL_1334;
  assign _EVAL_1942 = {{73'd0}, _EVAL_1876};
  assign _EVAL_1827 = _EVAL_291 ? _EVAL_1187 : _EVAL_2482;
  assign _EVAL_2202 = _EVAL_1141 | _EVAL_1830;
  assign _EVAL_250 = _EVAL_2535[7];
  assign _EVAL_798 = _EVAL_1628 | _EVAL_1169;
  assign _EVAL_1526 = _EVAL_151 == 12'h351;
  assign _EVAL_2504 = _EVAL_1551[16];
  assign _EVAL_1948 = _EVAL_113 == 12'hb92;
  assign _EVAL_1802 = _EVAL_1687 | _EVAL_1958;
  assign _EVAL_1332 = ~_EVAL_1187;
  assign _EVAL_1602 = _EVAL_1701 | _EVAL_2072;
  assign _EVAL_1066 = _EVAL_113 == 12'hb11;
  assign _EVAL_1693 = _EVAL_1198 | _EVAL_895;
  assign _EVAL_573 = _EVAL_1056 & _EVAL_2267;
  assign _EVAL_1758 = _EVAL_113 == 12'hb9f;
  assign _EVAL_2027 = _EVAL_2320 ? _EVAL_1399 : _EVAL_1534;
  assign _EVAL_902 = _EVAL_2009 | _EVAL_1090;
  assign _EVAL_1110 = _EVAL_1515 | _EVAL_1984;
  assign _EVAL_482 = _EVAL_1274 | _EVAL_2374;
  assign _EVAL_2414 = {_EVAL_1947,2'h0,_EVAL_1212,_EVAL_741,_EVAL_1867,_EVAL_1595,_EVAL_1064};
  assign _EVAL_1095 = _EVAL_2505 ? _EVAL_227 : 30'h0;
  assign _EVAL_314 = _EVAL_1750 | _EVAL_190;
  assign _EVAL_1245 = _EVAL_113 < 12'hc20;
  assign _EVAL_1600 = _EVAL_113 == 12'h337;
  assign _EVAL_1962 = _EVAL_151 == 12'hc04;
  assign _EVAL_233 = _EVAL_1215 & _EVAL_1096;
  assign _EVAL_1354 = _EVAL_587 | _EVAL_1529;
  assign _EVAL_582 = _EVAL_1551[22];
  assign _EVAL_674 = _EVAL_1790 | _EVAL_1806;
  assign _EVAL_2307 = &_EVAL_60;
  assign _EVAL_146 = ~_EVAL_2202;
  assign _EVAL_1887 = 8'h0;
  assign _EVAL_594 = _EVAL_2490 & 32'hf;
  assign _EVAL_199 = {{39'd0}, _EVAL_2445};
  assign _EVAL_1072 = _EVAL_2490[5];
  assign _EVAL_110 = _EVAL_1032;
  assign _EVAL_919 = _EVAL_1882 | _EVAL_737;
  assign _EVAL_717 = _EVAL_1893 | _EVAL_2397;
  assign _EVAL_2058 = {{30'd0}, _EVAL_321};
  assign _EVAL_440 = _EVAL_685 & _EVAL_2128;
  assign _EVAL_599 = _EVAL_230 ? 32'h1 : 32'h0;
  assign _EVAL_938 = _EVAL_781 | _EVAL_2196;
  assign _EVAL_1968 = _EVAL_1736 ? _EVAL_1038 : {{1'd0}, _EVAL_2342};
  assign _EVAL_2378 = _EVAL_395[0];
  assign _EVAL_311 = _EVAL_1739 | _EVAL_499;
  assign _EVAL_2179 = _EVAL_2272 | _EVAL_164;
  assign _EVAL_2363 = {4'h2,_EVAL_1686,14'h400,_EVAL_2191,_EVAL_671,2'h0,_EVAL_727,_EVAL_1940};
  assign _EVAL_348 = _EVAL_113 == 12'hb97;
  assign _EVAL_2404 = _EVAL_113 == 12'h3bb;
  assign _EVAL_821 = _EVAL_1983 ? _EVAL_535 : _EVAL_1262;
  assign _EVAL_1558 = _EVAL_2279 ? _EVAL_329 : _EVAL_1904;
  assign _EVAL_305 = _EVAL_687 ? 32'h4210324 : 32'h0;
  assign _EVAL_1905 = ~_EVAL_1662;
  assign _EVAL_112 = _EVAL_767;
  assign _EVAL_513 = _EVAL_113 == 12'hc0a;
  assign _EVAL_2405 = _EVAL_1177 ? 7'h7e : 7'h2;
  assign _EVAL_2442 = {_EVAL_540,_EVAL_2267};
  assign _EVAL_287 = _EVAL_2174 & _EVAL_1103;
  assign _EVAL_317 = _EVAL_1652 | _EVAL_1571;
  assign _EVAL_2153 = _EVAL_1335 | _EVAL_1347;
  assign _EVAL_1118 = _EVAL_1327[17];
  assign _EVAL_1202 = _EVAL_113 == 12'hb8a;
  assign _EVAL_1092 = _EVAL_1602 | _EVAL_2410;
  assign _EVAL_2184 = _EVAL_113 == 12'h300;
  assign _EVAL_2319 = _EVAL_1119 ? _EVAL_2028 : _EVAL_875;
  assign _EVAL_725 = _EVAL_1816 ? 5'h13 : _EVAL_1589;
  assign _EVAL_1841 = _EVAL_2210 & _EVAL_407;
  assign _EVAL_837 = {_EVAL_1782, 2'h0};
  assign _EVAL_240 = _EVAL_2074 | _EVAL_517;
  assign _EVAL_1041 = _EVAL_151 == 12'hb00;
  assign _EVAL_2454 = _EVAL_652 | _EVAL_867;
  assign _EVAL_1060 = _EVAL_1654 ? 5'h19 : _EVAL_2022;
  assign _EVAL_77 = _EVAL_825 | _EVAL_1607;
  assign _EVAL_459 = _EVAL_402[4];
  assign _EVAL_1927 = _EVAL_113 == 12'hb08;
  assign _EVAL_1997 = _EVAL_1485 & _EVAL_2127;
  assign _EVAL_1640 = _EVAL_1839 ? _EVAL_2099 : 32'h0;
  assign _EVAL_2436 = _EVAL_342 | _EVAL_1569;
  assign _EVAL_2120 = _EVAL_1808 | _EVAL_66;
  assign _EVAL_394 = _EVAL_113 >= 12'hc80;
  assign _EVAL_2487 = _EVAL_2490 & 32'h8000001f;
  assign _EVAL_1801 = _EVAL_113 == 12'h343;
  assign _EVAL_2336 = _EVAL_1019 ? _EVAL_293 : 32'h0;
  assign _EVAL_1210 = _EVAL_1732 | _EVAL_1143;
  assign _EVAL_710 = _EVAL_402[15];
  assign _EVAL_2046 = {{28'd0}, _EVAL_1913};
  assign _EVAL_236 = _EVAL_1150 & _EVAL_1395;
  assign _EVAL_1324 = _EVAL_523 | _EVAL_2131;
  assign _EVAL_2004 = _EVAL_2320 & _EVAL_1534;
  assign _EVAL_1778 = _EVAL_1759 | _EVAL_928;
  assign _EVAL_1386 = _EVAL_938 | _EVAL_2527;
  assign _EVAL_1807 = _EVAL_564[4:3];
  assign _EVAL_210 = {{73'd0}, _EVAL_403};
  assign _EVAL_2266 = _EVAL_1667 ? _EVAL_73 : 32'h0;
  assign _EVAL_116 = _EVAL_1556[31:0];
  assign _EVAL_2371 = _EVAL_1977 | _EVAL_102;
  assign _EVAL_2497 = {{63'd0}, _EVAL_1105};
  assign _EVAL_1482 = ~_EVAL_1537;
  assign _EVAL_298 = _EVAL_2478 | _EVAL_2016;
  assign _EVAL_1939 = _EVAL_394 & _EVAL_787;
  assign _EVAL_1874 = {_EVAL_2465,1'h0,1'h0,_EVAL_1620,_EVAL_1618,_EVAL_949,_EVAL_872};
  assign _EVAL_769 = _EVAL_2387 & _EVAL_2112;
  assign _EVAL_811 = _EVAL_384 & _EVAL_2435;
  assign _EVAL_2480 = _EVAL_1756 & _EVAL_1454;
  assign _EVAL_2160 = _EVAL_1332 | _EVAL_2058;
  assign _EVAL_2278 = _EVAL_402[9];
  assign _EVAL_2109 = ~_EVAL_2179;
  assign _EVAL_739 = {_EVAL_2251, 30'h0};
  assign _EVAL_1405 = 2'h1 == _EVAL_1541 ? _EVAL_1357 : _EVAL_2245;
  assign _EVAL_111 = _EVAL_1733[0];
  assign _EVAL_304 = _EVAL_1795 & _EVAL_835;
  assign _EVAL_232 = _EVAL_1860 | _EVAL_1448;
  assign _EVAL_1341 = _EVAL_2495 ? 5'h1b : _EVAL_1283;
  assign _EVAL_2015 = _EVAL_317 | _EVAL_771;
  assign _EVAL_1498 = _EVAL_2371 ? _EVAL_1976 : _EVAL_237;
  assign _EVAL_9 = _EVAL_1935;
  assign _EVAL_1348 = {{25'd0}, _EVAL_2405};
  assign _EVAL_2022 = _EVAL_1963 ? 5'h18 : _EVAL_283;
  assign _EVAL_2062 = _EVAL_113 == 12'hb03;
  assign _EVAL_1517 = _EVAL_1586 & _EVAL_45;
  assign _EVAL_1057 = _EVAL_1625 | _EVAL_353;
  assign _EVAL_560 = _EVAL_1439 + 34'h1;
  assign _EVAL_150 = _EVAL_1694;
  assign _EVAL_1933 = _EVAL_1112 ? 5'h3 : _EVAL_2114;
  assign _EVAL_2006 = ~_EVAL_1564;
  assign _EVAL_248 = _EVAL_1778 | _EVAL_692;
  assign _EVAL_6 = _EVAL_1920;
  assign _EVAL_768 = _EVAL_2280[7];
  assign _EVAL_215 = _EVAL_113 == 12'h326;
  assign _EVAL_1529 = _EVAL_113 == 12'hc09;
  assign _EVAL_2147 = _EVAL_343 | _EVAL_957;
  assign _EVAL_1833 = _EVAL_1029[63:6];
  assign _EVAL_1884 = _EVAL_625 | _EVAL_428;
  assign _EVAL_1381 = _EVAL_113 == 12'hb8f;
  assign _EVAL_830 = _EVAL_1246 | _EVAL_2484;
  assign _EVAL_2368 = _EVAL_1879 | _EVAL_530;
  assign _EVAL_2242 = {{71'd0}, _EVAL_935};
  assign _EVAL_1597 = _EVAL_1551[14];
  assign _EVAL_2265 = _EVAL_113 == 12'hc88;
  assign _EVAL_1407 = _EVAL_1689 ? _EVAL_629 : 32'h0;
  assign _EVAL_346 = _EVAL_113 == 12'h3bc;
  assign _EVAL_329 = _EVAL_1983 ? _EVAL_237 : _EVAL_1107;
  assign _EVAL_11 = _EVAL_1229;
  assign _EVAL_325 = _EVAL_1306 ? _EVAL_1565 : _EVAL_1187;
  assign _EVAL_2047 = _EVAL_113 == 12'h351;
  assign _EVAL_1991 = _EVAL_942 | 32'h1;
  assign _EVAL_1126 = _EVAL_1364 ? _EVAL_1369 : _EVAL_1439;
  assign _EVAL_568 = _EVAL_232 | _EVAL_670;
  assign _EVAL_1175 = 2'h2 == _EVAL_1541 ? _EVAL_617 : _EVAL_414;
  assign _EVAL_1990 = _EVAL_113 == 12'hb13;
  assign _EVAL_1664 = _EVAL_1062 + 58'h1;
  assign _EVAL_177 = _EVAL_679;
  assign _EVAL_734 = _EVAL_113 == 12'hc15;
  assign _EVAL_1860 = _EVAL_642 | _EVAL_1613;
  assign _EVAL_1073 = _EVAL_1069 ? 5'h14 : _EVAL_725;
  assign _EVAL_2137 = _EVAL_1306 ? _EVAL_893 : _EVAL_965;
  assign _EVAL_1783 = _EVAL_2024 ? _EVAL_1755 : {{1'd0}, _EVAL_498};
  assign _EVAL_129 = _EVAL_1534;
  assign _EVAL_156 = _EVAL_937;
  assign _EVAL_446 = _EVAL_1321 | _EVAL_1023;
  assign _EVAL_2457 = 2'h3 == _EVAL_1541 ? _EVAL_1878 : _EVAL_1175;
  assign _EVAL_2025 = _EVAL_2490 & 32'hfffffffd;
  assign _EVAL_2092 = _EVAL_113 == 12'h7b0;
  assign _EVAL_2423 = 2'h2 == _EVAL_1541 ? _EVAL_500 : _EVAL_333;
  assign _EVAL_474 = _EVAL_113 == 12'hb93;
  assign _EVAL_1116 = _EVAL_2371 ? _EVAL_1827 : _EVAL_1187;
  assign _EVAL_258 = _EVAL_113 == 12'hb9c;
  assign _EVAL_1015 = _EVAL_918 + 31'h1;
  assign _EVAL_185 = _EVAL_1867;
  assign _EVAL_124 = _EVAL_1734[31:0];
  assign _EVAL_1081 = _EVAL_1562[9];
  assign _EVAL_728 = _EVAL_1551[3];
  assign _EVAL_1901 = _EVAL_113 == 12'hc1d;
  assign _EVAL_585 = _EVAL_546 | _EVAL_246;
  assign _EVAL_13 = _EVAL_1525;
  assign _EVAL_169 = _EVAL_1357;
  assign _EVAL_1652 = _EVAL_322 | _EVAL_608;
  assign _EVAL_780 = _EVAL_1284 ? 4'h7 : _EVAL_2541;
  assign _EVAL_1037 = {{71'd0}, _EVAL_1140};
  assign _EVAL_874 = _EVAL_1916 | _EVAL_2130;
  assign _EVAL_1035 = _EVAL_1862 | _EVAL_880;
  assign _EVAL_1283 = _EVAL_2103 ? 5'h1a : _EVAL_1060;
  assign _EVAL_1768 = _EVAL_1872 | _EVAL_1630;
  assign _EVAL_402 = _EVAL_2537 ? _EVAL_466 : 32'h0;
  assign _EVAL_1645 = _EVAL_1329 | _EVAL_2181;
  assign _EVAL_1130 = ~_EVAL_1032;
  assign _EVAL_888 = _EVAL_1551[23];
  assign _EVAL_414 = 2'h1 == _EVAL_1541 ? _EVAL_872 : _EVAL_1463;
  assign _EVAL_443 = {4'h0,_EVAL_63,1'h0,2'h0,_EVAL_90,1'h0,2'h0,_EVAL_57,1'h0,2'h0};
  assign _EVAL_1627 = ~_EVAL_2073;
  assign _EVAL_447 = _EVAL_1597 ? 5'he : _EVAL_2477;
  assign _EVAL_1793 = _EVAL_1645 | _EVAL_728;
  assign _EVAL_1984 = _EVAL_113 == 12'hb8e;
  assign _EVAL_12 = _EVAL_949;
  assign _EVAL_1710 = _EVAL_713 & _EVAL_1157;
  assign _EVAL_1256 = _EVAL_113 == 12'hb9e;
  assign _EVAL_2327 = _EVAL_405 & _EVAL_430;
  assign _EVAL_238 = {_EVAL_2391,2'h0,_EVAL_312,_EVAL_795,_EVAL_2461,_EVAL_1383};
  assign _EVAL_42 = _EVAL_1155;
  assign _EVAL_1133 = ~_EVAL_1581;
  assign _EVAL_845 = _EVAL_882 ? _EVAL_1992 : {{33'd0}, _EVAL_2534};
  assign _EVAL_1926 = _EVAL_1519 & _EVAL_1468;
  assign _EVAL_506 = _EVAL_402[22];
  assign _EVAL_260 = _EVAL_537 | _EVAL_251;
  assign _EVAL_2390 = {_EVAL_2280,_EVAL_607};
  assign _EVAL_2549 = 32'h80000000 | _EVAL_1402;
  assign _EVAL_1737 = _EVAL_113 == 12'h3b3;
  assign _EVAL_2178 = _EVAL_1310 | _EVAL_553;
  assign _EVAL_437 = _EVAL_2124[63:6];
  assign _EVAL_1953 = _EVAL_1892 | _EVAL_1752;
  assign _EVAL_1851 = _EVAL_1525[0];
  assign _EVAL_963 = {_EVAL_18,_EVAL_135,_EVAL_141,_EVAL_126,_EVAL_120,_EVAL_84,_EVAL_49,_EVAL_88};
  assign _EVAL_878 = _EVAL_461[1];
  assign _EVAL_1481 = _EVAL_2328[31:0];
  assign _EVAL_1363 = _EVAL_694 | _EVAL_2055;
  assign _EVAL_885 = _EVAL_973 & _EVAL_1709;
  assign _EVAL_524 = _EVAL_531[4:0];
  assign _EVAL_792 = _EVAL_113 == 12'hc12;
  assign _EVAL_17 = _EVAL_2451;
  assign _EVAL_824 = 2'h3 == _EVAL_1541 ? _EVAL_647 : _EVAL_1961;
  assign _EVAL_853 = 2'h1 == _EVAL_1541 ? _EVAL_2163 : _EVAL_1113;
  assign _EVAL_973 = _EVAL_151 == 12'h3a1;
  assign _EVAL_871 = _EVAL_1880 ? 5'h1f : _EVAL_1729;
  assign _EVAL_2039 = {{71'd0}, _EVAL_1925};
  assign _EVAL_1107 = _EVAL_1753 ? _EVAL_965 : _EVAL_365;
  assign _EVAL_1535 = _EVAL_593 | _EVAL_2110;
  assign _EVAL_1121 = _EVAL_113 == 12'hb86;
  assign _EVAL_1002 = _EVAL_2393 & _EVAL_1266;
  assign _EVAL_2411 = _EVAL_113 == 12'hb98;
  assign _EVAL_1250 = _EVAL_113 == 12'h320;
  assign _EVAL_706 = _EVAL_747 | _EVAL_2344;
  assign _EVAL_1179 = _EVAL_2371 ? _EVAL_1592 : _EVAL_2329;
  assign _EVAL_763 = _EVAL_402[11];
  assign _EVAL_695 = {_EVAL_1001,_EVAL_1511,_EVAL_689,_EVAL_804,_EVAL_245,_EVAL_1761,_EVAL_2426,_EVAL_1514};
  assign _EVAL_2210 = _EVAL_134 == 3'h4;
  assign _EVAL_2041 = _EVAL_151 == 12'h323;
  assign _EVAL_1581 = _EVAL_665 | _EVAL_691;
  assign _EVAL_1042 = _EVAL_113 == 12'hb18;
  assign _EVAL_1287 = _EVAL_2481[1];
  assign _EVAL_997 = _EVAL_113 == 12'h328;
  assign _EVAL_907 = _EVAL_267 | _EVAL_1749;
  assign _EVAL_308 = _EVAL_1731 ? _EVAL_1810 : 8'h0;
  assign _EVAL_1690 = _EVAL_683 | _EVAL_723;
  assign _EVAL_1897 = _EVAL_973 & _EVAL_1130;
  assign _EVAL_1470 = _EVAL_113 == 12'hb0e;
  assign _EVAL_803 = _EVAL_113 == 12'hb85;
  assign _EVAL_476 = _EVAL_2468 | _EVAL_358;
  assign _EVAL_262 = _EVAL_1031 ? _EVAL_676 : 32'h0;
  assign _EVAL_2096 = _EVAL_113[11:10];
  assign _EVAL_131 = _EVAL_2521;
  assign _EVAL_2412 = _EVAL_2196 ? 5'hc : _EVAL_2150;
  assign _EVAL_1604 = _EVAL_402[5];
  assign _EVAL_1848 = _EVAL_697 | _EVAL_1256;
  assign _EVAL_1509 = _EVAL_113 == 12'h33e;
  assign _EVAL_909 = _EVAL_151 == 12'h301;
  assign _EVAL_1204 = _EVAL_1288 & _EVAL_1911;
  assign _EVAL_898 = 32'h0;
  assign _EVAL_48 = _EVAL_2177 | _EVAL_155;
  assign _EVAL_2091 = _EVAL_2126 + 4'h8;
  assign _EVAL_1798 = _EVAL_2277 ? _EVAL_2168 : _EVAL_1062;
  assign _EVAL_2503 = _EVAL_1947 | _EVAL_2325;
  assign _EVAL_1385 = _EVAL_2071 | _EVAL_1714;
  assign _EVAL_274 = _EVAL_1800 | _EVAL_1938;
  assign _EVAL_631 = _EVAL_380 & _EVAL_2272;
  assign _EVAL_332 = _EVAL_2361 & _EVAL_2272;
  assign _EVAL_2192 = _EVAL_151 == 12'h7b0;
  assign _EVAL_2232 = _EVAL_1753 ? _EVAL_2401 : _EVAL_1399;
  assign _EVAL_915 = _EVAL_1009 ? 5'h18 : _EVAL_1524;
  assign _EVAL_781 = _EVAL_2108 | _EVAL_817;
  assign _EVAL_2121 = _EVAL_2535[4];
  assign _EVAL_330 = _EVAL_204 ? 32'h3 : _EVAL_50;
  assign _EVAL_125 = _EVAL_1633;
  assign _EVAL_591 = _EVAL_800 | _EVAL_2132;
  assign _EVAL_1249 = _EVAL_113 == 12'hb06;
  assign _EVAL_577 = _EVAL_2032 | _EVAL_532;
  assign _EVAL_514 = _EVAL_2530 ? _EVAL_849 : 32'h0;
  assign _EVAL_713 = _EVAL_548 & _EVAL_2272;
  assign _EVAL_1058 = _EVAL_556 | _EVAL_1284;
  assign _EVAL_593 = _EVAL_825 | _EVAL_1905;
  assign _EVAL_760 = _EVAL_2279 ? _EVAL_821 : _EVAL_535;
  assign _EVAL_2045 = _EVAL_1929 ? 5'h11 : _EVAL_1792;
  assign _EVAL_1024 = _EVAL_113 == 12'hb9a;
  assign _EVAL_1970 = _EVAL_1311 ? _EVAL_2390 : _EVAL_845;
  assign _EVAL_2429 = {_EVAL_767,1'h0,1'h0,_EVAL_460,_EVAL_630,_EVAL_1967,_EVAL_1878};
  assign _EVAL_1124 = {_EVAL_2550,_EVAL_2248};
  assign _EVAL_1820 = _EVAL_113 == 12'hc85;
  assign _EVAL_1809 = _EVAL_1092 | _EVAL_565;
  assign _EVAL_1456 = _EVAL_2542 | _EVAL_2166;
  assign _EVAL_1732 = _EVAL_724 | _EVAL_506;
  assign _EVAL_1705 = _EVAL_1971 | _EVAL_2162;
  assign _EVAL_1635 = _EVAL_113 == 12'h3be;
  assign _EVAL_375 = _EVAL_2437 | _EVAL_381;
  assign _EVAL_78 = _EVAL_2301;
  assign _EVAL_1573 = _EVAL_485 & _EVAL_801;
  assign _EVAL_843 = _EVAL_113 == 12'h341;
  assign _EVAL_1749 = _EVAL_113 == 12'hc9c;
  assign _EVAL_136 = _EVAL_1206;
  assign _EVAL_351 = _EVAL_2279 ? _EVAL_2107 : _EVAL_192;
  assign _EVAL_2479 = _EVAL_113 == 12'hb8b;
  assign _EVAL_1392 = _EVAL_2320 ? _EVAL_2099 : _EVAL_531;
  assign _EVAL_1190 = {4'h2,_EVAL_282,14'h400,_EVAL_1478,1'h0,2'h0,_EVAL_1696,_EVAL_2429};
  assign _EVAL_575 = {{5'd0}, _EVAL_166};
  assign _EVAL_2028 = {_EVAL_2490,_EVAL_223};
  assign _EVAL_2113 = _EVAL_2393 ? _EVAL_2262 : 30'h0;
  assign _EVAL_59 = _EVAL_799;
  assign _EVAL_1308 = _EVAL_1690 | _EVAL_1452;
  assign _EVAL_721 = _EVAL_564[1];
  assign _EVAL_1340 = {{95'd0}, _EVAL_975};
  assign _EVAL_2466 = _EVAL_151 == 12'hc82;
  assign _EVAL_1583 = _EVAL_1090 ? 5'h5 : _EVAL_216;
  assign _EVAL_163 = _EVAL_1910;
  assign _EVAL_181 = _EVAL_1496 & _EVAL_1698;
  assign _EVAL_682 = _EVAL_1670[63:6];
  assign _EVAL_1016 = _EVAL_113 == 12'hb0d;
  assign _EVAL_1678 = _EVAL_714 | _EVAL_1654;
  assign _EVAL_1859 = _EVAL_2183 | _EVAL_1411;
  assign _EVAL_1531 = _EVAL_543 | _EVAL_2098;
  assign _EVAL_584 = _EVAL_113 == 12'hc1b;
  assign _EVAL_1566 = _EVAL_663 ? _EVAL_2490 : {{30'd0}, _EVAL_1541};
  assign _EVAL_958 = _EVAL_113 == 12'h335;
  assign _EVAL_2415 = _EVAL_441 & 32'h10100000;
  assign _EVAL_2501 = _EVAL_2093 & _EVAL_1245;
  assign _EVAL_1872 = _EVAL_807 | _EVAL_1683;
  assign _EVAL_639 = _EVAL_1416[63:32];
  assign _EVAL_2138 = _EVAL_1959 & 32'hfffffffe;
  assign _EVAL_160 = _EVAL_2418;
  assign _EVAL_1402 = {{30'd0}, _EVAL_2402};
  assign _EVAL_556 = _EVAL_326 | _EVAL_700;
  assign _EVAL_2328 = {_EVAL_1817,_EVAL_498};
  assign _EVAL_109 = _EVAL_1326;
  assign _EVAL_1662 = _EVAL_1308 | _EVAL_844;
  assign _EVAL_537 = _EVAL_1659 | _EVAL_958;
  assign _EVAL_1862 = _EVAL_1956 | _EVAL_1440;
  assign _EVAL_1010 = _EVAL_113 == 12'hc04;
  assign _EVAL_52 = _EVAL_207[31:0];
  assign _EVAL_2243 = _EVAL_1930 ? _EVAL_528 : 40'h0;
  assign _EVAL_553 = _EVAL_113 == 12'hc13;
  assign _EVAL_187 = _EVAL_2178 | _EVAL_474;
  assign _EVAL_1836 = _EVAL_1796 | _EVAL_417;
  assign _EVAL_596 = _EVAL_728 ? 5'h3 : _EVAL_2469;
  assign _EVAL_1533 = _EVAL_2511[30:0];
  assign _EVAL_1904 = _EVAL_2371 ? _EVAL_2347 : _EVAL_2182;
  assign _EVAL_1999 = _EVAL_2320 ? _EVAL_205 : _EVAL_1070;
  assign _EVAL_1230 = _EVAL_1371 | _EVAL_1009;
  assign _EVAL_1850 = _EVAL_2086 | _EVAL_459;
  assign _EVAL_2528 = _EVAL_113 == 12'hb17;
  assign _EVAL_1043 = ~_EVAL_2490;
  assign _EVAL_1484 = _EVAL_531[7:0];
  assign _EVAL_249 = _EVAL_483 | _EVAL_514;
  assign _EVAL_1327 = {{71'd0}, _EVAL_2490};
  assign _EVAL_945 = _EVAL_558 | _EVAL_2272;
  assign _EVAL_279 = _EVAL_113 == 12'hb1d;
  assign _EVAL_2249 = _EVAL_1312 | _EVAL_1906;
  assign _EVAL_1040 = _EVAL_1221 >> _EVAL_2182;
  assign _EVAL_1145 = _EVAL_204 ? 12'h800 : 12'h808;
  assign _EVAL_1613 = _EVAL_113 == 12'h3a0;
  assign _EVAL_2536 = 2'h2 == _EVAL_1541 ? _EVAL_417 : _EVAL_1228;
  assign _EVAL_1349 = _EVAL_1768 | _EVAL_327;
  assign _EVAL_2551 = _EVAL_1742 | _EVAL_2496;
  assign _EVAL_2064 = _EVAL_151 == 12'h7c1;
  assign _EVAL_1452 = _EVAL_113 == 12'hf11;
  assign _EVAL_2376 = _EVAL_2206 | _EVAL_1290;
  assign _EVAL_2305 = _EVAL_1186 | _EVAL_73;
  assign _EVAL_1395 = _EVAL_1738[0];
  assign _EVAL_1164 = _EVAL_291 ? _EVAL_1306 : _EVAL_1286;
  assign _EVAL_1700 = {_EVAL_2048,2'h3};
  assign _EVAL_1564 = _EVAL_395[1];
  assign _EVAL_268 = _EVAL_2490 & 32'h1;
  assign _EVAL_675 = _EVAL_2054 & _EVAL_2282;
  assign _EVAL_37 = &_EVAL_2096;
  assign _EVAL_1687 = _EVAL_815 | _EVAL_539;
  assign _EVAL_1022 = _EVAL_568 | _EVAL_1873;
  assign _EVAL_191 = _EVAL_402[19];
  assign _EVAL_541 = _EVAL_1208 | _EVAL_2260;
  assign _EVAL_1418 = _EVAL_1328 | _EVAL_2358;
  assign _EVAL_1720 = _EVAL_113 == 12'hc0c;
  assign _EVAL_2276 = _EVAL_113 == 12'h305;
  assign _EVAL_819 = _EVAL_1574[7:0];
  assign _EVAL_1342 = _EVAL_113 == 12'h332;
  assign _EVAL_2548 = _EVAL_1995 | _EVAL_997;
  assign _EVAL_850 = _EVAL_1378 | _EVAL_2195;
  assign _EVAL_2032 = _EVAL_480 | _EVAL_199;
  assign _EVAL_928 = _EVAL_113 == 12'hb91;
  assign _EVAL_208 = _EVAL_113 == 12'hb0c;
  assign _EVAL_362 = {_EVAL_1326,1'h0,1'h0,_EVAL_1300,_EVAL_500,_EVAL_2301,_EVAL_617};
  assign _EVAL_918 = {_EVAL_1813,_EVAL_212};
  assign _EVAL_2251 = _EVAL_1380 & _EVAL_1306;
  assign _EVAL_2089 = _EVAL_1983 ? _EVAL_1025 : _EVAL_400;
  assign _EVAL_2541 = _EVAL_2278 ? 4'h9 : _EVAL_1483;
  assign _EVAL_1830 = _EVAL_1503 & _EVAL_1178;
  assign _EVAL_1068 = _EVAL_1817 + 34'h1;
  assign _EVAL_486 = _EVAL_113 == 12'hc86;
  assign _EVAL_1712 = _EVAL_1032 | _EVAL_598;
  assign _EVAL_2468 = _EVAL_2294 | _EVAL_2140;
  assign _EVAL_200 = _EVAL_113 == 12'hc95;
  assign _EVAL_1767 = _EVAL_1884 | _EVAL_2121;
  assign _EVAL_2017 = _EVAL_1787[2];
  assign _EVAL_2189 = _EVAL_2270 | _EVAL_1316;
  assign _EVAL_863 = _EVAL_2283 | _EVAL_2377;
  assign _EVAL_2471 = _EVAL_1447 | _EVAL_1037;
  assign _EVAL_190 = _EVAL_402[8];
  assign _EVAL_726 = _EVAL_1771 & _EVAL_712;
  assign _EVAL_1958 = _EVAL_113 == 12'hc1c;
  assign _EVAL_1877 = _EVAL_2547 | _EVAL_189;
  assign _EVAL_483 = _EVAL_451 | _EVAL_1765;
  assign _EVAL_270 = _EVAL_679[0];
  assign _EVAL_2244 = _EVAL_2214 | _EVAL_1336;
  assign _EVAL_2132 = _EVAL_113 == 12'h33a;
  assign _EVAL_736 = _EVAL_113 == 12'hc94;
  assign _EVAL_1894 = _EVAL_701 ? _EVAL_2328 : 40'h0;
  assign _EVAL_450 = _EVAL_2174 | _EVAL_917;
  assign _EVAL_1064 = {_EVAL_665,2'h0,_EVAL_1525,_EVAL_1027,_EVAL_668,_EVAL_1920};
  assign _EVAL_2320 = _EVAL_2256 & _EVAL_924;
  assign _EVAL_2343 = _EVAL_151 == 12'h7a2;
  assign _EVAL_711 = _EVAL_354 | _EVAL_1189;
  assign _EVAL_2490 = _EVAL_2303 & _EVAL_490;
  assign _EVAL_809 = _EVAL_1518 & _EVAL_1028;
  assign _EVAL_2257 = _EVAL_1705 | _EVAL_444;
  assign _EVAL_1109 = _EVAL_1132 | _EVAL_1640;
  assign _EVAL_1119 = _EVAL_151 == 12'hb80;
  assign _EVAL_2164 = {_EVAL_735,_EVAL_2490};
  assign _EVAL_1691 = _EVAL_2493 & _EVAL_212;
  assign _EVAL_2369 = _EVAL_113 == 12'hc84;
  assign _EVAL_2463 = _EVAL_1373 | _EVAL_1863;
  assign _EVAL_1639 = _EVAL_1804 ? 5'h5 : _EVAL_495;
  assign _EVAL_7 = _EVAL_2422;
  assign _EVAL_2448 = _EVAL_209 ? _EVAL_2490 : {{2'd0}, _EVAL_227};
  assign _EVAL_1546 = _EVAL_710 ? 4'hf : _EVAL_2502;
  assign _EVAL_392 = {{1'd0}, _EVAL_1280};
  assign _EVAL_1560 = _EVAL_113 == 12'h33d;
  assign _EVAL_145 = _EVAL_2042;
  assign _EVAL_1445 = {_EVAL_359,_EVAL_452};
  assign _EVAL_2296 = _EVAL_929[0];
  assign _EVAL_2303 = _EVAL_364 | _EVAL_73;
  assign _EVAL_1316 = _EVAL_113 == 12'hb8c;
  assign _EVAL_320 = _EVAL_1349 | _EVAL_2226;
  assign _EVAL_225 = 2'h2 == _EVAL_1541 ? _EVAL_2075 : _EVAL_484;
  assign _EVAL_426 = _EVAL_1315 | _EVAL_2307;
  assign _EVAL_408 = _EVAL_1922[30:0];
  assign _EVAL_95 = _EVAL_2075;
  assign _EVAL_2417 = _EVAL_424 & _EVAL_2272;
  assign _EVAL_2267 = _EVAL_461[0];
  assign _EVAL_999 = _EVAL_151 == 12'h3b4;
  assign _EVAL_2527 = _EVAL_2535[11];
  assign _EVAL_2339 = _EVAL_1551[30];
  assign _EVAL_2170 = _EVAL_704 ? 5'hc : _EVAL_1764;
  assign _EVAL_429 = _EVAL_2442 + 31'h1;
  assign _EVAL_1854 = _EVAL_1551[28];
  assign _EVAL_712 = _EVAL_2409 | _EVAL_2272;
  assign _EVAL_652 = _EVAL_2033 | _EVAL_346;
  assign _EVAL_315 = _EVAL_2061 ? _EVAL_2490 : {{2'd0}, _EVAL_2418};
  assign _EVAL_1374 = _EVAL_1562[8];
  assign _EVAL_431 = _EVAL_2253 | _EVAL_947;
  assign _EVAL_1670 = {_EVAL_2029,_EVAL_2490};
  assign _EVAL_783 = _EVAL_2085[30:0];
  assign _EVAL_1170 = _EVAL_1923 ? 5'h19 : _EVAL_915;
  assign _EVAL_1137 = {{5'd0}, _EVAL_121};
  assign _EVAL_2460 = _EVAL_619 | _EVAL_1748;
  assign _EVAL_2392 = _EVAL_2371 ? _EVAL_2543 : _EVAL_2315;
  assign _EVAL_2514 = _EVAL_113 == 12'h338;
  assign _EVAL_1701 = _EVAL_465 | _EVAL_1202;
  assign _EVAL_504 = _EVAL_676 >> _EVAL_1776;
  assign _EVAL_405 = {_EVAL_2418,_EVAL_1851};
  assign _EVAL_1568 = _EVAL_1017 | _EVAL_2500;
  assign _EVAL_1839 = _EVAL_151 == 12'h342;
  assign _EVAL_1816 = _EVAL_1551[19];
  assign _EVAL_293 = {_EVAL_1161,2'h0,_EVAL_461,_EVAL_2422,_EVAL_1955,_EVAL_1504,_EVAL_1883,_EVAL_1593};
  assign _EVAL_2003 = _EVAL_2490[8:7];
  assign _EVAL_967 = _EVAL_1854 ? 5'h1c : _EVAL_1934;
  assign _EVAL_2469 = _EVAL_2456 ? 5'h7 : _EVAL_2134;
  assign _EVAL_1950 = ~_EVAL_2285;
  assign _EVAL_214 = _EVAL_1306 ? 1'h0 : _EVAL_1306;
  assign _EVAL_1265 = _EVAL_1002 ? _EVAL_2490 : {{2'd0}, _EVAL_2262};
  assign _EVAL_1556 = {_EVAL_2327,2'h3};
  assign _EVAL_2180 = _EVAL_1962 ? _EVAL_2328 : 40'h0;
  assign _EVAL_355 = _EVAL_2451 | _EVAL_1345;
  assign _EVAL_2169 = _EVAL_2210 & _EVAL_337;
  assign _EVAL_1313 = _EVAL_291 ? {{1'd0}, _EVAL_1280} : _EVAL_755;
  assign _EVAL_791 = _EVAL_113 == 12'hc8c;
  assign _EVAL_165 = _EVAL_1959;
  assign _EVAL_26 = _EVAL_312;
  assign _EVAL_82 = _EVAL_722;
  assign _EVAL_1940 = {_EVAL_2349,1'h0,1'h0,_EVAL_1718,_EVAL_2171,_EVAL_420,_EVAL_2457};
  assign _EVAL_469 = _EVAL_582 ? 5'h16 : _EVAL_2208;
  assign _EVAL_2350 = _EVAL_847 | _EVAL_350;
  assign _EVAL_1401 = _EVAL_1575 & _EVAL_1851;
  assign _EVAL_2112 = _EVAL_113[7];
  assign _EVAL_2347 = _EVAL_291 ? _EVAL_2035 : _EVAL_1007;
  assign _EVAL_271 = _EVAL_113 == 12'h7a0;
  assign _EVAL_2144 = _EVAL_1203 ? 4'hd : _EVAL_2077;
  assign _EVAL_286 = _EVAL_2274 | _EVAL_2145;
  assign _EVAL_1931 = _EVAL_332 | _EVAL_1964;
  assign _EVAL_1458 = _EVAL_1230 | _EVAL_888;
  assign _EVAL_161 = _EVAL_2279 ? _EVAL_2498 : _EVAL_1594;
  assign _EVAL_691 = _EVAL_1947 & _EVAL_1691;
  assign _EVAL_445 = _EVAL_715 | _EVAL_1737;
  assign _EVAL_1771 = 2'h0 == _EVAL_1541;
  assign _EVAL_602 = _EVAL_2165 ? 5'h3 : _EVAL_1273;
  assign _EVAL_381 = _EVAL_954 ? _EVAL_1870 : 32'h0;
  assign _EVAL_122 = _EVAL_1213;
  assign _EVAL_64 = _EVAL_525 ? {{28'd0}, _EVAL_1599} : _EVAL_330;
  assign _EVAL_1274 = ~_EVAL_440;
  assign _EVAL_2014 = _EVAL_876 | _EVAL_2339;
  assign _EVAL_1880 = _EVAL_402[31];
  assign _EVAL_1350 = _EVAL_1131 & _EVAL_2024;
  assign _EVAL_2122 = _EVAL_320 | _EVAL_654;
  assign _EVAL_2020 = _EVAL_2119 & _EVAL_1803;
  assign _EVAL_955 = {{73'd0}, _EVAL_1095};
  assign _EVAL_1169 = _EVAL_2246 ? _EVAL_2363 : 32'h0;
  assign _EVAL_651 = _EVAL_1386 | _EVAL_1112;
  assign _EVAL_1235 = _EVAL_2063 ? _EVAL_1334 : 32'h0;
  assign _EVAL_189 = _EVAL_1562[0];
  assign _EVAL_1745 = _EVAL_113 == 12'h301;
  assign _EVAL_380 = _EVAL_1554[27];
  assign _EVAL_1028 = _EVAL_1484 == 8'he;
  assign _EVAL_1051 = _EVAL_441 & 32'h30000000;
  assign _EVAL_621 = _EVAL_1531 | _EVAL_2416;
  assign _EVAL_76 = _EVAL_370;
  assign _EVAL_382 = _EVAL_990 & _EVAL_270;
  assign _EVAL_65 = _EVAL_313;
  assign _EVAL_2250 = _EVAL_1423 | _EVAL_2396;
  assign _EVAL_1659 = _EVAL_1192 | _EVAL_736;
  assign _EVAL_1228 = 2'h1 == _EVAL_1541 ? _EVAL_985 : _EVAL_1796;
  assign _EVAL_2280 = _EVAL_2490[7:0];
  assign _EVAL_966 = {_EVAL_136,_EVAL_156,_EVAL_60,_EVAL_176,_EVAL_31,_EVAL_125,_EVAL_55,_EVAL_117,_EVAL_931};
  assign _EVAL_1030 = _EVAL_1081 ? 5'h9 : _EVAL_2198;
  assign _EVAL_1279 = _EVAL_1065 ? _EVAL_2319 : {{57'd0}, _EVAL_1944};
  assign _EVAL_604 = _EVAL_1041 ? _EVAL_1124 : 64'h0;
  assign _EVAL_732 = _EVAL_1251 ? _EVAL_2490 : {{2'd0}, _EVAL_359};
  assign _EVAL_29 = _EVAL_1027;
  assign _EVAL_1821 = _EVAL_1422 | _EVAL_1527;
  assign _EVAL_981 = _EVAL_113 == 12'hc8e;
  assign _EVAL_472 = _EVAL_2463 | _EVAL_1153;
  assign _EVAL_861 = _EVAL_531[31];
  assign _EVAL_1380 = _EVAL_748 & _EVAL_66;
  assign _EVAL_865 = {{63'd0}, _EVAL_2180};
  assign _EVAL_277 = _EVAL_291 ? _EVAL_1534 : _EVAL_2004;
  assign _EVAL_1183 = _EVAL_1540 | _EVAL_2039;
  assign _EVAL_1421 = ~_EVAL_1712;
  assign _EVAL_1215 = _EVAL_234[6];
  assign _EVAL_1111 = _EVAL_1255 | _EVAL_279;
  assign _EVAL_1589 = _EVAL_2060 ? 5'h12 : _EVAL_661;
  assign _EVAL_1114 = _EVAL_2320 ? _EVAL_2329 : _EVAL_1565;
  assign _EVAL_403 = _EVAL_999 ? _EVAL_2418 : 30'h0;
  assign _EVAL_1790 = _EVAL_2052 | _EVAL_1801;
  assign _EVAL_2135 = _EVAL_1689 ? _EVAL_810 : 32'h0;
  assign _EVAL_356 = _EVAL_113 == 12'hb94;
  assign _EVAL_1493 = _EVAL_113 == 12'hb0f;
  assign _EVAL_2292 = _EVAL_531[30];
  assign _EVAL_2193 = ~_EVAL_2102;
  assign _EVAL_744 = _EVAL_1760 | _EVAL_2432;
  assign _EVAL_323 = _EVAL_113 == 12'hc99;
  assign _EVAL_1254 = _EVAL_1936 | _EVAL_1553;
  assign _EVAL_2520 = _EVAL_650 | _EVAL_2495;
  assign _EVAL_418 = _EVAL_233 ? _EVAL_572 : _EVAL_2550;
  assign _EVAL_1142 = _EVAL_113 == 12'hc9e;
  assign _EVAL_1 = _EVAL_1124[31:0];
  assign _EVAL_810 = {4'h2,_EVAL_2366,14'h400,_EVAL_2075,_EVAL_417,2'h0,_EVAL_2082,_EVAL_362};
  assign _EVAL_2060 = _EVAL_1551[18];
  assign _EVAL_1764 = _EVAL_2181 ? 5'hb : _EVAL_596;
  assign _EVAL_930 = _EVAL_428 ? 5'h0 : _EVAL_555;
  assign _EVAL_494 = |_EVAL_440;
  assign _EVAL_251 = _EVAL_113 == 12'hb15;
  assign _EVAL_1808 = _EVAL_550 | _EVAL_2371;
  assign _EVAL_1444 = _EVAL_852 | _EVAL_1501;
  assign _EVAL_2397 = _EVAL_113 == 12'hc89;
  assign _EVAL_779 = _EVAL_113 == 12'h7b1;
  assign _EVAL_697 = _EVAL_2147 | _EVAL_2440;
  assign _EVAL_1489 = _EVAL_113 == 12'h3b6;
  assign _EVAL_2124 = {_EVAL_2490,_EVAL_1490};
  assign _EVAL_361 = _EVAL_2513 | _EVAL_1816;
  assign _EVAL_2034 = _EVAL_113 == 12'hc06;
  assign _EVAL_438 = _EVAL_2084[30:0];
  assign _EVAL_2143 = _EVAL_113 == 12'hb89;
  assign _EVAL_2452 = _EVAL_121 | _EVAL_2371;
  assign _EVAL_1191 = _EVAL_113 == 12'hb07;
  assign _EVAL_1838 = _EVAL_1945 | _EVAL_2062;
  assign _EVAL_1637 = _EVAL_1005 | _EVAL_2268;
  assign _EVAL_1069 = _EVAL_1551[20];
  assign _EVAL_2133 = _EVAL_2390[39:6];
  assign _EVAL_288 = &_EVAL_125;
  assign _EVAL_2055 = _EVAL_113 == 12'h32c;
  assign _EVAL_471 = _EVAL_113 == 12'h7a1;
  assign _EVAL_543 = _EVAL_2350 | _EVAL_1824;
  assign _EVAL_1425 = _EVAL_2371 ? _EVAL_796 : _EVAL_2272;
  assign _EVAL_2478 = _EVAL_1993 | _EVAL_1209;
  assign _EVAL_1883 = {_EVAL_2451,2'h0,_EVAL_1738,_EVAL_891,_EVAL_1788,_EVAL_1849};
  assign _EVAL_1857 = ~_EVAL_2335;
  assign _EVAL_851 = _EVAL_113 == 12'h3b4;
  assign _EVAL_172 = _EVAL_1231;
  assign _EVAL_1782 = _EVAL_929[31:2];
  assign _EVAL_1822 = _EVAL_1702 ? _EVAL_2476 : 103'h0;
  assign _EVAL_2345 = _EVAL_1065 ? _EVAL_1970 : {{33'd0}, _EVAL_2534};
  assign _EVAL_571 = _EVAL_2122 | _EVAL_1600;
  assign _EVAL_2223 = {{73'd0}, _EVAL_1046};
  assign _EVAL_684 = _EVAL_1210 | _EVAL_1924;
  assign _EVAL_2093 = _EVAL_113 >= 12'hc00;
  assign _EVAL_995 = _EVAL_2244 | _EVAL_569;
  assign _EVAL_1122 = {{73'd0}, _EVAL_655};
  assign _EVAL_1309 = _EVAL_481 ? 5'hf : _EVAL_447;
  assign _EVAL_175 = 1'h0;
  assign _EVAL_2217 = _EVAL_113 == 12'h3b7;
  assign _EVAL_2488 = _EVAL_1551[17];
  assign _EVAL_956 = _EVAL_2371 ? _EVAL_1969 : _EVAL_1978;
  assign _EVAL_216 = _EVAL_2271 ? 5'h8 : _EVAL_930;
  assign _EVAL_552 = {{71'd0}, _EVAL_413};
  assign _EVAL_1536 = _EVAL_2444 + _EVAL_943;
  assign _EVAL_183 = _EVAL_793;
  assign _EVAL_2029 = _EVAL_1124[63:32];
  assign _EVAL_3 = _EVAL_795;
  assign _EVAL_1787 = _EVAL_1888[7:0];
  assign _EVAL_1359 = _EVAL_1048 ? 5'h4 : _EVAL_1259;
  assign _EVAL_1063 = _EVAL_1275 | _EVAL_2514;
  assign _EVAL_1378 = _EVAL_367 | _EVAL_1122;
  assign _EVAL_2087 = _EVAL_134 == 3'h5;
  assign _EVAL_1599 = _EVAL_2091[3:0];
  assign _EVAL_555 = _EVAL_2121 ? 5'h4 : _EVAL_253;
  assign _EVAL_2508 = _EVAL_2376 | _EVAL_1381;
  assign _EVAL_1969 = _EVAL_291 ? _EVAL_1612 : _EVAL_1978;
  assign _EVAL_1697 = _EVAL_189 ? 5'h0 : _EVAL_1359;
  assign _EVAL_625 = _EVAL_902 | _EVAL_2271;
  assign _EVAL_654 = _EVAL_113 == 12'hc96;
  assign _EVAL_670 = _EVAL_113 == 12'h3a2;
  assign _EVAL_1539 = _EVAL_1738[1];
  assign _EVAL_1741 = _EVAL_1567 ? _EVAL_1416 : 64'h0;
  assign _EVAL_1668 = _EVAL_375 | _EVAL_959;
  assign _EVAL_817 = _EVAL_2535[13];
  assign _EVAL_536 = _EVAL_2343 ? _EVAL_824 : 32'h0;
  assign _EVAL_546 = _EVAL_2189 | _EVAL_791;
  assign _EVAL_1315 = &_EVAL_176;
  assign _EVAL_2258 = _EVAL_2346 | _EVAL_2411;
  assign _EVAL_873 = _EVAL_2279 ? _EVAL_2089 : _EVAL_1025;
  assign _EVAL_531 = _EVAL_525 ? {{28'd0}, _EVAL_1599} : _EVAL_330;
  assign _EVAL_2416 = _EVAL_1551[8];
  assign _EVAL_197 = _EVAL_832 | _EVAL_73;
  assign _EVAL_40 = _EVAL_227;
  assign _EVAL_53 = _EVAL_1947;
  assign _EVAL_2134 = _EVAL_350 ? 5'h9 : _EVAL_2321;
  assign _EVAL_1689 = _EVAL_134[1];
  assign _EVAL_1248 = _EVAL_410 | _EVAL_1404;
  assign _EVAL_1896 = _EVAL_830 | _EVAL_1024;
  assign _EVAL_1485 = _EVAL_151 == 12'h3b5;
  assign _EVAL_281 = _EVAL_2535[9];
  assign _EVAL_204 = _EVAL_2210 & _EVAL_519;
  assign _EVAL_673 = _EVAL_297 | _EVAL_1052;
  assign _EVAL_1722 = _EVAL_134 == 3'h7;
  assign _EVAL_424 = _EVAL_1890[27];
  assign _EVAL_1698 = ~_EVAL_2272;
  assign _EVAL_1629 = _EVAL_1119 ? _EVAL_502 : 32'h0;
  assign _EVAL_1450 = _EVAL_1261[31:1];
  assign _EVAL_1177 = _EVAL_387[0];
  assign _EVAL_2314 = _EVAL_2041 ? _EVAL_1217 : 32'h0;
  assign _EVAL_2049 = _EVAL_1043 | 32'h1;
  assign _EVAL_2338 = _EVAL_151 == 12'h3b0;
  assign _EVAL_1601 = _EVAL_778 | _EVAL_775;
  assign _EVAL_477 = _EVAL_2258 | _EVAL_242;
  assign _EVAL_702 = _EVAL_1460 | _EVAL_2433;
  assign _EVAL_2434 = _EVAL_1050 ? 2'h3 : _EVAL_427;
  assign _EVAL_2188 = _EVAL_113 <= 12'h343;
  assign _EVAL_1912 = _EVAL_151 == 12'hb84;
  assign _EVAL_223 = _EVAL_1124[31:0];
  assign _EVAL_2359 = _EVAL_151 == 12'h343;
  assign _EVAL_1048 = _EVAL_1562[4];
  assign _EVAL_80 = _EVAL_665;
  assign _EVAL_322 = _EVAL_2197 | _EVAL_2313;
  assign _EVAL_2321 = _EVAL_1824 ? 5'h1 : _EVAL_1855;
  assign _EVAL_2513 = _EVAL_1818 | _EVAL_1069;
  assign _EVAL_802 = _EVAL_151 == 12'h300;
  assign _EVAL_951 = _EVAL_1510 | _EVAL_1384;
  assign _EVAL_1699 = _EVAL_113 == 12'hc97;
  assign _EVAL_856 = _EVAL_819[4:3];
  assign _EVAL_2208 = _EVAL_2326 ? 5'h15 : _EVAL_1073;
  assign _EVAL_97 = _EVAL_991[31:0];
  assign _EVAL_770 = _EVAL_1006 | _EVAL_865;
  assign _EVAL_1792 = _EVAL_2151 ? 5'h10 : {{1'd0}, _EVAL_1546};
  assign _EVAL_397 = _EVAL_113 == 12'h323;
  assign _EVAL_1636 = _EVAL_441 & 32'h20200000;
  assign _EVAL_2036 = 2'h1 == _EVAL_1541 ? _EVAL_1017 : _EVAL_962;
  assign _EVAL_2538 = _EVAL_187 | _EVAL_398;
  assign _EVAL_1952 = _EVAL_564[7];
  assign _EVAL_663 = _EVAL_151 == 12'h7a0;
  assign _EVAL_2253 = _EVAL_295 | _EVAL_1549;
  assign _EVAL_1882 = _EVAL_614 & 32'h1005;
  assign _EVAL_132 = _EVAL_1918;
  assign _EVAL_32 = _EVAL_820;
  assign _EVAL_1881 = _EVAL_657 | _EVAL_776;
  assign _EVAL_2191 = 2'h3 == _EVAL_1541 ? _EVAL_1478 : _EVAL_225;
  assign _EVAL_1794 = _EVAL_1018 & _EVAL_1410;
  assign _EVAL_1651 = _EVAL_1753 ? _EVAL_754 : _EVAL_439;
  assign _EVAL_1888 = _EVAL_2490[31:16];
  assign _EVAL_650 = _EVAL_1214 | _EVAL_730;
  assign _EVAL_1510 = _EVAL_2015 | _EVAL_2497;
  assign _EVAL_1393 = _EVAL_1168 == 32'h0;
  assign _EVAL_154 = _EVAL_1383;
  assign _EVAL_2171 = 2'h3 == _EVAL_1541 ? _EVAL_630 : _EVAL_2423;
  assign _EVAL_1144 = ~_EVAL_1072;
  assign _EVAL_1994 = _EVAL_1484 == 8'hc;
  assign _EVAL_306 = _EVAL_2490[1:0];
  assign _EVAL_676 = _EVAL_765;
  assign _EVAL_897 = _EVAL_113 == 12'hb00;
  assign _EVAL_926 = _EVAL_663 ? _EVAL_1541 : 2'h0;
  assign _EVAL_1724 = _EVAL_2037 | _EVAL_672;
  assign _EVAL_2018 = _EVAL_1065 ? _EVAL_533 : _EVAL_760;
  assign _EVAL_1239 = _EVAL_1311 ? _EVAL_1810 : 8'h0;
  assign _EVAL_353 = _EVAL_1562[11];
  assign _EVAL_968 = _EVAL_757 ? 5'h1 : _EVAL_1583;
  assign _EVAL_2110 = _EVAL_1708 & _EVAL_1719;
  assign _EVAL_1360 = _EVAL_1306 | _EVAL_515;
  assign _EVAL_626 = _EVAL_1406 ? 5'hc : _EVAL_1609;
  assign _EVAL_1410 = _EVAL_819[0];
  assign _EVAL_1013 = _EVAL_2416 ? 5'h8 : _EVAL_1954;
  assign _EVAL_2056 = {_EVAL_21,_EVAL_51,_EVAL_23,_EVAL_10,_EVAL_62,_EVAL_5,_EVAL_153,_EVAL_167,_EVAL_963,_EVAL_443};
  assign _EVAL_1461 = _EVAL_300[6];
  assign _EVAL_1192 = _EVAL_1254 | _EVAL_356;
  assign _EVAL_1080 = _EVAL_151 == 12'h3b7;
  assign _EVAL_1501 = _EVAL_113 == 12'hb02;
  assign _EVAL_1194 = _EVAL_1161 | _EVAL_1012;
  assign _EVAL_1716 = _EVAL_134[1:0];
  assign _EVAL_378 = _EVAL_191 ? 5'h13 : _EVAL_1200;
  assign _EVAL_1993 = _EVAL_798 | _EVAL_536;
  assign _EVAL_1157 = _EVAL_962 | _EVAL_936;
  assign _EVAL_947 = _EVAL_113 == 12'h331;
  assign _EVAL_634 = _EVAL_1983 ? _EVAL_2401 : _EVAL_2232;
  assign _EVAL_1373 = _EVAL_951 | _EVAL_473;
  assign _EVAL_2379 = {_EVAL_67,_EVAL_143,_EVAL_35,_EVAL_82,_EVAL_69,_EVAL_9,_EVAL_132,_EVAL_59};
  assign _EVAL_2084 = _EVAL_384 + 31'h1;
  assign _EVAL_870 = _EVAL_2447 ? _EVAL_1616 : 32'h0;
  assign _EVAL_2011 = _EVAL_2272 ? _EVAL_1145 : 12'h800;
  assign _EVAL_221 = _EVAL_113 == 12'h339;
  assign _EVAL_2 = _EVAL_2272;
  assign _EVAL_140 = _EVAL_1536[31:0];
  assign _EVAL_2239 = _EVAL_271 | _EVAL_471;
  assign _EVAL_2372 = _EVAL_921 | _EVAL_1121;
  assign _EVAL_1981 = _EVAL_1324 | _EVAL_2494;
  assign _EVAL_1800 = _EVAL_2372 | _EVAL_486;
  assign _EVAL_484 = 2'h1 == _EVAL_1541 ? _EVAL_820 : _EVAL_1344;
  assign _EVAL_1777 = _EVAL_1339 ? _EVAL_2490 : {{2'd0}, _EVAL_540};
  assign _EVAL_640 = _EVAL_2490 & 32'h80000003;
  assign _EVAL_1516 = _EVAL_2020 ? _EVAL_1100 : _EVAL_837;
  assign _EVAL_1658 = _EVAL_833 | _EVAL_2184;
  assign _EVAL_1914 = _EVAL_1065 ? _EVAL_315 : {{2'd0}, _EVAL_2418};
  assign _EVAL_646 = _EVAL_2065 | _EVAL_2219;
  assign _EVAL_991 = {_EVAL_2480,2'h3};
  assign _EVAL_1623 = ~_EVAL_1194;
  assign _EVAL_1047 = _EVAL_2280[4:3];
  assign _EVAL_1903 = _EVAL_1896 | _EVAL_658;
  assign _EVAL_244 = ~_EVAL_181;
  assign _EVAL_1628 = {{30'd0}, _EVAL_926};
  assign _EVAL_1765 = _EVAL_2192 ? _EVAL_695 : 32'h0;
  assign _EVAL_106 = _EVAL_1344;
  assign _EVAL_2310 = _EVAL_113 == 12'h3b8;
  assign _EVAL_1178 = _EVAL_113 <= 12'h143;
  assign _EVAL_1014 = _EVAL_2146 | _EVAL_412;
  assign _EVAL_895 = _EVAL_1562[1];
  assign _EVAL_622 = _EVAL_2135 | _EVAL_73;
  assign _EVAL_1924 = _EVAL_402[20];
  assign _EVAL_1415 = _EVAL_402[23];
  assign _EVAL_1503 = _EVAL_113 >= 12'h140;
  assign _EVAL_36 = _EVAL_196 | _EVAL_1627;
  assign _EVAL_1915 = _EVAL_1003 | _EVAL_1346;
  assign _EVAL_1497 = _EVAL_1924 ? 5'h14 : _EVAL_378;
  assign _EVAL_1492 = ~_EVAL_2049;
  assign _EVAL_1086 = _EVAL_929[31:7];
  assign _EVAL_1125 = _EVAL_113 == 12'hb99;
  assign _EVAL_1681 = _EVAL_701 ? _EVAL_2164 : {{33'd0}, _EVAL_1783};
  assign _EVAL_2489 = _EVAL_1693 | _EVAL_1804;
  assign _EVAL_400 = _EVAL_1753 ? _EVAL_1025 : 2'h0;
  assign _EVAL_2512 = _EVAL_2320 ? _EVAL_2315 : _EVAL_101;
  assign _EVAL_597 = _EVAL_2371 ? _EVAL_2382 : _EVAL_2099;
  assign _EVAL_1321 = _EVAL_989 | _EVAL_1597;
  assign _EVAL_1029 = {_EVAL_639,_EVAL_2490};
  assign _EVAL_1413 = _EVAL_1644 ? 1'h0 : _EVAL_937;
  assign _EVAL_1244 = _EVAL_265 | _EVAL_857;
  assign _EVAL_1123 = _EVAL_444 ? 5'h1a : _EVAL_1170;
  assign _EVAL_1091 = _EVAL_1866 | _EVAL_566;
  assign _EVAL_1661 = _EVAL_470 ? _EVAL_502 : 32'h0;
  assign _EVAL_1766 = 32'h0;
  assign _EVAL_2462 = _EVAL_1821 | _EVAL_792;
  assign _EVAL_2241 = ~_EVAL_665;
  assign _EVAL_1025 = _EVAL_2371 ? _EVAL_1825 : _EVAL_365;
  assign _EVAL_46 = _EVAL_647;
  assign _EVAL_54 = _EVAL_1788;
  assign _EVAL_2131 = _EVAL_113 == 12'hc07;
  assign _EVAL_507 = _EVAL_2320 ? _EVAL_365 : _EVAL_893;
  assign _EVAL_2102 = _EVAL_454 | _EVAL_598;
  assign _EVAL_2389 = _EVAL_1733[4];
  assign _EVAL_1561 = _EVAL_113 == 12'hc03;
  assign _EVAL_1132 = _EVAL_1668 | _EVAL_2013;
  assign _EVAL_989 = _EVAL_2467 | _EVAL_481;
  assign _EVAL_1490 = _EVAL_1416[31:0];
  assign _EVAL_1725 = {_EVAL_2425,1'h0,1'h0,_EVAL_1657,_EVAL_2331,_EVAL_1075,_EVAL_1463};
  assign _EVAL_179 = _EVAL_2391;
  assign _EVAL_349 = _EVAL_1891 & _EVAL_1698;
  assign _EVAL_465 = _EVAL_311 | _EVAL_513;
  assign _EVAL_1755 = _EVAL_498 + _EVAL_1563;
  assign _EVAL_243 = _EVAL_918 & _EVAL_2394;
  assign _EVAL_174 = _EVAL_2532;
  assign _EVAL_2330 = _EVAL_431 | _EVAL_1066;
  assign _EVAL_1442 = _EVAL_113 >= 12'h340;
  assign _EVAL_2190 = _EVAL_2021 | _EVAL_1036;
  assign _EVAL_523 = _EVAL_274 | _EVAL_1191;
  assign _EVAL_2061 = _EVAL_999 & _EVAL_1133;
  assign _EVAL_964 = ~_EVAL_1348;
  assign _EVAL_1567 = _EVAL_151 == 12'hb02;
  assign _EVAL_1298 = _EVAL_113 == 12'hb88;
  assign _EVAL_386 = _EVAL_904 == 32'h20000000;
  assign _EVAL_2177 = _EVAL_121 > 1'h0;
  assign _EVAL_2183 = _EVAL_1129 | _EVAL_1621;
  assign _EVAL_1989 = _EVAL_1698 ? _EVAL_893 : _EVAL_237;
  assign _EVAL_2377 = _EVAL_402[14];
  assign _EVAL_289 = _EVAL_1912 ? _EVAL_1441 : _EVAL_1681;
  assign _EVAL_1756 = {_EVAL_2262,_EVAL_2378};
  assign _EVAL_1776 = _EVAL_113[4:0];
  assign _EVAL_61 = _EVAL_1878;
  assign _EVAL_230 = _EVAL_151 == 12'hf12;
  assign _EVAL_2195 = {{73'd0}, _EVAL_2113};
  assign _EVAL_2357 = _EVAL_113 == 12'hc9d;
  assign _EVAL_857 = {{71'd0}, _EVAL_305};
  assign _EVAL_2291 = _EVAL_151 == 12'h3b3;
  assign _EVAL_2033 = _EVAL_2190 | _EVAL_2404;
  assign _EVAL_1916 = _EVAL_688 | _EVAL_809;
  assign _EVAL_1129 = _EVAL_249 | _EVAL_1762;
  assign _EVAL_935 = _EVAL_1859 | _EVAL_2117;
  assign _EVAL_256 = _EVAL_1065 ? _EVAL_289 : {{33'd0}, _EVAL_1783};
  assign _EVAL_2294 = _EVAL_2428 | _EVAL_1429;
  assign _EVAL_784 = _EVAL_674 | _EVAL_369;
  assign _EVAL_2511 = _EVAL_2054 + 31'h1;
  assign _EVAL_300 = _EVAL_1505 + _EVAL_575;
  assign _EVAL_1893 = _EVAL_1354 | _EVAL_2143;
  assign _EVAL_620 = _EVAL_1890[12];
  assign _EVAL_384 = {_EVAL_1155,_EVAL_270};
  assign _EVAL_75 = _EVAL_741;
  assign _EVAL_69 = _EVAL_1120;
  assign _EVAL_343 = _EVAL_1856 | _EVAL_1509;
  assign _EVAL_157 = _EVAL_417;
  assign _EVAL_1665 = _EVAL_113 == 12'h3b9;
  assign _EVAL_377 = _EVAL_419 ? _EVAL_2128 : 32'h0;
  assign _EVAL_957 = _EVAL_113 == 12'hb1e;
  assign _EVAL_2344 = _EVAL_402[18];
  assign _EVAL_1136 = _EVAL_151 == 12'h341;
  assign _EVAL_1977 = _EVAL_525 | _EVAL_204;
  assign _EVAL_527 = _EVAL_2279 ? _EVAL_1413 : _EVAL_937;
  assign _EVAL_1088 = _EVAL_2280[0];
  assign _EVAL_687 = _EVAL_151 == 12'hf13;
  assign _EVAL_1090 = _EVAL_2535[5];
  assign _EVAL_207 = {_EVAL_243,2'h3};
  assign _EVAL_2522 = _EVAL_545 | _EVAL_2058;
  assign _EVAL_2145 = _EVAL_113 == 12'h33f;
  assign _EVAL_924 = _EVAL_1270 | _EVAL_1994;
  assign _EVAL_653 = _EVAL_113 == 12'h3b0;
  assign _EVAL_590 = _EVAL_391[0];
  assign _EVAL_267 = _EVAL_1802 | _EVAL_258;
  assign _EVAL_724 = _EVAL_1634 | _EVAL_1415;
  assign _EVAL_1371 = _EVAL_2257 | _EVAL_1923;
  assign _EVAL_1083 = _EVAL_1567 ? _EVAL_1029 : {{57'd0}, _EVAL_1968};
  assign _EVAL_1379 = {{71'd0}, _EVAL_2399};
  assign _EVAL_2518 = _EVAL_1502 | _EVAL_2488;
  assign _EVAL_327 = _EVAL_113 == 12'hc16;
  assign _EVAL_2059 = _EVAL_1688 | _EVAL_2449;
  assign _EVAL_1351 = 2'h2 == _EVAL_1541 ? _EVAL_1300 : _EVAL_2524;
  assign _EVAL_1759 = _EVAL_2330 | _EVAL_883;
  assign _EVAL_2475 = _EVAL_1551[0];
  assign _EVAL_2485 = _EVAL_1733[0];
  assign _EVAL_1310 = _EVAL_673 | _EVAL_1990;
  assign _EVAL_2200 = _EVAL_913 & _EVAL_2193;
  assign _EVAL_1483 = _EVAL_1391 ? 4'h1 : _EVAL_2031;
  assign _EVAL_867 = _EVAL_113 == 12'h3bd;
  assign _EVAL_439 = ~_EVAL_1823;
  assign _EVAL_1944 = _EVAL_1096 ? _EVAL_234 : {{1'd0}, _EVAL_2248};
  assign _EVAL_39 = _EVAL_1300;
  assign _EVAL_860 = _EVAL_1485 ? _EVAL_1813 : 30'h0;
  assign _EVAL_2065 = _EVAL_2436 | _EVAL_899;
  assign _EVAL_1318 = _EVAL_1180 & _EVAL_2500;
  assign _EVAL_72 = _EVAL_743;
  assign _EVAL_2080 = _EVAL_1110 | _EVAL_981;
  assign _EVAL_708 = _EVAL_1022 | _EVAL_653;
  assign _EVAL_2073 = _EVAL_280[5];
  assign _EVAL_2154 = {{71'd0}, _EVAL_262};
  assign _EVAL_2219 = _EVAL_113 == 12'hc02;
  assign _EVAL_2270 = _EVAL_666 | _EVAL_1720;
  assign _EVAL_1328 = _EVAL_1797 | _EVAL_1880;
  assign _EVAL_485 = 2'h3 == _EVAL_1541;
  assign _EVAL_345 = _EVAL_706 | _EVAL_1929;
  assign _EVAL_1742 = _EVAL_2454 | _EVAL_1635;
  assign _EVAL_1160 = _EVAL_850 | _EVAL_955;
  assign _EVAL_1715 = _EVAL_1019 & _EVAL_1094;
  assign _EVAL_495 = _EVAL_1374 ? 5'h8 : _EVAL_1697;
  assign _EVAL_782 = ~_EVAL_2451;
  assign _EVAL_1835 = _EVAL_2320 ? _EVAL_2137 : _EVAL_965;
  assign _EVAL_490 = ~_EVAL_2266;
  assign _EVAL_1540 = _EVAL_2460 | _EVAL_616;
  assign _EVAL_705 = _EVAL_2490 & 32'hffff0888;
  assign _EVAL_2435 = ~_EVAL_438;
  assign _EVAL_737 = _EVAL_280 & 32'hffffeffa;
  assign _EVAL_1046 = _EVAL_2291 ? _EVAL_540 : 30'h0;
  assign _EVAL_389 = _EVAL_113 == 12'h304;
  assign _EVAL_60 = _EVAL_877;
  assign _EVAL_618 = _EVAL_2305 & _EVAL_490;
  assign _EVAL_360 = _EVAL_1091 | _EVAL_707;
  assign _EVAL_2063 = _EVAL_151 == 12'h324;
  assign _EVAL_1084 = _EVAL_151 == 12'h305;
  assign _EVAL_800 = _EVAL_2030 | _EVAL_323;
  assign _EVAL_364 = _EVAL_1689 ? _EVAL_103 : 32'h0;
  assign _EVAL_228 = _EVAL_2280[2];
  assign _EVAL_1335 = _EVAL_2239 | _EVAL_2365;
  assign _EVAL_419 = _EVAL_151 == 12'h304;
  assign _EVAL_2168 = _EVAL_1664[57:0];
  assign _EVAL_34 = _EVAL_1700[31:0];
  assign _EVAL_1211 = _EVAL_594 | _EVAL_2172;
  assign _EVAL_1921 = _EVAL_651 | _EVAL_250;
  assign _EVAL_1819 = _EVAL_2490[0];
  assign _EVAL_1625 = _EVAL_1285 | _EVAL_1406;
  assign _EVAL_159 = _EVAL_872;
  assign _EVAL_456 = _EVAL_113 == 12'hc0b;
  assign _EVAL_934 = 2'h2 == _EVAL_1541 ? _EVAL_1326 : _EVAL_1417;
  assign _EVAL_1551 = _EVAL_2322 ? _EVAL_2078 : 32'h0;
  assign _EVAL_542 = _EVAL_175 & _EVAL_36;
  assign _EVAL_2493 = ~_EVAL_1495;
  assign _EVAL_933 = _EVAL_113 == 12'h33c;
  assign _EVAL_516 = _EVAL_2452 | _EVAL_2069;
  assign _EVAL_2024 = ~_EVAL_2389;
  assign _EVAL_2349 = 2'h3 == _EVAL_1541 ? _EVAL_767 : _EVAL_934;
  assign _EVAL_1580 = _EVAL_1065 ? _EVAL_1777 : {{2'd0}, _EVAL_540};
  assign _EVAL_96 = _EVAL_426 | _EVAL_288;
  assign _EVAL_1319 = _EVAL_151[7];
  assign _EVAL_1824 = _EVAL_1551[1];
  assign _EVAL_1563 = {{5'd0}, _EVAL_86};
  assign _EVAL_1643 = _EVAL_493 | _EVAL_2479;
  assign _EVAL_1609 = _EVAL_353 ? 5'hb : _EVAL_602;
  assign _EVAL_363 = ~_EVAL_2329;
  assign _EVAL_635 = _EVAL_700 ? 4'h3 : _EVAL_780;
  assign _EVAL_1440 = _EVAL_113 == 12'hb82;
  assign _EVAL_68 = _EVAL_834;
  assign _EVAL_99 = _EVAL_668;
  assign _EVAL_658 = _EVAL_113 == 12'hc9a;
  assign _EVAL_1682 = _EVAL_113 == 12'hb1a;
  assign _EVAL_2130 = _EVAL_1457 & _EVAL_2053;
  assign _EVAL_470 = _EVAL_151 == 12'hc80;
  assign _EVAL_876 = _EVAL_2199 | _EVAL_2517;
  assign _EVAL_291 = _EVAL_874 | _EVAL_2272;
  assign _EVAL_831 = _EVAL_2182 < 2'h1;
  assign _EVAL_180 = _EVAL_1065 & _EVAL_1147;
  assign _EVAL_31 = _EVAL_365;
  assign _EVAL_2225 = _EVAL_932 | _EVAL_1820;
  assign _EVAL_2052 = _EVAL_1385 | _EVAL_843;
  assign _EVAL_1290 = _EVAL_113 == 12'hc0f;
  assign _EVAL_2500 = ~_EVAL_985;
  assign _EVAL_55 = _EVAL_1280;
  assign _EVAL_1261 = _EVAL_2320 ? _EVAL_27 : _EVAL_133;
  assign _EVAL_1301 = _EVAL_360 | _EVAL_2047;
  assign _EVAL_1524 = _EVAL_888 ? 5'h17 : _EVAL_469;
  assign _EVAL_1586 = _EVAL_151 == 12'hf14;
  assign _EVAL_1964 = ~_EVAL_1017;
  assign _EVAL_533 = _EVAL_1702 ? _EVAL_1360 : _EVAL_760;
  assign _EVAL_25 = _EVAL_1595;
  assign _EVAL_943 = {{27'd0}, _EVAL_1264};
  assign _EVAL_754 = ~_EVAL_2160;
  assign _EVAL_2445 = _EVAL_2398 ? _EVAL_1124 : 64'h0;
  assign _EVAL_103 = _EVAL_1244[31:0];
  assign _EVAL_2437 = _EVAL_1456 | _EVAL_377;
  assign _EVAL_1151 = _EVAL_130[1];
  assign _EVAL_410 = _EVAL_863 | _EVAL_1203;
  assign _EVAL_2529 = _EVAL_1964 | _EVAL_2272;
  assign _EVAL_2212 = _EVAL_1005 & _EVAL_620;
  assign _EVAL_2211 = _EVAL_1525[1];
  assign _EVAL_1909 = 32'h80000000 + _EVAL_1181;
  assign _EVAL_1186 = _EVAL_1689 ? _EVAL_2486 : 32'h0;
  assign _EVAL_2326 = _EVAL_1551[21];
  assign _EVAL_2086 = _EVAL_314 | _EVAL_512;
  assign _EVAL_1648 = {{73'd0}, _EVAL_860};
  assign _EVAL_1988 = _EVAL_2066 | _EVAL_1758;
  assign _EVAL_862 = _EVAL_432 | _EVAL_2316;
  assign _EVAL_444 = _EVAL_1551[26];
  assign _EVAL_1795 = ~_EVAL_1287;
  assign _EVAL_295 = _EVAL_1953 | _EVAL_1430;
  assign _EVAL_1647 = _EVAL_151 == 12'h7b2;
  assign _EVAL_1660 = _EVAL_1015[30:0];
  assign _EVAL_2456 = _EVAL_1551[7];
  assign _EVAL_2030 = _EVAL_627 | _EVAL_1125;
  assign _EVAL_1495 = _EVAL_1212[1];
  assign _EVAL_2057 = _EVAL_2462 | _EVAL_1948;
  assign _EVAL_714 = _EVAL_2520 | _EVAL_2103;
  assign _EVAL_4 = _EVAL_2245;
  assign _EVAL_1739 = _EVAL_717 | _EVAL_503;
  assign _EVAL_2000 = _EVAL_113 == 12'h33b;
  assign _EVAL_1810 = _EVAL_528[39:32];
  assign _EVAL_1336 = _EVAL_113 == 12'hc0d;
  assign _EVAL_390 = _EVAL_1775 & _EVAL_2185;
  assign _EVAL_598 = _EVAL_1032 & _EVAL_382;
  assign _EVAL_1760 = _EVAL_445 | _EVAL_851;
  assign _EVAL_929 = _EVAL_387 & _EVAL_964;
  assign _EVAL_368 = _EVAL_113 == 12'h352;
  assign _EVAL_1832 = _EVAL_217 | _EVAL_210;
  assign _EVAL_171 = _EVAL_1696;
  assign _EVAL_723 = _EVAL_113 == 12'hf12;
  assign _EVAL_899 = _EVAL_113 == 12'hc00;
  assign _EVAL_1823 = _EVAL_363 | _EVAL_2058;
  assign _EVAL_1803 = _EVAL_1730 == 3'h0;
  assign _EVAL_666 = _EVAL_1363 | _EVAL_208;
  assign _EVAL_265 = _EVAL_910 | _EVAL_552;
  assign _EVAL_558 = ~_EVAL_2366;
  assign _EVAL_1946 = _EVAL_291 ? _EVAL_965 : _EVAL_1835;
  assign _EVAL_354 = _EVAL_477 | _EVAL_221;
  assign _EVAL_2421 = _EVAL_571 | _EVAL_2528;
  assign _EVAL_307 = _EVAL_1039 ? _EVAL_1733 : 5'h0;
  assign _EVAL_1532 = _EVAL_1535 | _EVAL_349;
  assign _EVAL_797 = {{71'd0}, _EVAL_599};
  assign _EVAL_847 = _EVAL_1793 | _EVAL_2456;
  assign _EVAL_818 = _EVAL_1407 | _EVAL_73;
  assign _EVAL_699 = _EVAL_679[1];
  assign _EVAL_1692 = _EVAL_2028[63:6];
  assign _EVAL_2140 = _EVAL_113 == 12'hc83;
  assign _EVAL_1730 = _EVAL_1484[7:5];
  assign _EVAL_1885 = _EVAL_113 == 12'hb80;
  assign _EVAL_1099 = _EVAL_113 == 12'hb9b;
  assign _EVAL_1612 = _EVAL_1698 ? _EVAL_1565 : _EVAL_1978;
  assign _EVAL_2361 = _EVAL_618[27];
  assign _EVAL_2209 = {_EVAL_113, 20'h0};
  assign _EVAL_1527 = _EVAL_113 == 12'hb12;
  assign _EVAL_1273 = _EVAL_517 ? 5'h7 : _EVAL_1030;
  assign _EVAL_196 = _EVAL_176 == 2'h0;
  assign _EVAL_1987 = _EVAL_1058 | _EVAL_2278;
  assign _EVAL_1050 = _EVAL_861 & _EVAL_1028;
  assign _EVAL_1218 = _EVAL_980 | _EVAL_2079;
  assign _EVAL_1634 = _EVAL_1678 | _EVAL_1963;
  assign _EVAL_637 = _EVAL_113 == 12'h32f;
  assign _EVAL_480 = _EVAL_1233 | _EVAL_2154;
  assign _EVAL_2409 = ~_EVAL_962;
  assign _EVAL_43 = _EVAL_2481;
  assign _EVAL_1208 = _EVAL_995 | _EVAL_952;
  assign _EVAL_1007 = _EVAL_2320 ? _EVAL_659 : 2'h3;
  assign _EVAL_38 = _EVAL_1557;
  assign _EVAL_100 = _EVAL_2182;
  assign _EVAL_188 = _EVAL_1111 | _EVAL_1901;
  assign _EVAL_807 = _EVAL_2249 | _EVAL_200;
  assign _EVAL_835 = _EVAL_2481[0];
  assign _EVAL_2142 = _EVAL_1562[13];
  assign _EVAL_1200 = _EVAL_2344 ? 5'h12 : _EVAL_2045;
  assign _EVAL_1398 = _EVAL_188 | _EVAL_2295;
  assign _EVAL_1222 = _EVAL_2304 == 32'h20000000;
  assign _EVAL_1971 = _EVAL_1723 | _EVAL_1854;
  assign _EVAL_2031 = _EVAL_1604 ? 4'h5 : _EVAL_1684;
  assign _EVAL_372 = _EVAL_2280[1];
  assign _EVAL_1976 = _EVAL_291 ? _EVAL_1989 : _EVAL_237;
  assign _EVAL_1863 = {{95'd0}, _EVAL_308};
  assign _EVAL_1203 = _EVAL_402[13];
  assign _EVAL_1683 = _EVAL_113 == 12'h336;
  assign _EVAL_704 = _EVAL_1551[12];
  assign _EVAL_2226 = _EVAL_113 == 12'hb96;
  assign _EVAL_2173 = {_EVAL_1707,2'h3};
  assign _EVAL_1255 = _EVAL_907 | _EVAL_1560;
  assign _EVAL_1806 = _EVAL_113 == 12'h342;
  assign _EVAL_2127 = ~_EVAL_2503;
  assign _EVAL_319 = _EVAL_1014 | _EVAL_1471;
  assign _EVAL_659 = _EVAL_1306 ? 2'h3 : _EVAL_2182;
  assign _EVAL_2476 = {84'h0,6'h0,_EVAL_965,2'h0,2'h0,2'h0,1'h0,_EVAL_1306,3'h0};
  assign _EVAL_2214 = _EVAL_585 | _EVAL_1016;
  assign _EVAL_655 = _EVAL_2338 ? _EVAL_359 : 30'h0;
  assign _EVAL_696 = _EVAL_1147 ? _EVAL_1959 : 32'h0;
  assign _EVAL_1686 = 2'h3 == _EVAL_1541 ? _EVAL_282 : _EVAL_1431;
  assign _EVAL_1852 = _EVAL_831 | _EVAL_390;
  assign _EVAL_2316 = _EVAL_113 == 12'hb1b;
  assign _EVAL_939 = _EVAL_1068[33:0];
  assign _EVAL_1779 = _EVAL_1080 & _EVAL_1421;
  assign _EVAL_2313 = {{98'd0}, _EVAL_307};
  assign _EVAL_297 = _EVAL_2057 | _EVAL_2309;
  assign _EVAL_1330 = _EVAL_2490[3];
  assign _EVAL_787 = _EVAL_113 < 12'hca0;
  assign _EVAL_2398 = _EVAL_151 == 12'hc00;
  assign _EVAL_2234 = _EVAL_2490 & 32'h7ff03;
  assign _EVAL_19 = _EVAL_531[31];
  assign _EVAL_1631 = _EVAL_113 == 12'hc17;
  assign _EVAL_638 = _EVAL_2490[6];
  assign _EVAL_142 = _EVAL_1620;
  assign _EVAL_757 = _EVAL_2535[1];
  assign _EVAL_2491 = _EVAL_2279 ? _EVAL_634 : _EVAL_2401;
  assign _EVAL_567 = _EVAL_2371 ? _EVAL_1946 : _EVAL_965;
  assign _EVAL_448 = _EVAL_113 == 12'hc0e;
  assign _EVAL_1472 = _EVAL_113 == 12'h7c0;
  assign _EVAL_629 = {4'h2,_EVAL_1017,14'h400,_EVAL_820,_EVAL_985,2'h0,_EVAL_2163,_EVAL_1874};
  assign _EVAL_1616 = _EVAL_1416[63:32];
  assign _EVAL_1826 = _EVAL_770 | _EVAL_1340;
  assign _EVAL_155 = _EVAL_2371;
  assign _EVAL_2077 = _EVAL_1404 ? 4'hc : _EVAL_2105;
  assign _EVAL_954 = _EVAL_151 == 12'h340;
  assign _EVAL_1684 = _EVAL_190 ? 4'h8 : {{1'd0}, _EVAL_379};
  assign _EVAL_2285 = _EVAL_429[30:0];
  assign _EVAL_2340 = _EVAL_1787[4:3];
  assign _EVAL_1388 = _EVAL_1710 & _EVAL_436;
  assign _EVAL_1422 = _EVAL_248 | _EVAL_1342;
  assign _EVAL_162 = _EVAL_2163;
  assign _EVAL_1861 = _EVAL_541 | _EVAL_1470;
  assign _EVAL_337 = _EVAL_1636 == 32'h20000000;
  assign _EVAL_138 = _EVAL_1478;
  assign _EVAL_759 = _EVAL_858 | _EVAL_388;
  assign _EVAL_2279 = _EVAL_2210 & _EVAL_386;
  assign _EVAL_1856 = _EVAL_1398 | _EVAL_2357;
  assign _EVAL_1220 = _EVAL_2026 & _EVAL_2500;
  assign _EVAL_1789 = _EVAL_402[29];
  assign _EVAL_1416 = {_EVAL_1062,_EVAL_2342};
  assign _EVAL_497 = _EVAL_2169 | _EVAL_2420;
  assign _EVAL_1264 = _EVAL_2108 ? 5'he : _EVAL_1436;
  assign _EVAL_1005 = _EVAL_2417 & _EVAL_1568;
  assign _EVAL_299 = _EVAL_1019 & _EVAL_782;
  assign _EVAL_33 = _EVAL_1618;
  assign _EVAL_379 = _EVAL_512 ? 3'h0 : 3'h4;
  assign _EVAL_2016 = _EVAL_802 ? _EVAL_1260 : 32'h0;
  assign _EVAL_1706 = {{31'd0}, _EVAL_1517};
  assign _EVAL_1431 = 2'h2 == _EVAL_1541 ? _EVAL_2366 : _EVAL_2036;
  assign _EVAL_1709 = ~_EVAL_1947;
  assign _EVAL_2374 = 32'h0;
  assign _EVAL_509 = _EVAL_2371 ? _EVAL_1313 : {{1'd0}, _EVAL_1280};
  assign _EVAL_195 = _EVAL_1350 ? _EVAL_939 : _EVAL_1817;
  assign _EVAL_2074 = _EVAL_1057 | _EVAL_2165;
  assign _EVAL_144 = _EVAL_540;
  assign _EVAL_14 = _EVAL_1113;
  assign _EVAL_1983 = _EVAL_823 & _EVAL_1319;
  assign _EVAL_79 = _EVAL_1955;
  assign _EVAL_2449 = {{73'd0}, _EVAL_401};
  assign _EVAL_1886 = _EVAL_2538 | _EVAL_1829;
  assign _EVAL_0 = _EVAL_395;
  assign _EVAL_2484 = _EVAL_113 == 12'hc1a;
  assign _EVAL_1598 = _EVAL_1921 | _EVAL_281;
  assign _EVAL = _EVAL_1532 | _EVAL_542;
  assign _EVAL_1995 = _EVAL_1981 | _EVAL_1735;
  assign _EVAL_661 = _EVAL_2488 ? 5'h11 : _EVAL_889;
  assign _EVAL_694 = _EVAL_1643 | _EVAL_1291;
  assign _EVAL_1056 = ~_EVAL_878;
  assign _EVAL_2037 = ~_EVAL_1151;
  assign _EVAL_94 = _EVAL_1998[31:0];
  assign _EVAL_1866 = _EVAL_1424 | _EVAL_779;
  assign _EVAL_1748 = {{71'd0}, _EVAL_870};
  assign _EVAL_1873 = _EVAL_113 == 12'h3a3;
  assign _EVAL_373 = ~_EVAL_1319;
  assign _EVAL_2510 = _EVAL_2550 + 58'h1;
  assign _EVAL_1181 = {{1'd0}, _EVAL_739};
  assign _EVAL_2477 = _EVAL_1023 ? 5'hd : _EVAL_2170;
  assign _EVAL_1594 = _EVAL_291 ? {{20'd0}, _EVAL_2011} : _EVAL_1293;
  assign _EVAL_1669 = {{71'd0}, _EVAL_1629};
  assign _EVAL_499 = _EVAL_113 == 12'hb0a;
  assign _EVAL_2166 = _EVAL_1487 ? _EVAL_685 : 32'h0;
  assign _EVAL_30 = _EVAL_2159;
  assign _EVAL_773 = _EVAL_113[10];
  assign _EVAL_212 = _EVAL_1212[0];
  assign _EVAL_1262 = _EVAL_1753 | _EVAL_535;
  assign _EVAL_1275 = _EVAL_1957 | _EVAL_1699;
  assign _EVAL_1219 = _EVAL_2200 ? _EVAL_2490 : {{2'd0}, _EVAL_1910};
  assign _EVAL_936 = ~_EVAL_1796;
  assign _EVAL_2410 = _EVAL_113 == 12'h32b;
  assign _EVAL_1928 = ~_EVAL_2391;
  assign _EVAL_91 = _EVAL_2331;
  assign _EVAL_1355 = _EVAL_291 ? _EVAL_1070 : _EVAL_1999;
  assign _EVAL_2148 = _EVAL_1065 ? _EVAL_1455 : {{2'd0}, _EVAL_1813};
  assign _EVAL_2396 = _EVAL_113 == 12'hb84;
  assign _EVAL_234 = _EVAL_2248 + _EVAL_488;
  assign _EVAL_1845 = _EVAL_580 & _EVAL_2516;
  assign _EVAL_549 = _EVAL_1327[7];
  assign _EVAL_1436 = _EVAL_817 ? 5'hd : _EVAL_2412;
  assign _EVAL_1677 = _EVAL_222 + 31'h1;
  assign _EVAL_8 = _EVAL_454;
  assign _EVAL_2026 = _EVAL_1890[11];
  assign _EVAL_2269 = _EVAL_1318 & _EVAL_1931;
  assign _EVAL_316 = _EVAL_319 | _EVAL_1550;
  assign _EVAL_735 = _EVAL_2328[39:32];
  assign _EVAL_607 = _EVAL_528[31:0];
  assign _EVAL_217 = _EVAL_1160 | _EVAL_2223;
  assign _EVAL_388 = _EVAL_113 == 12'hc08;
  assign _EVAL_595 = _EVAL_973 & _EVAL_357;
  assign _EVAL_688 = _EVAL_2069 | _EVAL_1050;
  assign _EVAL_1427 = _EVAL_476 | _EVAL_628;
  assign _EVAL_1773 = {_EVAL_2,_EVAL_164,_EVAL_68,_EVAL_56,_EVAL_24,_EVAL_100,_EVAL_96,_EVAL_122,_EVAL_2379,_EVAL_966};
  assign _EVAL_1285 = _EVAL_1767 | _EVAL_2142;
  assign _EVAL_1891 = _EVAL_1085 == 12'h410;
  assign _EVAL_1744 = _EVAL_1065 ? _EVAL_1219 : {{2'd0}, _EVAL_1910};
  assign _EVAL_1038 = _EVAL_2342 + _EVAL_1137;
  assign _EVAL_58 = _EVAL_1796;
  assign _EVAL_775 = _EVAL_504[0];
  assign _EVAL_318 = _EVAL_1183 | _EVAL_2413;
  assign _EVAL_1565 = ~_EVAL_1991;
  assign _EVAL_123 = _EVAL_1212;
  assign _EVAL_2146 = _EVAL_2250 | _EVAL_2369;
  assign _EVAL_2196 = _EVAL_2535[12];
  assign _EVAL_1266 = ~_EVAL_450;
  assign _EVAL_616 = {{71'd0}, _EVAL_1661};
  assign _EVAL_554 = _EVAL_1019 & _EVAL_1928;
  assign _EVAL_2365 = _EVAL_113 == 12'h7a2;
  assign _EVAL_1812 = _EVAL_1172 ? _EVAL_521 : 8'h0;
  assign _EVAL_1358 = _EVAL_113 == 12'hb14;
  assign _EVAL_2399 = _EVAL_973 ? _EVAL_592 : 32'h0;
  assign _EVAL_1019 = _EVAL_151 == 12'h3a0;
  assign _EVAL_2172 = _EVAL_2042 & 32'hfffffff0;
  assign _EVAL_539 = _EVAL_113 == 12'hb1c;
  assign _EVAL_632 = _EVAL_2421 | _EVAL_1631;
  assign _EVAL_118 = _EVAL_1217;
  assign _EVAL_892 = _EVAL_1753 ? _EVAL_192 : 1'h1;
  assign _EVAL_1141 = _EVAL_1442 & _EVAL_2188;
  assign _EVAL_2048 = _EVAL_222 & _EVAL_1857;
  assign _EVAL_2432 = _EVAL_113 == 12'h3b5;
  assign _EVAL_836 = _EVAL_1019 & _EVAL_563;
  assign _EVAL_350 = _EVAL_1551[9];
  assign _EVAL_2323 = _EVAL_564[0];
  assign _EVAL_1695 = _EVAL_2182 <= 2'h1;
  assign _EVAL_720 = _EVAL_1039 ? _EVAL_2025 : {{27'd0}, _EVAL_1733};
  assign _EVAL_565 = _EVAL_113 == 12'hb0b;
  assign _EVAL_1406 = _EVAL_1562[12];
  assign _EVAL_357 = ~_EVAL_454;
  assign _EVAL_1762 = _EVAL_1647 ? _EVAL_1159 : 32'h0;
  assign _EVAL_548 = _EVAL_2427[27];
  assign _EVAL_1172 = _EVAL_151 == 12'hc84;
  assign _EVAL_1345 = _EVAL_1161 & _EVAL_573;
  assign _EVAL_1936 = _EVAL_1886 | _EVAL_1358;
  assign _EVAL_182 = _EVAL_630;
  assign _EVAL_2066 = _EVAL_1182 | _EVAL_1898;
  assign _EVAL_1537 = _EVAL_1733[3];
  assign _EVAL_139 = _EVAL_461;
  assign _EVAL_2282 = ~_EVAL_1533;
  assign _EVAL_2119 = _EVAL_2296 & _EVAL_861;
  assign _EVAL_1233 = _EVAL_1826 | _EVAL_2255;
  assign _EVAL_535 = _EVAL_2371 ? _EVAL_1164 : _EVAL_1306;
  assign _EVAL_143 = 2'h1;
  assign _EVAL_2271 = _EVAL_2535[8];
  assign _EVAL_2247 = _EVAL_1038[6];
  assign _EVAL_2495 = _EVAL_402[27];
  assign _EVAL_1688 = _EVAL_1479 | _EVAL_1942;
  assign _EVAL_1323 = _EVAL_151 == 12'h352;
  assign _EVAL_882 = _EVAL_151 == 12'hb03;
  assign _EVAL_2367 = _EVAL_1065 ? _EVAL_732 : {{2'd0}, _EVAL_359};
  assign _EVAL_178 = _EVAL_985;
  assign _EVAL_921 = _EVAL_2104 | _EVAL_2034;
  assign _EVAL_2021 = _EVAL_1082 | _EVAL_1665;
  assign _EVAL_1911 = _EVAL_1554[12];
  assign _EVAL_832 = _EVAL_1689 ? _EVAL_1190 : 32'h0;
  assign _EVAL_1396 = _EVAL_281 ? 5'h9 : _EVAL_968;
  assign _EVAL_209 = _EVAL_2505 & _EVAL_1663;
  assign _EVAL_579 = _EVAL_1558[0];
  assign _EVAL_1919 = _EVAL_937 & _EVAL_1698;
  assign _EVAL_580 = _EVAL_2427[11];
  assign _EVAL_2333 = _EVAL_1445 + 31'h1;
  assign _EVAL_2535 = {_EVAL_20, 14'h0};
  assign _EVAL_1270 = _EVAL_1484 == 8'hd;
  assign _EVAL_2007 = _EVAL_113 == 12'hc19;
  assign _EVAL_1735 = _EVAL_113 == 12'hc87;
  assign _EVAL_1438 = _EVAL_819[7];
  assign _EVAL_2277 = _EVAL_2247 & _EVAL_1736;
  assign _EVAL_701 = _EVAL_151 == 12'hb04;
  assign _EVAL_1097 = _EVAL_1710 | _EVAL_558;
  assign _EVAL_1214 = _EVAL_1418 | _EVAL_1789;
  assign _EVAL_2547 = _EVAL_2489 | _EVAL_1374;
  assign _EVAL_833 = _EVAL_2153 | _EVAL_1745;
  assign _EVAL_2255 = {{95'd0}, _EVAL_1812};
  assign _EVAL_1487 = _EVAL_151 == 12'h344;
  assign _EVAL_1221 = {_EVAL_804,_EVAL_245,_EVAL_1761,_EVAL_2426};
  assign _EVAL_173 = _EVAL_1227;
  assign _EVAL_2304 = _EVAL_2209 & 32'h20400000;
  assign _EVAL_1168 = _EVAL_441 & 32'h20100000;
  assign _EVAL_1312 = _EVAL_260 | _EVAL_734;
  assign _EVAL_2467 = _EVAL_2518 | _EVAL_2504;
  assign _EVAL_2043 = _EVAL_506 ? 5'h16 : _EVAL_1512;
  assign _EVAL_194 = _EVAL_2490[1];
  assign _EVAL_515 = _EVAL_1327[3];
  assign _EVAL_2088 = ~_EVAL_417;
  assign _EVAL_391 = _EVAL_1327[12:11];
  assign _EVAL_879 = _EVAL_2442 & _EVAL_1950;
  assign _EVAL_128 = _EVAL_2425;
  assign _EVAL_747 = _EVAL_684 | _EVAL_191;
  assign _EVAL_505 = _EVAL_1779 ? _EVAL_2490 : {{2'd0}, _EVAL_1155};
  assign _EVAL_906 = _EVAL_564[2];
  assign _EVAL_358 = _EVAL_113 == 12'h324;
  assign _EVAL_404 = _EVAL_819[2];
  assign _EVAL_1304 = _EVAL_2447 ? _EVAL_2124 : _EVAL_1083;
  assign _EVAL_2400 = _EVAL_113 == 12'hc82;
  assign _EVAL_671 = 2'h3 == _EVAL_1541 ? 1'h0 : _EVAL_2536;
  assign _EVAL_683 = _EVAL_1289 | _EVAL_1476;
  assign _EVAL_572 = _EVAL_2510[57:0];
  assign _EVAL_1707 = _EVAL_1445 & _EVAL_1985;
  assign _EVAL_473 = {{95'd0}, _EVAL_1239};
  assign _EVAL_1502 = _EVAL_361 | _EVAL_2060;
  assign _EVAL_222 = {_EVAL_227,_EVAL_1395};
  assign _EVAL_1723 = _EVAL_2014 | _EVAL_2544;
  assign _EVAL_283 = _EVAL_1415 ? 5'h17 : _EVAL_2043;
  assign _EVAL_844 = _EVAL_113 == 12'hf13;
  assign _EVAL_1621 = _EVAL_2306 ? _EVAL_855 : 32'h0;
  assign _EVAL_119 = _EVAL_1849;
  assign _EVAL_413 = _EVAL_881 ? 32'h489 : 32'h0;
  assign _EVAL_1922 = _EVAL_1756 + 31'h1;
  assign _EVAL_2498 = _EVAL_1983 ? _EVAL_849 : _EVAL_1651;
  assign _EVAL_1031 = _EVAL_151 == 12'h306;
  assign _EVAL_1322 = _EVAL_2182[0];
  assign _EVAL_481 = _EVAL_1551[15];
  assign _EVAL_1131 = _EVAL_1755[6];
  assign _EVAL_2206 = _EVAL_2221 | _EVAL_1493;
  assign _EVAL_2537 = _EVAL_1306 & _EVAL_1852;
  assign _EVAL_1708 = _EVAL_2501 | _EVAL_1939;
  assign _EVAL_74 = _EVAL_2465;
  assign _EVAL_2486 = {4'h2,_EVAL_962,14'h400,_EVAL_1344,_EVAL_1796,2'h0,_EVAL_1113,_EVAL_1725};
  assign _EVAL_2246 = _EVAL_151 == 12'h7a1;
  assign _EVAL_302 = _EVAL_1065 ? _EVAL_1304 : {{57'd0}, _EVAL_1968};
  assign _EVAL_564 = _EVAL_2490[31:24];
  assign _EVAL_910 = _EVAL_2471 | _EVAL_797;
  assign _EVAL_715 = _EVAL_1102 | _EVAL_1721;
  assign _EVAL_2150 = _EVAL_2527 ? 5'hb : _EVAL_1933;
  assign _EVAL_336 = _EVAL_1789 ? 5'h1d : _EVAL_1770;
  assign _EVAL_1654 = _EVAL_402[25];
  assign _EVAL_218 = _EVAL_1220 & _EVAL_1637;
  assign _EVAL_972 = _EVAL_1987 | _EVAL_1391;
  assign _EVAL_2283 = _EVAL_239 | _EVAL_710;
  assign _EVAL_1329 = _EVAL_446 | _EVAL_704;
  assign _EVAL_1289 = _EVAL_2551 | _EVAL_1472;
  assign _EVAL_334 = _EVAL_113 == 12'hc9f;
  assign _EVAL_2098 = _EVAL_1551[5];
  assign _EVAL_753 = _EVAL_2366 | _EVAL_2088;
  assign _EVAL_1012 = _EVAL_665 & _EVAL_1401;
  assign _EVAL_2502 = _EVAL_2377 ? 4'he : _EVAL_2144;
  assign _EVAL_1923 = _EVAL_1551[25];
  assign _EVAL_239 = _EVAL_345 | _EVAL_2151;
  assign _EVAL_1424 = _EVAL_784 | _EVAL_2092;
  assign _EVAL_2117 = _EVAL_1323 ? _EVAL_1070 : 32'h0;
  assign _EVAL_2427 = _EVAL_818 & _EVAL_490;
  assign _EVAL_727 = 2'h3 == _EVAL_1541 ? _EVAL_1696 : _EVAL_1451;
  assign _EVAL_657 = _EVAL_275 | _EVAL_1099;
  assign _EVAL_436 = _EVAL_2427[12];
  assign _EVAL_1036 = _EVAL_113 == 12'h3ba;
  assign _EVAL_532 = {{39'd0}, _EVAL_2175};
  assign _EVAL_707 = _EVAL_113 == 12'h350;
  assign _EVAL_1006 = _EVAL_472 | _EVAL_1941;
  assign _EVAL_2524 = 2'h1 == _EVAL_1541 ? _EVAL_1620 : _EVAL_1657;
  assign _EVAL_932 = _EVAL_316 | _EVAL_803;
  assign _EVAL_2072 = _EVAL_113 == 12'hc8a;
  assign _EVAL_2393 = _EVAL_151 == 12'h3b1;
  assign _EVAL_2268 = ~_EVAL_282;
  assign _EVAL_1898 = _EVAL_113 == 12'hc1f;
  always @(posedge _EVAL_85) begin
    _EVAL_227 <= _EVAL_254[29:0];
    if (_EVAL_83) begin
      _EVAL_237 <= 2'h3;
    end else if (_EVAL_1065) begin
      if (_EVAL_2192) begin
        if (_EVAL_983) begin
          _EVAL_237 <= 2'h3;
        end else begin
          _EVAL_237 <= 2'h0;
        end
      end else begin
        _EVAL_237 <= _EVAL_1498;
      end
    end else begin
      _EVAL_237 <= _EVAL_1498;
    end
    if (_EVAL_83) begin
      _EVAL_245 <= 1'h0;
    end
    if (_EVAL_83) begin
      _EVAL_280 <= 32'h40901105;
    end else if (_EVAL_1065) begin
      if (_EVAL_909) begin
        if (_EVAL_1724) begin
          _EVAL_280 <= _EVAL_919;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_282 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_1573) begin
        if (_EVAL_2246) begin
          _EVAL_282 <= _EVAL_1288;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_312 <= 2'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_554) begin
        _EVAL_312 <= _EVAL_1047;
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_836) begin
        _EVAL_313 <= _EVAL_1410;
      end
    end
    _EVAL_359 <= _EVAL_2367[29:0];
    if (_EVAL_83) begin
      _EVAL_365 <= 2'h3;
    end else if (_EVAL_1065) begin
      if (_EVAL_802) begin
        if (_EVAL_590) begin
          _EVAL_365 <= 2'h3;
        end else begin
          _EVAL_365 <= 2'h0;
        end
      end else begin
        _EVAL_365 <= _EVAL_873;
      end
    end else begin
      _EVAL_365 <= _EVAL_873;
    end
    if (_EVAL_83) begin
      _EVAL_366 <= 1'h0;
    end
    if (_EVAL_1065) begin
      if (_EVAL_595) begin
        _EVAL_370 <= _EVAL_1926;
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_2284) begin
        if (_EVAL_2343) begin
          _EVAL_385 <= _EVAL_2490;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_387 <= 32'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_1084) begin
        _EVAL_387 <= _EVAL_2490;
      end
    end
    if (_EVAL_83) begin
      _EVAL_395 <= 2'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_836) begin
        _EVAL_395 <= _EVAL_856;
      end
    end
    if (_EVAL_83) begin
      _EVAL_417 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_2284) begin
        if (_EVAL_2246) begin
          _EVAL_417 <= _EVAL_218;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_454 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_595) begin
        _EVAL_454 <= _EVAL_912;
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_1573) begin
        if (_EVAL_2246) begin
          _EVAL_460 <= _EVAL_1330;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_461 <= 2'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_1715) begin
        _EVAL_461 <= _EVAL_1807;
      end
    end
    _EVAL_498 <= _EVAL_256[5:0];
    if (_EVAL_83) begin
      _EVAL_500 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_2284) begin
        if (_EVAL_2246) begin
          _EVAL_500 <= _EVAL_672;
        end
      end
    end
    _EVAL_540 <= _EVAL_1580[29:0];
    if (_EVAL_83) begin
      _EVAL_611 <= 1'h0;
    end
    if (_EVAL_83) begin
      _EVAL_617 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_2284) begin
        if (_EVAL_2246) begin
          _EVAL_617 <= _EVAL_1819;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_630 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_1573) begin
        if (_EVAL_2246) begin
          _EVAL_630 <= _EVAL_672;
        end
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_1573) begin
        if (_EVAL_2343) begin
          _EVAL_647 <= _EVAL_2490;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_665 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_612) begin
        _EVAL_665 <= _EVAL_768;
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_612) begin
        _EVAL_668 <= _EVAL_1907;
      end
    end
    if (_EVAL_83) begin
      _EVAL_679 <= 2'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_1897) begin
        _EVAL_679 <= _EVAL_1807;
      end
    end
    if (_EVAL_83) begin
      _EVAL_689 <= 12'h0;
    end
    if (_EVAL_83) begin
      _EVAL_722 <= 8'h0;
    end
    if (_EVAL_83) begin
      _EVAL_740 <= 3'h0;
    end else if (_EVAL_2371) begin
      if (_EVAL_291) begin
        if (_EVAL_1698) begin
          _EVAL_740 <= _EVAL_2385;
        end
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_885) begin
        _EVAL_741 <= _EVAL_404;
      end
    end
    if (_EVAL_83) begin
      _EVAL_743 <= 1'h0;
    end
    if (_EVAL_1065) begin
      if (_EVAL_1573) begin
        if (_EVAL_2246) begin
          _EVAL_767 <= _EVAL_638;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_793 <= 1'h0;
    end
    if (_EVAL_1065) begin
      if (_EVAL_554) begin
        _EVAL_795 <= _EVAL_228;
      end
    end
    if (_EVAL_83) begin
      _EVAL_799 <= 1'h0;
    end
    if (_EVAL_83) begin
      _EVAL_804 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_2192) begin
        _EVAL_804 <= _EVAL_501;
      end
    end
    if (_EVAL_83) begin
      _EVAL_820 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_1588) begin
        if (_EVAL_2246) begin
          _EVAL_820 <= _EVAL_1388;
        end
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_2306) begin
        _EVAL_855 <= _EVAL_2490;
      end
    end
    if (_EVAL_83) begin
      _EVAL_872 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_1588) begin
        if (_EVAL_2246) begin
          _EVAL_872 <= _EVAL_1819;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_877 <= 2'h0;
    end
    if (_EVAL_83) begin
      _EVAL_890 <= 2'h0;
    end
    if (_EVAL_1065) begin
      if (_EVAL_299) begin
        _EVAL_891 <= _EVAL_2017;
      end
    end
    if (_EVAL_83) begin
      _EVAL_905 <= 1'h0;
    end
    if (_EVAL_83) begin
      _EVAL_937 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_802) begin
        _EVAL_937 <= _EVAL_1118;
      end else begin
        _EVAL_937 <= _EVAL_527;
      end
    end else begin
      _EVAL_937 <= _EVAL_527;
    end
    if (_EVAL_83) begin
      _EVAL_949 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_1588) begin
        if (_EVAL_2246) begin
          _EVAL_949 <= _EVAL_194;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_962 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_726) begin
        if (_EVAL_2246) begin
          _EVAL_962 <= _EVAL_332;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_965 <= 2'h3;
    end else if (_EVAL_1065) begin
      if (_EVAL_1702) begin
        if (_EVAL_590) begin
          _EVAL_965 <= 2'h3;
        end else begin
          _EVAL_965 <= 2'h0;
        end
      end else begin
        _EVAL_965 <= _EVAL_567;
      end
    end else begin
      _EVAL_965 <= _EVAL_567;
    end
    if (_EVAL_83) begin
      _EVAL_985 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_1588) begin
        if (_EVAL_2246) begin
          _EVAL_985 <= _EVAL_324;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_1001 <= 2'h1;
    end
    if (_EVAL_83) begin
      _EVAL_1017 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_1588) begin
        if (_EVAL_2246) begin
          _EVAL_1017 <= _EVAL_1710;
        end
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_612) begin
        _EVAL_1027 <= _EVAL_228;
      end
    end
    if (_EVAL_83) begin
      _EVAL_1032 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_1897) begin
        _EVAL_1032 <= _EVAL_1952;
      end
    end
    if (_EVAL_83) begin
      _EVAL_1059 <= 2'h0;
    end
    if (_EVAL_83) begin
      _EVAL_1062 <= 58'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_2447) begin
        _EVAL_1062 <= _EVAL_437;
      end else if (_EVAL_1567) begin
        _EVAL_1062 <= _EVAL_1833;
      end else begin
        _EVAL_1062 <= _EVAL_1798;
      end
    end else begin
      _EVAL_1062 <= _EVAL_1798;
    end
    if (_EVAL_83) begin
      _EVAL_1070 <= 32'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_1323) begin
        _EVAL_1070 <= _EVAL_640;
      end else begin
        _EVAL_1070 <= _EVAL_1297;
      end
    end else begin
      _EVAL_1070 <= _EVAL_1297;
    end
    if (_EVAL_83) begin
      _EVAL_1075 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_726) begin
        if (_EVAL_2246) begin
          _EVAL_1075 <= _EVAL_194;
        end
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_726) begin
        if (_EVAL_2246) begin
          _EVAL_1113 <= _EVAL_2003;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_1120 <= 1'h0;
    end
    _EVAL_1155 <= _EVAL_1389[29:0];
    if (_EVAL_1065) begin
      if (_EVAL_1647) begin
        _EVAL_1159 <= _EVAL_2490;
      end
    end
    if (_EVAL_83) begin
      _EVAL_1161 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_1715) begin
        _EVAL_1161 <= _EVAL_1952;
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_1526) begin
        _EVAL_1187 <= _EVAL_1492;
      end else begin
        _EVAL_1187 <= _EVAL_1116;
      end
    end else begin
      _EVAL_1187 <= _EVAL_1116;
    end
    if (_EVAL_83) begin
      _EVAL_1206 <= 1'h0;
    end
    if (_EVAL_83) begin
      _EVAL_1212 <= 2'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_885) begin
        _EVAL_1212 <= _EVAL_856;
      end
    end
    if (_EVAL_83) begin
      _EVAL_1213 <= 27'h0;
    end
    if (_EVAL_83) begin
      _EVAL_1217 <= 32'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_2041) begin
        _EVAL_1217 <= _EVAL_2234;
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_836) begin
        _EVAL_1227 <= _EVAL_1794;
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_1897) begin
        _EVAL_1229 <= _EVAL_906;
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_595) begin
        _EVAL_1231 <= _EVAL_2017;
      end
    end
    if (_EVAL_83) begin
      _EVAL_1280 <= 1'h0;
    end else begin
      _EVAL_1280 <= _EVAL_509[0];
    end
    if (_EVAL_1065) begin
      if (_EVAL_2284) begin
        if (_EVAL_2246) begin
          _EVAL_1300 <= _EVAL_1330;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_1302 <= 32'h0;
    end
    _EVAL_1306 <= _EVAL_83 | _EVAL_2018;
    if (_EVAL_1065) begin
      if (_EVAL_2284) begin
        if (_EVAL_2246) begin
          _EVAL_1326 <= _EVAL_638;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_1334 <= 32'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_2063) begin
        _EVAL_1334 <= _EVAL_2234;
      end
    end
    if (_EVAL_83) begin
      _EVAL_1344 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_726) begin
        if (_EVAL_2246) begin
          _EVAL_1344 <= _EVAL_1201;
        end
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_1588) begin
        if (_EVAL_2343) begin
          _EVAL_1357 <= _EVAL_2490;
        end
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_554) begin
        _EVAL_1383 <= _EVAL_1088;
      end
    end
    if (_EVAL_83) begin
      _EVAL_1399 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_802) begin
        _EVAL_1399 <= _EVAL_549;
      end else begin
        _EVAL_1399 <= _EVAL_351;
      end
    end else begin
      _EVAL_1399 <= _EVAL_351;
    end
    if (_EVAL_1065) begin
      if (_EVAL_1311) begin
        _EVAL_1439 <= _EVAL_2133;
      end else if (_EVAL_882) begin
        _EVAL_1439 <= _EVAL_1834;
      end else begin
        _EVAL_1439 <= _EVAL_1126;
      end
    end else begin
      _EVAL_1439 <= _EVAL_1126;
    end
    if (_EVAL_83) begin
      _EVAL_1463 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_726) begin
        if (_EVAL_2246) begin
          _EVAL_1463 <= _EVAL_1819;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_1478 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_1573) begin
        if (_EVAL_2246) begin
          _EVAL_1478 <= _EVAL_1204;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_1496 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_2192) begin
        _EVAL_1496 <= _EVAL_672;
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_1715) begin
        _EVAL_1504 <= _EVAL_2323;
      end
    end
    _EVAL_1505 <= _EVAL_2345[5:0];
    if (_EVAL_83) begin
      _EVAL_1511 <= 2'h0;
    end
    if (_EVAL_83) begin
      _EVAL_1525 <= 2'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_612) begin
        _EVAL_1525 <= _EVAL_1047;
      end
    end
    if (_EVAL_83) begin
      _EVAL_1534 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_802) begin
        _EVAL_1534 <= _EVAL_515;
      end else begin
        _EVAL_1534 <= _EVAL_2491;
      end
    end else begin
      _EVAL_1534 <= _EVAL_2491;
    end
    _EVAL_1541 <= _EVAL_2446[1:0];
    if (_EVAL_83) begin
      _EVAL_1545 <= 1'h0;
    end
    if (_EVAL_1065) begin
      if (_EVAL_836) begin
        _EVAL_1557 <= _EVAL_404;
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_885) begin
        _EVAL_1595 <= _EVAL_1410;
      end
    end
    if (_EVAL_83) begin
      _EVAL_1618 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_1588) begin
        if (_EVAL_2246) begin
          _EVAL_1618 <= _EVAL_672;
        end
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_1588) begin
        if (_EVAL_2246) begin
          _EVAL_1620 <= _EVAL_1330;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_1633 <= 2'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_802) begin
        _EVAL_1633 <= 2'h0;
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_726) begin
        if (_EVAL_2246) begin
          _EVAL_1657 <= _EVAL_1330;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_1672 <= 1'h0;
    end
    if (_EVAL_1065) begin
      if (_EVAL_1897) begin
        _EVAL_1694 <= _EVAL_1869;
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_1573) begin
        if (_EVAL_2246) begin
          _EVAL_1696 <= _EVAL_2003;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_1733 <= 5'h0;
    end else begin
      _EVAL_1733 <= _EVAL_896[4:0];
    end
    if (_EVAL_83) begin
      _EVAL_1738 <= 2'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_299) begin
        _EVAL_1738 <= _EVAL_2340;
      end
    end
    if (_EVAL_83) begin
      _EVAL_1757 <= 1'h0;
    end
    if (_EVAL_83) begin
      _EVAL_1761 <= 1'h0;
    end
    if (_EVAL_1065) begin
      if (_EVAL_299) begin
        _EVAL_1788 <= _EVAL_1926;
      end
    end
    if (_EVAL_83) begin
      _EVAL_1796 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_726) begin
        if (_EVAL_2246) begin
          _EVAL_1796 <= _EVAL_2269;
        end
      end
    end
    _EVAL_1813 <= _EVAL_2148[29:0];
    if (_EVAL_1065) begin
      if (_EVAL_1912) begin
        _EVAL_1817 <= _EVAL_2334;
      end else if (_EVAL_701) begin
        _EVAL_1817 <= _EVAL_589;
      end else begin
        _EVAL_1817 <= _EVAL_195;
      end
    end else begin
      _EVAL_1817 <= _EVAL_195;
    end
    if (_EVAL_83) begin
      _EVAL_1828 <= 2'h0;
    end
    _EVAL_1847 <= _EVAL_1847;
    if (_EVAL_1065) begin
      if (_EVAL_299) begin
        _EVAL_1849 <= _EVAL_1468;
      end
    end
    if (_EVAL_83) begin
      _EVAL_1858 <= 2'h0;
    end
    if (_EVAL_1065) begin
      if (_EVAL_885) begin
        _EVAL_1867 <= _EVAL_1794;
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_954) begin
        _EVAL_1870 <= _EVAL_2490;
      end
    end
    if (_EVAL_83) begin
      _EVAL_1878 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_1573) begin
        if (_EVAL_2246) begin
          _EVAL_1878 <= _EVAL_1819;
        end
      end
    end
    _EVAL_1910 <= _EVAL_1744[29:0];
    if (_EVAL_83) begin
      _EVAL_1918 <= 1'h0;
    end
    if (_EVAL_1065) begin
      if (_EVAL_612) begin
        _EVAL_1920 <= _EVAL_1088;
      end
    end
    if (_EVAL_83) begin
      _EVAL_1935 <= 1'h0;
    end
    if (_EVAL_83) begin
      _EVAL_1947 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_885) begin
        _EVAL_1947 <= _EVAL_1438;
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_1715) begin
        _EVAL_1955 <= _EVAL_1869;
      end
    end
    if (_EVAL_83) begin
      _EVAL_1959 <= 32'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_1147) begin
        _EVAL_1959 <= _EVAL_2263;
      end
    end
    if (_EVAL_83) begin
      _EVAL_1967 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_1573) begin
        if (_EVAL_2246) begin
          _EVAL_1967 <= _EVAL_194;
        end
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_2530) begin
        _EVAL_1978 <= _EVAL_1492;
      end else begin
        _EVAL_1978 <= _EVAL_956;
      end
    end else begin
      _EVAL_1978 <= _EVAL_956;
    end
    if (_EVAL_83) begin
      _EVAL_2042 <= 32'hf;
    end else if (_EVAL_1065) begin
      if (_EVAL_2064) begin
        _EVAL_2042 <= _EVAL_1211;
      end
    end
    if (_EVAL_244) begin
      _EVAL_2069 <= 1'h0;
    end else begin
      _EVAL_2069 <= _EVAL_516;
    end
    if (_EVAL_83) begin
      _EVAL_2075 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_2284) begin
        if (_EVAL_2246) begin
          _EVAL_2075 <= _EVAL_2212;
        end
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_2284) begin
        if (_EVAL_2246) begin
          _EVAL_2082 <= _EVAL_2003;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_2099 <= 32'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_1839) begin
        _EVAL_2099 <= _EVAL_2487;
      end else begin
        _EVAL_2099 <= _EVAL_597;
      end
    end else begin
      _EVAL_2099 <= _EVAL_597;
    end
    if (_EVAL_1065) begin
      if (_EVAL_419) begin
        _EVAL_2128 <= _EVAL_705;
      end
    end
    if (_EVAL_83) begin
      _EVAL_2149 <= 1'h0;
    end
    if (_EVAL_1065) begin
      if (_EVAL_595) begin
        _EVAL_2159 <= _EVAL_1468;
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_1588) begin
        if (_EVAL_2246) begin
          _EVAL_2163 <= _EVAL_2003;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_2174 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_836) begin
        _EVAL_2174 <= _EVAL_1438;
      end
    end
    if (_EVAL_83) begin
      _EVAL_2182 <= 2'h3;
    end else if (_EVAL_579) begin
      _EVAL_2182 <= 2'h3;
    end else begin
      _EVAL_2182 <= 2'h0;
    end
    if (_EVAL_83) begin
      _EVAL_2185 <= 1'h0;
    end
    if (_EVAL_1065) begin
      if (_EVAL_726) begin
        if (_EVAL_2343) begin
          _EVAL_2245 <= _EVAL_2490;
        end
      end
    end
    _EVAL_2262 <= _EVAL_2441[29:0];
    if (_EVAL_83) begin
      _EVAL_2272 <= 1'h0;
    end else if (_EVAL_2279) begin
      if (_EVAL_1983) begin
        _EVAL_2272 <= 1'h0;
      end else begin
        _EVAL_2272 <= _EVAL_1425;
      end
    end else begin
      _EVAL_2272 <= _EVAL_1425;
    end
    if (_EVAL_1919) begin
      _EVAL_2297 <= _EVAL_365;
    end else begin
      _EVAL_2297 <= _EVAL_2182;
    end
    if (_EVAL_83) begin
      _EVAL_2301 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_2284) begin
        if (_EVAL_2246) begin
          _EVAL_2301 <= _EVAL_194;
        end
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_2359) begin
        _EVAL_2315 <= _EVAL_2490;
      end else begin
        _EVAL_2315 <= _EVAL_2392;
      end
    end else begin
      _EVAL_2315 <= _EVAL_2392;
    end
    if (_EVAL_1065) begin
      if (_EVAL_1136) begin
        _EVAL_2329 <= _EVAL_1492;
      end else begin
        _EVAL_2329 <= _EVAL_1179;
      end
    end else begin
      _EVAL_2329 <= _EVAL_1179;
    end
    if (_EVAL_83) begin
      _EVAL_2331 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_726) begin
        if (_EVAL_2246) begin
          _EVAL_2331 <= _EVAL_672;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_2342 <= 6'h0;
    end else begin
      _EVAL_2342 <= _EVAL_302[5:0];
    end
    if (_EVAL_83) begin
      _EVAL_2352 <= 3'h0;
    end
    if (_EVAL_83) begin
      _EVAL_2366 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_2284) begin
        if (_EVAL_2246) begin
          _EVAL_2366 <= _EVAL_1005;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_2391 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_554) begin
        _EVAL_2391 <= _EVAL_768;
      end
    end
    _EVAL_2418 <= _EVAL_1914[29:0];
    if (_EVAL_83) begin
      _EVAL_2420 <= 1'h0;
    end else begin
      _EVAL_2420 <= _EVAL_497;
    end
    if (_EVAL_1065) begin
      if (_EVAL_1715) begin
        _EVAL_2422 <= _EVAL_906;
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_726) begin
        if (_EVAL_2246) begin
          _EVAL_2425 <= _EVAL_638;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_2426 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_2192) begin
        _EVAL_2426 <= _EVAL_1785;
      end
    end
    if (_EVAL_83) begin
      _EVAL_2451 <= 1'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_299) begin
        _EVAL_2451 <= _EVAL_912;
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_554) begin
        _EVAL_2461 <= _EVAL_1907;
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_1588) begin
        if (_EVAL_2246) begin
          _EVAL_2465 <= _EVAL_638;
        end
      end
    end
    if (_EVAL_83) begin
      _EVAL_2481 <= 2'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_595) begin
        _EVAL_2481 <= _EVAL_2340;
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_1031) begin
        _EVAL_2492 <= _EVAL_2490;
      end
    end
    if (_EVAL_1065) begin
      if (_EVAL_1897) begin
        _EVAL_2521 <= _EVAL_2323;
      end
    end
    if (_EVAL_83) begin
      _EVAL_2532 <= 1'h0;
    end
  end
  always @(posedge _EVAL_41) begin
    if (_EVAL_83) begin
      _EVAL_834 <= 1'h0;
    end else if (_EVAL_2120) begin
      _EVAL_834 <= 1'h0;
    end else begin
      _EVAL_834 <= _EVAL_213;
    end
    if (_EVAL_83) begin
      _EVAL_2248 <= 6'h0;
    end else begin
      _EVAL_2248 <= _EVAL_1279[5:0];
    end
    if (_EVAL_83) begin
      _EVAL_2550 <= 58'h0;
    end else if (_EVAL_1065) begin
      if (_EVAL_1119) begin
        _EVAL_2550 <= _EVAL_1692;
      end else if (_EVAL_1041) begin
        _EVAL_2550 <= _EVAL_682;
      end else begin
        _EVAL_2550 <= _EVAL_418;
      end
    end else begin
      _EVAL_2550 <= _EVAL_418;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_227 = _RAND_0[29:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_237 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_245 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_280 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_282 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_312 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_313 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_359 = _RAND_7[29:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_365 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_366 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_370 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_385 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_387 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_395 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_417 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_454 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_460 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _EVAL_461 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  _EVAL_498 = _RAND_18[5:0];
  _RAND_19 = {1{`RANDOM}};
  _EVAL_500 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  _EVAL_540 = _RAND_20[29:0];
  _RAND_21 = {1{`RANDOM}};
  _EVAL_611 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  _EVAL_617 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  _EVAL_630 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  _EVAL_647 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  _EVAL_665 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  _EVAL_668 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  _EVAL_679 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  _EVAL_689 = _RAND_28[11:0];
  _RAND_29 = {1{`RANDOM}};
  _EVAL_722 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  _EVAL_740 = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  _EVAL_741 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  _EVAL_743 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  _EVAL_767 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  _EVAL_793 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  _EVAL_795 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  _EVAL_799 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  _EVAL_804 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  _EVAL_820 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  _EVAL_834 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  _EVAL_855 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  _EVAL_872 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  _EVAL_877 = _RAND_42[1:0];
  _RAND_43 = {1{`RANDOM}};
  _EVAL_890 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  _EVAL_891 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  _EVAL_905 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  _EVAL_937 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  _EVAL_949 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  _EVAL_962 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  _EVAL_965 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  _EVAL_985 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  _EVAL_1001 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  _EVAL_1017 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  _EVAL_1027 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  _EVAL_1032 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  _EVAL_1059 = _RAND_55[1:0];
  _RAND_56 = {2{`RANDOM}};
  _EVAL_1062 = _RAND_56[57:0];
  _RAND_57 = {1{`RANDOM}};
  _EVAL_1070 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  _EVAL_1075 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  _EVAL_1113 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  _EVAL_1120 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  _EVAL_1155 = _RAND_61[29:0];
  _RAND_62 = {1{`RANDOM}};
  _EVAL_1159 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  _EVAL_1161 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  _EVAL_1187 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  _EVAL_1206 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  _EVAL_1212 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  _EVAL_1213 = _RAND_67[26:0];
  _RAND_68 = {1{`RANDOM}};
  _EVAL_1217 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  _EVAL_1227 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  _EVAL_1229 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  _EVAL_1231 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  _EVAL_1280 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  _EVAL_1300 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  _EVAL_1302 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  _EVAL_1306 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  _EVAL_1326 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  _EVAL_1334 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  _EVAL_1344 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  _EVAL_1357 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  _EVAL_1383 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  _EVAL_1399 = _RAND_81[0:0];
  _RAND_82 = {2{`RANDOM}};
  _EVAL_1439 = _RAND_82[33:0];
  _RAND_83 = {1{`RANDOM}};
  _EVAL_1463 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  _EVAL_1478 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  _EVAL_1496 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  _EVAL_1504 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  _EVAL_1505 = _RAND_87[5:0];
  _RAND_88 = {1{`RANDOM}};
  _EVAL_1511 = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  _EVAL_1525 = _RAND_89[1:0];
  _RAND_90 = {1{`RANDOM}};
  _EVAL_1534 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  _EVAL_1541 = _RAND_91[1:0];
  _RAND_92 = {1{`RANDOM}};
  _EVAL_1545 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  _EVAL_1557 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  _EVAL_1595 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  _EVAL_1618 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  _EVAL_1620 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  _EVAL_1633 = _RAND_97[1:0];
  _RAND_98 = {1{`RANDOM}};
  _EVAL_1657 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  _EVAL_1672 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  _EVAL_1694 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  _EVAL_1696 = _RAND_101[1:0];
  _RAND_102 = {1{`RANDOM}};
  _EVAL_1733 = _RAND_102[4:0];
  _RAND_103 = {1{`RANDOM}};
  _EVAL_1738 = _RAND_103[1:0];
  _RAND_104 = {1{`RANDOM}};
  _EVAL_1757 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  _EVAL_1761 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  _EVAL_1788 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  _EVAL_1796 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  _EVAL_1813 = _RAND_108[29:0];
  _RAND_109 = {2{`RANDOM}};
  _EVAL_1817 = _RAND_109[33:0];
  _RAND_110 = {1{`RANDOM}};
  _EVAL_1828 = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  _EVAL_1847 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  _EVAL_1849 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  _EVAL_1858 = _RAND_113[1:0];
  _RAND_114 = {1{`RANDOM}};
  _EVAL_1867 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  _EVAL_1870 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  _EVAL_1878 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  _EVAL_1910 = _RAND_117[29:0];
  _RAND_118 = {1{`RANDOM}};
  _EVAL_1918 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  _EVAL_1920 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  _EVAL_1935 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  _EVAL_1947 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  _EVAL_1955 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  _EVAL_1959 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  _EVAL_1967 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  _EVAL_1978 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  _EVAL_2042 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  _EVAL_2069 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  _EVAL_2075 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  _EVAL_2082 = _RAND_129[1:0];
  _RAND_130 = {1{`RANDOM}};
  _EVAL_2099 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  _EVAL_2128 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  _EVAL_2149 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  _EVAL_2159 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  _EVAL_2163 = _RAND_134[1:0];
  _RAND_135 = {1{`RANDOM}};
  _EVAL_2174 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  _EVAL_2182 = _RAND_136[1:0];
  _RAND_137 = {1{`RANDOM}};
  _EVAL_2185 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  _EVAL_2245 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  _EVAL_2248 = _RAND_139[5:0];
  _RAND_140 = {1{`RANDOM}};
  _EVAL_2262 = _RAND_140[29:0];
  _RAND_141 = {1{`RANDOM}};
  _EVAL_2272 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  _EVAL_2297 = _RAND_142[1:0];
  _RAND_143 = {1{`RANDOM}};
  _EVAL_2301 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  _EVAL_2315 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  _EVAL_2329 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  _EVAL_2331 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  _EVAL_2342 = _RAND_147[5:0];
  _RAND_148 = {1{`RANDOM}};
  _EVAL_2352 = _RAND_148[2:0];
  _RAND_149 = {1{`RANDOM}};
  _EVAL_2366 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  _EVAL_2391 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  _EVAL_2418 = _RAND_151[29:0];
  _RAND_152 = {1{`RANDOM}};
  _EVAL_2420 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  _EVAL_2422 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  _EVAL_2425 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  _EVAL_2426 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  _EVAL_2451 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  _EVAL_2461 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  _EVAL_2465 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  _EVAL_2481 = _RAND_159[1:0];
  _RAND_160 = {1{`RANDOM}};
  _EVAL_2492 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  _EVAL_2521 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  _EVAL_2532 = _RAND_162[0:0];
  _RAND_163 = {2{`RANDOM}};
  _EVAL_2550 = _RAND_163[57:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
