//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_5_assert(
  input         _EVAL,
  input         _EVAL_0,
  input  [3:0]  _EVAL_1,
  input         _EVAL_2,
  input  [3:0]  _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  input  [1:0]  _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input  [3:0]  _EVAL_11,
  input  [31:0] _EVAL_12,
  input  [2:0]  _EVAL_13,
  input  [3:0]  _EVAL_14,
  input  [2:0]  _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  input  [3:0]  _EVAL_18
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire [32:0] _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire [6:0] _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire [5:0] _EVAL_35;
  wire  _EVAL_36;
  wire [31:0] _EVAL_37;
  wire [7:0] _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire [8:0] _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire [22:0] _EVAL_48;
  wire [7:0] _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_54;
  wire [15:0] _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire [32:0] _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  reg [8:0] _EVAL_67;
  wire [31:0] _EVAL_68;
  wire [7:0] _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire [8:0] _EVAL_75;
  wire [32:0] _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire [32:0] _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire [5:0] _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire [15:0] _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire [32:0] _EVAL_112;
  wire [5:0] _EVAL_113;
  wire  _EVAL_114;
  reg [2:0] _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire [31:0] _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_126;
  wire [3:0] _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire [32:0] _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire [2:0] _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire [6:0] _EVAL_149;
  wire [32:0] _EVAL_150;
  wire [32:0] _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire [7:0] _EVAL_156;
  wire  _EVAL_157;
  wire [32:0] _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire [32:0] _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire [32:0] _EVAL_174;
  wire  _EVAL_175;
  reg [3:0] _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire [15:0] _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire [15:0] _EVAL_187;
  wire  _EVAL_188;
  wire [3:0] _EVAL_189;
  wire [5:0] _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire [5:0] _EVAL_193;
  wire [32:0] _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire [8:0] _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire [31:0] _EVAL_206;
  wire  _EVAL_207;
  wire [32:0] _EVAL_208;
  wire  _EVAL_209;
  reg [1:0] _EVAL_210;
  wire [8:0] _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  reg [2:0] _EVAL_215;
  wire  _EVAL_216;
  wire [2:0] _EVAL_217;
  wire  _EVAL_218;
  wire [6:0] _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  reg [5:0] _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire [1:0] _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_245;
  reg [3:0] _EVAL_246;
  wire  _EVAL_247;
  reg  _EVAL_248;
  wire [31:0] _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire [8:0] _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  wire [1:0] _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire [8:0] _EVAL_262;
  reg [2:0] _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire [32:0] _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire [6:0] _EVAL_271;
  wire  _EVAL_272;
  reg [3:0] _EVAL_273;
  wire  _EVAL_274;
  wire [22:0] _EVAL_275;
  reg [5:0] _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire [8:0] _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire [32:0] _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  reg [5:0] _EVAL_286;
  wire [5:0] _EVAL_287;
  wire  _EVAL_288;
  wire [3:0] _EVAL_289;
  wire  _EVAL_290;
  wire [31:0] _EVAL_291;
  reg [31:0] _EVAL_292;
  wire  _EVAL_293;
  wire [32:0] _EVAL_294;
  wire  _EVAL_295;
  wire [32:0] _EVAL_296;
  wire  _EVAL_297;
  wire [31:0] _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire [31:0] _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_304;
  wire  _EVAL_305;
  reg [3:0] _EVAL_306;
  wire [32:0] _EVAL_307;
  wire  _EVAL_308;
  wire  _EVAL_310;
  wire  _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_315;
  wire [8:0] _EVAL_317;
  reg [31:0] _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_320;
  wire  _EVAL_321;
  wire [32:0] _EVAL_322;
  wire  _EVAL_323;
  wire [32:0] _EVAL_324;
  wire  _EVAL_325;
  wire  _EVAL_327;
  wire [32:0] _EVAL_328;
  wire [31:0] _EVAL_329;
  wire  _EVAL_330;
  wire  _EVAL_331;
  wire  _EVAL_332;
  wire  _EVAL_333;
  wire  _EVAL_334;
  wire  _EVAL_335;
  wire  _EVAL_336;
  wire  _EVAL_337;
  wire  _EVAL_338;
  reg [5:0] _EVAL_339;
  wire  _EVAL_340;
  wire  _EVAL_341;
  wire  _EVAL_342;
  wire  _EVAL_344;
  wire [31:0] _EVAL_345;
  wire  _EVAL_346;
  wire [3:0] _EVAL_347;
  wire [32:0] _EVAL_348;
  wire  _EVAL_349;
  wire  _EVAL_350;
  wire  _EVAL_351;
  wire  _EVAL_352;
  wire  _EVAL_353;
  wire  _EVAL_354;
  wire  _EVAL_355;
  wire  _EVAL_356;
  wire  _EVAL_357;
  reg  _EVAL_358;
  wire  _EVAL_359;
  wire  _EVAL_360;
  wire  _EVAL_361;
  wire  _EVAL_362;
  wire [32:0] _EVAL_363;
  wire  _EVAL_364;
  wire  _EVAL_365;
  wire [32:0] _EVAL_366;
  wire  _EVAL_367;
  wire [32:0] _EVAL_368;
  wire  _EVAL_369;
  wire  _EVAL_370;
  wire  _EVAL_371;
  wire  _EVAL_372;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_61 = _EVAL_5 & _EVAL_270;
  assign _EVAL_78 = _EVAL_242 | _EVAL_17;
  assign _EVAL_27 = ~_EVAL_234;
  assign _EVAL_201 = _EVAL_0 & _EVAL_226;
  assign _EVAL_191 = _EVAL_5 & _EVAL_41;
  assign _EVAL_188 = _EVAL_8 != 2'h2;
  assign _EVAL_307 = $signed(_EVAL_150) & -33'sh10000;
  assign _EVAL_91 = _EVAL_301 | _EVAL_17;
  assign _EVAL_204 = ~_EVAL_78;
  assign _EVAL_348 = _EVAL_294;
  assign _EVAL_38 = ~_EVAL_156;
  assign _EVAL_197 = _EVAL_0 & _EVAL_82;
  assign _EVAL_363 = _EVAL_322;
  assign _EVAL_141 = _EVAL_258[1];
  assign _EVAL_151 = {1'b0,$signed(_EVAL_68)};
  assign _EVAL_366 = _EVAL_328;
  assign _EVAL_126 = _EVAL_228 | _EVAL_17;
  assign _EVAL_42 = _EVAL_262 >> _EVAL_1;
  assign _EVAL_69 = _EVAL_275[7:0];
  assign _EVAL_72 = _EVAL_5 & _EVAL_50;
  assign _EVAL_291 = {{24'd0}, _EVAL_49};
  assign _EVAL_120 = _EVAL_148 | _EVAL_207;
  assign _EVAL_196 = _EVAL_172 & _EVAL_220;
  assign _EVAL_99 = _EVAL_13 == 3'h5;
  assign _EVAL_199 = _EVAL_0 & _EVAL_247;
  assign _EVAL_131 = _EVAL_186 | _EVAL_58;
  assign _EVAL_136 = $signed(_EVAL_158) & -33'sh4000;
  assign _EVAL_274 = _EVAL_295 | _EVAL_164;
  assign _EVAL_119 = _EVAL_289 == 4'h0;
  assign _EVAL_347 = ~_EVAL_189;
  assign _EVAL_242 = _EVAL == _EVAL_248;
  assign _EVAL_237 = _EVAL_251 | _EVAL_17;
  assign _EVAL_161 = ~_EVAL_236;
  assign _EVAL_182 = _EVAL_3[0];
  assign _EVAL_146 = 4'h2 == _EVAL_3;
  assign _EVAL_171 = ~_EVAL_320;
  assign _EVAL_156 = _EVAL_48[7:0];
  assign _EVAL_349 = _EVAL_167 | _EVAL_17;
  assign _EVAL_353 = _EVAL_147 | _EVAL_133;
  assign _EVAL_325 = _EVAL_259 | _EVAL_277;
  assign _EVAL_82 = ~_EVAL_23;
  assign _EVAL_149 = _EVAL_339 - 6'h1;
  assign _EVAL_225 = ~_EVAL_238;
  assign _EVAL_142 = _EVAL_12 == _EVAL_318;
  assign _EVAL_84 = _EVAL_89 & _EVAL_107;
  assign _EVAL_113 = _EVAL_32[5:0];
  assign _EVAL_64 = ~_EVAL_288;
  assign _EVAL_56 = 16'h1 << _EVAL_1;
  assign _EVAL_202 = _EVAL_67 | _EVAL_253;
  assign _EVAL_46 = _EVAL_13 == 3'h1;
  assign _EVAL_360 = _EVAL_127 == 4'h0;
  assign _EVAL_194 = $signed(_EVAL_296) & -33'sh1000;
  assign _EVAL_65 = ~_EVAL_152;
  assign _EVAL_337 = _EVAL_25 & _EVAL_173;
  assign _EVAL_183 = ~_EVAL_29;
  assign _EVAL_205 = _EVAL_13[0];
  assign _EVAL_338 = _EVAL_8 == 2'h0;
  assign _EVAL_344 = _EVAL_28 | _EVAL_17;
  assign _EVAL_362 = ~_EVAL_43;
  assign _EVAL_195 = _EVAL_14 == _EVAL_306;
  assign _EVAL_342 = ~_EVAL_178;
  assign _EVAL_81 = _EVAL_1 == _EVAL_176;
  assign _EVAL_354 = plusarg_reader_out == 32'h0;
  assign _EVAL_123 = _EVAL_25 & _EVAL_288;
  assign _EVAL_66 = _EVAL_216 | _EVAL_17;
  assign _EVAL_293 = _EVAL_5 & _EVAL_64;
  assign _EVAL_86 = _EVAL_119 | _EVAL_17;
  assign _EVAL_167 = ~_EVAL_10;
  assign _EVAL_209 = _EVAL_3 <= 4'h8;
  assign _EVAL_40 = ~_EVAL_355;
  assign _EVAL_350 = ~_EVAL_237;
  assign _EVAL_303 = _EVAL_249 == 32'h0;
  assign _EVAL_238 = _EVAL_264 | _EVAL_17;
  assign _EVAL_31 = _EVAL_200 | _EVAL_87;
  assign _EVAL_179 = ~_EVAL_284;
  assign _EVAL_47 = ~_EVAL_104;
  assign _EVAL_203 = _EVAL_15 == 3'h0;
  assign _EVAL_370 = _EVAL_172 & _EVAL_311;
  assign _EVAL_132 = _EVAL_3 <= 4'h6;
  assign _EVAL_313 = _EVAL_217 <= 3'h6;
  assign _EVAL_208 = {1'b0,$signed(_EVAL_345)};
  assign _EVAL_103 = _EVAL_7 <= 3'h2;
  assign _EVAL_45 = _EVAL_132 & _EVAL_214;
  assign _EVAL_290 = _EVAL_5 & _EVAL_124;
  assign _EVAL_30 = _EVAL_371 | _EVAL_58;
  assign _EVAL_122 = _EVAL_8 <= 2'h2;
  assign _EVAL_87 = _EVAL_14 == 4'h8;
  assign _EVAL_287 = _EVAL_149[5:0];
  assign _EVAL_147 = _EVAL_70 | _EVAL_280;
  assign _EVAL_264 = _EVAL_7 <= 3'h1;
  assign _EVAL_260 = _EVAL_15[2];
  assign _EVAL_52 = _EVAL_5 & _EVAL_85;
  assign _EVAL_312 = _EVAL_5 & _EVAL_334;
  assign _EVAL_135 = _EVAL_132 & _EVAL_231;
  assign _EVAL_184 = ~_EVAL_154;
  assign _EVAL_323 = _EVAL_103 | _EVAL_17;
  assign _EVAL_240 = _EVAL_15 == 3'h3;
  assign _EVAL_166 = ~_EVAL_321;
  assign _EVAL_98 = _EVAL_357 & _EVAL_222;
  assign _EVAL_112 = {1'b0,$signed(_EVAL_12)};
  assign _EVAL_315 = _EVAL_147 | _EVAL_196;
  assign _EVAL_158 = {1'b0,$signed(_EVAL_118)};
  assign _EVAL_231 = _EVAL_351 | _EVAL_164;
  assign _EVAL_294 = $signed(_EVAL_268) & -33'sh4000;
  assign _EVAL_297 = ~_EVAL_130;
  assign _EVAL_213 = _EVAL_25 | _EVAL_254;
  assign _EVAL_70 = _EVAL_3 >= 4'h2;
  assign _EVAL_227 = ~_EVAL_314;
  assign _EVAL_174 = {1'b0,$signed(_EVAL_37)};
  assign _EVAL_261 = _EVAL_14[3];
  assign _EVAL_74 = _EVAL_142 | _EVAL_17;
  assign _EVAL_29 = _EVAL_120 | _EVAL_17;
  assign _EVAL_89 = _EVAL_254 & _EVAL_93;
  assign _EVAL_157 = _EVAL_0 & _EVAL_102;
  assign _EVAL_285 = ~_EVAL_305;
  assign _EVAL_39 = _EVAL_13 == _EVAL_115;
  assign _EVAL_319 = _EVAL_356 | _EVAL_17;
  assign _EVAL_280 = _EVAL_141 & _EVAL_47;
  assign _EVAL_336 = _EVAL_209 & _EVAL_116;
  assign _EVAL_19 = _EVAL_12[0];
  assign _EVAL_178 = _EVAL_97 | _EVAL_17;
  assign _EVAL_359 = _EVAL_222 | _EVAL_17;
  assign _EVAL_255 = _EVAL_5 & _EVAL_240;
  assign _EVAL_58 = $signed(_EVAL_348) == 33'sh0;
  assign _EVAL_137 = ~_EVAL_20;
  assign _EVAL_270 = _EVAL_15 == 3'h2;
  assign _EVAL_104 = _EVAL_12[1];
  assign _EVAL_24 = ~_EVAL_71;
  assign _EVAL_259 = _EVAL_131 | _EVAL_304;
  assign _EVAL_296 = {1'b0,$signed(_EVAL_206)};
  assign _EVAL_145 = _EVAL_325 | _EVAL_162;
  assign _EVAL_200 = _EVAL_346 & _EVAL_313;
  assign _EVAL_90 = ~_EVAL_17;
  assign _EVAL_155 = _EVAL_2 == _EVAL_358;
  assign _EVAL_159 = ~_EVAL_367;
  assign _EVAL_109 = ~_EVAL_163;
  assign _EVAL_265 = _EVAL_54 | _EVAL_17;
  assign _EVAL_59 = _EVAL_185 | _EVAL_17;
  assign _EVAL_308 = _EVAL_332 | _EVAL_17;
  assign _EVAL_63 = _EVAL_7 == 3'h0;
  assign _EVAL_76 = $signed(_EVAL_208) & -33'sh400000;
  assign _EVAL_219 = _EVAL_276 - 6'h1;
  assign _EVAL_321 = _EVAL_297 | _EVAL_17;
  assign _EVAL_224 = _EVAL_295 | _EVAL_162;
  assign _EVAL_311 = _EVAL_104 & _EVAL_245;
  assign _EVAL_212 = ~_EVAL_308;
  assign _EVAL_162 = $signed(_EVAL_366) == 33'sh0;
  assign _EVAL_295 = _EVAL_241 | _EVAL_277;
  assign _EVAL_214 = _EVAL_162 | _EVAL_252;
  assign _EVAL_150 = {1'b0,$signed(_EVAL_302)};
  assign _EVAL_257 = ~_EVAL_218;
  assign _EVAL_334 = _EVAL_15 == 3'h1;
  assign _EVAL_310 = _EVAL_360 | _EVAL_17;
  assign _EVAL_320 = _EVAL_192 | _EVAL_17;
  assign _EVAL_129 = _EVAL_254 & _EVAL_23;
  assign _EVAL_365 = _EVAL_145 | _EVAL_164;
  assign _EVAL_198 = _EVAL_266 | _EVAL_17;
  assign _EVAL_153 = _EVAL_165 | _EVAL_364;
  assign _EVAL_364 = _EVAL_172 & _EVAL_143;
  assign _EVAL_164 = $signed(_EVAL_80) == 33'sh0;
  assign _EVAL_211 = _EVAL_67 >> _EVAL_14;
  assign _EVAL_367 = _EVAL_250 | _EVAL_17;
  assign _EVAL_187 = _EVAL_84 ? _EVAL_56 : 16'h0;
  assign _EVAL_271 = _EVAL_286 - 6'h1;
  assign _EVAL_324 = _EVAL_307;
  assign _EVAL_278 = ~_EVAL_106;
  assign _EVAL_88 = _EVAL_111 & _EVAL_96;
  assign _EVAL_356 = _EVAL_13 <= 3'h6;
  assign _EVAL_160 = _EVAL_47 & _EVAL_245;
  assign _EVAL_21 = ~_EVAL_349;
  assign _EVAL_277 = $signed(_EVAL_368) == 33'sh0;
  assign _EVAL_118 = _EVAL_12 ^ 32'h80000000;
  assign _EVAL_23 = _EVAL_276 == 6'h0;
  assign _EVAL_140 = _EVAL_1[2:0];
  assign _EVAL_333 = _EVAL_11 >= 4'h2;
  assign _EVAL_371 = $signed(_EVAL_363) == 33'sh0;
  assign _EVAL_268 = {1'b0,$signed(_EVAL_329)};
  assign _EVAL_28 = _EVAL_3 == _EVAL_246;
  assign _EVAL_322 = $signed(_EVAL_112) & -33'sh5000;
  assign _EVAL_172 = _EVAL_258[0];
  assign _EVAL_96 = _EVAL_51 & _EVAL_365;
  assign _EVAL_258 = _EVAL_233 | 2'h1;
  assign _EVAL_335 = _EVAL_140 <= 3'h6;
  assign _EVAL_275 = 23'hff << _EVAL_3;
  assign _EVAL_80 = _EVAL_136;
  assign _EVAL_372 = _EVAL_39 | _EVAL_17;
  assign _EVAL_25 = _EVAL_16 & _EVAL_5;
  assign _EVAL_169 = $signed(_EVAL_151) & -33'sh2000;
  assign _EVAL_173 = _EVAL_286 == 6'h0;
  assign _EVAL_304 = $signed(_EVAL_324) == 33'sh0;
  assign _EVAL_193 = _EVAL_219[5:0];
  assign _EVAL_328 = $signed(_EVAL_174) & -33'sh2000;
  assign _EVAL_165 = _EVAL_70 | _EVAL_138;
  assign _EVAL_134 = _EVAL_88 | _EVAL_17;
  assign _EVAL_189 = {_EVAL_153,_EVAL_341,_EVAL_315,_EVAL_353};
  assign _EVAL_108 = _EVAL_340 & _EVAL_87;
  assign _EVAL_221 = _EVAL_269 & _EVAL_335;
  assign _EVAL_60 = _EVAL_292 + 32'h1;
  assign _EVAL_148 = _EVAL_362 | _EVAL_354;
  assign _EVAL_51 = _EVAL_3 <= 4'h2;
  assign _EVAL_245 = ~_EVAL_19;
  assign _EVAL_152 = _EVAL_31 | _EVAL_17;
  assign _EVAL_298 = _EVAL_60[31:0];
  assign _EVAL_85 = _EVAL_15 == 3'h5;
  assign _EVAL_105 = _EVAL_337 ? _EVAL_180 : 16'h0;
  assign _EVAL_368 = _EVAL_76;
  assign _EVAL_54 = _EVAL_336 | _EVAL_139;
  assign _EVAL_226 = _EVAL_13 == 3'h6;
  assign _EVAL_314 = _EVAL_283 | _EVAL_17;
  assign _EVAL_247 = _EVAL_13 == 3'h4;
  assign _EVAL_43 = |_EVAL_67;
  assign _EVAL_111 = _EVAL_146 & _EVAL_200;
  assign _EVAL_48 = 23'hff << _EVAL_11;
  assign _EVAL_130 = _EVAL_211[0];
  assign _EVAL_262 = _EVAL_253 | _EVAL_67;
  assign _EVAL_357 = _EVAL_51 & _EVAL_200;
  assign _EVAL_26 = _EVAL_169;
  assign _EVAL_101 = ~_EVAL_73;
  assign _EVAL_41 = _EVAL_15 == 3'h6;
  assign _EVAL_94 = _EVAL_38[7:2];
  assign _EVAL_49 = ~_EVAL_69;
  assign _EVAL_57 = ~_EVAL_59;
  assign _EVAL_332 = _EVAL_221 | _EVAL_117;
  assign _EVAL_352 = ~_EVAL_331;
  assign _EVAL_110 = ~_EVAL_260;
  assign _EVAL_32 = _EVAL_230 - 6'h1;
  assign _EVAL_229 = _EVAL_336 | _EVAL_45;
  assign _EVAL_330 = ~_EVAL_323;
  assign _EVAL_37 = _EVAL_12 ^ 32'h20000000;
  assign _EVAL_207 = _EVAL_292 < plusarg_reader_out;
  assign _EVAL_253 = _EVAL_105[8:0];
  assign _EVAL_92 = _EVAL_0 & _EVAL_46;
  assign _EVAL_33 = _EVAL_0 & _EVAL_99;
  assign _EVAL_216 = _EVAL_7 <= 3'h4;
  assign _EVAL_345 = _EVAL_12 ^ 32'hc000000;
  assign _EVAL_282 = _EVAL_194;
  assign _EVAL_228 = _EVAL_369 | _EVAL_256;
  assign _EVAL_124 = _EVAL_15 == 3'h4;
  assign _EVAL_100 = ~_EVAL_223;
  assign _EVAL_272 = ~_EVAL_310;
  assign _EVAL_369 = _EVAL_253 != _EVAL_279;
  assign _EVAL_181 = ~_EVAL_91;
  assign _EVAL_234 = _EVAL_77 | _EVAL_17;
  assign _EVAL_340 = 4'h6 == _EVAL_3;
  assign _EVAL_251 = _EVAL_7 != 3'h0;
  assign _EVAL_250 = _EVAL_18 == _EVAL_189;
  assign _EVAL_116 = $signed(_EVAL_282) == 33'sh0;
  assign _EVAL_284 = _EVAL_81 | _EVAL_17;
  assign _EVAL_163 = _EVAL_333 | _EVAL_17;
  assign _EVAL_79 = ~_EVAL_232;
  assign _EVAL_128 = ~_EVAL_319;
  assign _EVAL_127 = _EVAL_18 & _EVAL_347;
  assign _EVAL_355 = _EVAL_170 | _EVAL_17;
  assign _EVAL_243 = _EVAL_13 == 3'h2;
  assign _EVAL_222 = _EVAL_336 | _EVAL_135;
  assign _EVAL_206 = _EVAL_12 ^ 32'h3000;
  assign _EVAL_267 = ~_EVAL_66;
  assign _EVAL_305 = _EVAL_98 | _EVAL_17;
  assign _EVAL_97 = _EVAL_357 | _EVAL_108;
  assign _EVAL_351 = _EVAL_224 | _EVAL_252;
  assign _EVAL_317 = ~_EVAL_279;
  assign _EVAL_233 = 2'h1 << _EVAL_182;
  assign _EVAL_22 = ~_EVAL_265;
  assign _EVAL_168 = ~_EVAL_359;
  assign _EVAL_107 = ~_EVAL_226;
  assign _EVAL_180 = 16'h1 << _EVAL_14;
  assign _EVAL_223 = _EVAL_229 | _EVAL_17;
  assign _EVAL_36 = _EVAL_188 | _EVAL_17;
  assign _EVAL_114 = _EVAL_5 & _EVAL_203;
  assign _EVAL_192 = _EVAL_7 <= 3'h3;
  assign _EVAL_218 = _EVAL_122 | _EVAL_17;
  assign _EVAL_300 = ~_EVAL_86;
  assign _EVAL_331 = _EVAL_361 | _EVAL_17;
  assign _EVAL_269 = ~_EVAL_62;
  assign _EVAL_139 = _EVAL_132 & _EVAL_274;
  assign _EVAL_232 = _EVAL_338 | _EVAL_17;
  assign _EVAL_175 = ~_EVAL_134;
  assign _EVAL_236 = _EVAL_195 | _EVAL_17;
  assign _EVAL_289 = ~_EVAL_18;
  assign _EVAL_71 = _EVAL_303 | _EVAL_17;
  assign _EVAL_154 = _EVAL_70 | _EVAL_17;
  assign _EVAL_241 = _EVAL_30 | _EVAL_304;
  assign _EVAL_177 = ~_EVAL_372;
  assign _EVAL_95 = |_EVAL_253;
  assign _EVAL_117 = _EVAL_1 == 4'h8;
  assign _EVAL_302 = _EVAL_12 ^ 32'h2000000;
  assign _EVAL_50 = _EVAL_15 == 3'h7;
  assign _EVAL_121 = _EVAL_7 == _EVAL_263;
  assign _EVAL_102 = _EVAL_13 == 3'h0;
  assign _EVAL_329 = _EVAL_12 ^ 32'h1800000;
  assign _EVAL_327 = ~_EVAL_126;
  assign _EVAL_252 = $signed(_EVAL_26) == 33'sh0;
  assign _EVAL_185 = _EVAL_11 == _EVAL_273;
  assign _EVAL_279 = _EVAL_187[8:0];
  assign _EVAL_75 = _EVAL_202 & _EVAL_317;
  assign _EVAL_346 = ~_EVAL_261;
  assign _EVAL_73 = _EVAL_121 | _EVAL_17;
  assign _EVAL_62 = _EVAL_1[3];
  assign _EVAL_34 = _EVAL_0 & _EVAL_243;
  assign _EVAL_235 = ~_EVAL_36;
  assign _EVAL_68 = _EVAL_12 ^ 32'h40000000;
  assign _EVAL_93 = _EVAL_230 == 6'h0;
  assign _EVAL_220 = _EVAL_47 & _EVAL_19;
  assign _EVAL_256 = ~_EVAL_95;
  assign _EVAL_170 = _EVAL_361 | _EVAL_10;
  assign _EVAL_144 = ~_EVAL_344;
  assign _EVAL_254 = _EVAL_6 & _EVAL_0;
  assign _EVAL_106 = _EVAL_63 | _EVAL_17;
  assign _EVAL_301 = _EVAL_42[0];
  assign _EVAL_249 = _EVAL_12 & _EVAL_291;
  assign _EVAL_35 = _EVAL_49[7:2];
  assign _EVAL_299 = ~_EVAL_198;
  assign _EVAL_143 = _EVAL_104 & _EVAL_19;
  assign _EVAL_20 = _EVAL_155 | _EVAL_17;
  assign _EVAL_361 = ~_EVAL_2;
  assign _EVAL_283 = ~_EVAL_9;
  assign _EVAL_217 = _EVAL_14[2:0];
  assign _EVAL_281 = ~_EVAL_74;
  assign _EVAL_190 = _EVAL_271[5:0];
  assign _EVAL_138 = _EVAL_141 & _EVAL_104;
  assign _EVAL_186 = _EVAL_371 | _EVAL_116;
  assign _EVAL_133 = _EVAL_172 & _EVAL_160;
  assign _EVAL_77 = _EVAL_8 == _EVAL_210;
  assign _EVAL_288 = _EVAL_339 == 6'h0;
  assign _EVAL_341 = _EVAL_165 | _EVAL_370;
  assign _EVAL_266 = _EVAL_15 == _EVAL_215;
  always @(posedge _EVAL_4) begin
    if (_EVAL_17) begin
      _EVAL_67 <= 9'h0;
    end else begin
      _EVAL_67 <= _EVAL_75;
    end
    if (_EVAL_129) begin
      _EVAL_115 <= _EVAL_13;
    end
    if (_EVAL_129) begin
      _EVAL_176 <= _EVAL_1;
    end
    if (_EVAL_129) begin
      _EVAL_210 <= _EVAL_8;
    end
    if (_EVAL_123) begin
      _EVAL_215 <= _EVAL_15;
    end
    if (_EVAL_17) begin
      _EVAL_230 <= 6'h0;
    end else if (_EVAL_254) begin
      if (_EVAL_93) begin
        if (_EVAL_205) begin
          _EVAL_230 <= _EVAL_94;
        end else begin
          _EVAL_230 <= 6'h0;
        end
      end else begin
        _EVAL_230 <= _EVAL_113;
      end
    end
    if (_EVAL_123) begin
      _EVAL_246 <= _EVAL_3;
    end
    if (_EVAL_129) begin
      _EVAL_248 <= _EVAL;
    end
    if (_EVAL_123) begin
      _EVAL_263 <= _EVAL_7;
    end
    if (_EVAL_129) begin
      _EVAL_273 <= _EVAL_11;
    end
    if (_EVAL_17) begin
      _EVAL_276 <= 6'h0;
    end else if (_EVAL_254) begin
      if (_EVAL_23) begin
        if (_EVAL_205) begin
          _EVAL_276 <= _EVAL_94;
        end else begin
          _EVAL_276 <= 6'h0;
        end
      end else begin
        _EVAL_276 <= _EVAL_193;
      end
    end
    if (_EVAL_17) begin
      _EVAL_286 <= 6'h0;
    end else if (_EVAL_25) begin
      if (_EVAL_173) begin
        if (_EVAL_110) begin
          _EVAL_286 <= _EVAL_35;
        end else begin
          _EVAL_286 <= 6'h0;
        end
      end else begin
        _EVAL_286 <= _EVAL_190;
      end
    end
    if (_EVAL_17) begin
      _EVAL_292 <= 32'h0;
    end else if (_EVAL_213) begin
      _EVAL_292 <= 32'h0;
    end else begin
      _EVAL_292 <= _EVAL_298;
    end
    if (_EVAL_123) begin
      _EVAL_306 <= _EVAL_14;
    end
    if (_EVAL_123) begin
      _EVAL_318 <= _EVAL_12;
    end
    if (_EVAL_17) begin
      _EVAL_339 <= 6'h0;
    end else if (_EVAL_25) begin
      if (_EVAL_288) begin
        if (_EVAL_110) begin
          _EVAL_339 <= _EVAL_35;
        end else begin
          _EVAL_339 <= 6'h0;
        end
      end else begin
        _EVAL_339 <= _EVAL_287;
      end
    end
    if (_EVAL_129) begin
      _EVAL_358 <= _EVAL_2;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_350) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acbd44f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ddabf03d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f28f4218)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_330) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a198419)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2ee27a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39cb7569)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_168) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6a06f0d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71413ee4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e65abe03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7dd6a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_327) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_312 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1663006c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27ecfad2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6570d12e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51452a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bea9af9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(860b197a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61759e0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1927606)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bcd7232d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a293672)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_257) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_257) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71999145)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(316d321c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96a8f8ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_330) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a700aad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_342) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(142a0b19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49712a73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5fc36f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_312 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_342) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_299) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e713341d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_312 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(842d4bf1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a27a1d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96a6a128)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(279626e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbf363d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b36eafa6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_168) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f37a1db4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(386098f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_312 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96a41ab0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_330) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7c017a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_312 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73ae149f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_312 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a732c949)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91f03f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f3cbe8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4416c426)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f74e3fe6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(623ff71d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(820c883f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_352) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98b4f897)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_300) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa8145c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c8112f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_299) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5117f1cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11c1b3cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e2d8891)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_327) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68837a78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_330) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9a6707f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4032f527)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be706813)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(465f0382)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b3b8f56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf21173e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_285) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(618a79b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba77d190)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ef1f833)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e032a96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ded31237)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_300) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(198a2eef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_257) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e4ecef5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(644051d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1981649)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ab73f6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(806b3bd9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4fb18662)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c483e2e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a76b9d19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1523b0e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da9cb69e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_312 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86b78232)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_312 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(588ce535)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b32081e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf21173e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_312 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e68f4b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0826b11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_281) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d33386ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a17ae11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_312 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(229fed1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_352) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_300) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7215a6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb3eea2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_312 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d43d8082)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_199 & _EVAL_257) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7732d1d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f57ce0a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_281) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88c2055)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_312 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a7c0b24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_300) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_337 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ac33c30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_350) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af2dbf1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_285) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_337 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cbe291d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_67 = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_115 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_176 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_210 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_215 = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_230 = _RAND_5[5:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_246 = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_248 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_263 = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_273 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_276 = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_286 = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_292 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_306 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_318 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_339 = _RAND_15[5:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_358 = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
