//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000


module XSquasher #(parameter WIDTH=32) (
  input valid,
  input [WIDTH-1:0] inp,
  output [WIDTH-1:0] outp
);
                    


  reg [WIDTH-1:0] squashed_inp;
  genvar i;
  generate
    for (i=0;i<WIDTH;i++) begin
      always @(inp[i]) begin
        if (inp[i] === 1'b1) squashed_inp[i] = 1'b1;
        else if (inp[i] === 1'b0) squashed_inp[i] = 1'b0;
        else squashed_inp[i] = bit'($random());
      end
    end
  endgenerate
                        
  assign outp = valid ? squashed_inp : inp;
                                         
endmodule
                    