//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_174_assert(
  input  [2:0] _EVAL,
  input        _EVAL_0,
  input  [1:0] _EVAL_1,
  input  [2:0] _EVAL_2,
  input  [8:0] _EVAL_3,
  input        _EVAL_4,
  input        _EVAL_5,
  input        _EVAL_6,
  input        _EVAL_7,
  input        _EVAL_8,
  input        _EVAL_9,
  input        _EVAL_10,
  input  [1:0] _EVAL_11,
  input  [2:0] _EVAL_12,
  input  [3:0] _EVAL_13,
  input        _EVAL_14
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_15;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire [9:0] _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire [1:0] _EVAL_28;
  wire  _EVAL_29;
  reg  _EVAL_30;
  wire [1:0] _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire [31:0] plusarg_reader_out;
  wire [3:0] _EVAL_38;
  reg [2:0] _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_43;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire [1:0] _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire [1:0] _EVAL_52;
  wire  _EVAL_53;
  wire [1:0] _EVAL_54;
  wire [1:0] _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire [9:0] _EVAL_67;
  wire  _EVAL_68;
  wire [3:0] _EVAL_69;
  reg [31:0] _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire [1:0] _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire [8:0] _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire [9:0] _EVAL_87;
  wire  _EVAL_88;
  wire [8:0] _EVAL_89;
  reg  _EVAL_90;
  wire  _EVAL_91;
  reg  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  reg  _EVAL_109;
  wire  _EVAL_110;
  wire [8:0] _EVAL_111;
  wire  _EVAL_112;
  wire [9:0] _EVAL_113;
  wire [8:0] _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire [9:0] _EVAL_117;
  wire [9:0] _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire [31:0] _EVAL_129;
  wire  _EVAL_130;
  wire [8:0] _EVAL_131;
  wire  _EVAL_132;
  wire [32:0] _EVAL_133;
  wire [4:0] _EVAL_134;
  reg [2:0] _EVAL_135;
  wire [8:0] _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  reg [1:0] _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  reg  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire [1:0] _EVAL_158;
  reg [2:0] _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire [1:0] _EVAL_175;
  wire [9:0] _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire [3:0] _EVAL_183;
  wire [9:0] _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire [1:0] _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire [9:0] _EVAL_192;
  wire  _EVAL_193;
  wire [9:0] _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire [9:0] _EVAL_202;
  wire [9:0] _EVAL_204;
  wire [9:0] _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire [9:0] _EVAL_208;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire [3:0] _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_216;
  reg  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire [9:0] _EVAL_229;
  wire  _EVAL_230;
  reg [1:0] _EVAL_231;
  wire [9:0] _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire [9:0] _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire [8:0] _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire [1:0] _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  reg  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire [1:0] _EVAL_265;
  reg [8:0] _EVAL_266;
  wire  _EVAL_267;
  wire [9:0] _EVAL_268;
  wire  _EVAL_269;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_249 = _EVAL_8 & _EVAL_61;
  assign _EVAL_33 = ~_EVAL_37;
  assign _EVAL_149 = _EVAL_141 & _EVAL_110;
  assign _EVAL_232 = {1'b0,$signed(_EVAL_89)};
  assign _EVAL_229 = _EVAL_192;
  assign _EVAL_108 = ~_EVAL_92;
  assign _EVAL_197 = _EVAL_112 | _EVAL_150;
  assign _EVAL_61 = _EVAL_2 == 3'h5;
  assign _EVAL_219 = ~_EVAL_193;
  assign _EVAL_221 = _EVAL_25 & _EVAL_51;
  assign _EVAL_186 = _EVAL_11 == _EVAL_139;
  assign _EVAL_188 = _EVAL_230 | _EVAL_4;
  assign _EVAL_181 = ~_EVAL_132;
  assign _EVAL_45 = _EVAL_13 == _EVAL_183;
  assign _EVAL_173 = _EVAL_5 & _EVAL_46;
  assign _EVAL_97 = _EVAL_1 >= 2'h2;
  assign _EVAL_211 = _EVAL_2 == 3'h6;
  assign _EVAL_83 = _EVAL_182 | _EVAL_4;
  assign _EVAL_115 = ~_EVAL_91;
  assign _EVAL_254 = _EVAL_2 == 3'h1;
  assign _EVAL_31 = 2'h1 << _EVAL_10;
  assign _EVAL_29 = _EVAL_106 & _EVAL_120;
  assign _EVAL_118 = $signed(_EVAL_235) & -10'sh100;
  assign _EVAL_56 = _EVAL_36 | _EVAL_4;
  assign _EVAL_259 = _EVAL_86 | _EVAL_4;
  assign _EVAL_212 = ~_EVAL_13;
  assign _EVAL_162 = _EVAL_45 | _EVAL_4;
  assign _EVAL_89 = _EVAL_3 ^ 9'h58;
  assign _EVAL_95 = _EVAL <= 3'h3;
  assign _EVAL_86 = _EVAL <= 3'h1;
  assign _EVAL_58 = _EVAL_25 & _EVAL_29;
  assign _EVAL_65 = ~_EVAL_130;
  assign _EVAL_246 = ~_EVAL_138;
  assign _EVAL_226 = _EVAL_34 | _EVAL_58;
  assign _EVAL_199 = ~_EVAL_10;
  assign _EVAL_25 = _EVAL_55[0];
  assign _EVAL_17 = ~_EVAL_109;
  assign _EVAL_19 = $signed(_EVAL_205) == 10'sh0;
  assign _EVAL_129 = _EVAL_133[31:0];
  assign _EVAL_43 = _EVAL_150 & _EVAL_255;
  assign _EVAL_16 = _EVAL_112 & _EVAL_108;
  assign _EVAL_37 = _EVAL_12 == 3'h6;
  assign _EVAL_169 = _EVAL_2 == 3'h0;
  assign _EVAL_202 = $signed(_EVAL_176) & -10'sh40;
  assign _EVAL_68 = _EVAL_265[0];
  assign _EVAL_62 = _EVAL_85 | _EVAL_23;
  assign _EVAL_85 = _EVAL_198 | _EVAL_19;
  assign _EVAL_74 = _EVAL_243 & _EVAL_267;
  assign _EVAL_47 = _EVAL_92 - 1'h1;
  assign _EVAL_236 = 2'h2 == _EVAL_1;
  assign _EVAL_75 = _EVAL_134[1:0];
  assign _EVAL_222 = _EVAL <= 3'h2;
  assign _EVAL_154 = ~_EVAL_190;
  assign _EVAL_73 = _EVAL_43 & _EVAL_33;
  assign _EVAL_239 = ~_EVAL_218;
  assign _EVAL_240 = _EVAL_8 & _EVAL_200;
  assign _EVAL_27 = ~_EVAL_56;
  assign _EVAL_195 = _EVAL_62 | _EVAL_40;
  assign _EVAL_193 = _EVAL_252 | _EVAL_4;
  assign _EVAL_71 = _EVAL_149 | _EVAL_4;
  assign _EVAL_51 = _EVAL_243 & _EVAL_120;
  assign _EVAL_185 = _EVAL_12 == _EVAL_135;
  assign _EVAL_269 = _EVAL_25 & _EVAL_74;
  assign _EVAL_18 = ~_EVAL_126;
  assign _EVAL_94 = _EVAL_10 == _EVAL_90;
  assign _EVAL_134 = 5'h3 << _EVAL_1;
  assign _EVAL_223 = _EVAL_30 | _EVAL_168;
  assign _EVAL_142 = ~_EVAL_71;
  assign _EVAL_36 = _EVAL_114 == 9'h0;
  assign _EVAL_124 = ~_EVAL_49;
  assign _EVAL_263 = _EVAL_47[0];
  assign _EVAL_251 = _EVAL_172 | _EVAL_151;
  assign _EVAL_208 = $signed(_EVAL_204) & -10'sh20;
  assign _EVAL_262 = _EVAL_12 == 3'h2;
  assign _EVAL_225 = _EVAL_222 | _EVAL_4;
  assign _EVAL_234 = ~_EVAL_179;
  assign _EVAL_214 = plusarg_reader_out == 32'h0;
  assign _EVAL_133 = _EVAL_70 + 32'h1;
  assign _EVAL_204 = {1'b0,$signed(_EVAL_111)};
  assign _EVAL_224 = _EVAL_8 & _EVAL_211;
  assign _EVAL_28 = _EVAL_109 - 1'h1;
  assign _EVAL_264 = ~_EVAL_81;
  assign _EVAL_218 = _EVAL_97 | _EVAL_4;
  assign _EVAL_164 = $signed(_EVAL_229) == 10'sh0;
  assign _EVAL_245 = _EVAL_8 & _EVAL_122;
  assign _EVAL_172 = _EVAL_234 | _EVAL_214;
  assign _EVAL_123 = _EVAL_171 | _EVAL_4;
  assign _EVAL_50 = ~_EVAL_6;
  assign _EVAL_267 = _EVAL_3[0];
  assign _EVAL_148 = ~_EVAL_83;
  assign _EVAL_117 = _EVAL_113;
  assign _EVAL_136 = _EVAL_3 ^ 9'h44;
  assign _EVAL_171 = _EVAL_212 == 4'h0;
  assign _EVAL_191 = ~_EVAL_76;
  assign _EVAL_125 = _EVAL_34 | _EVAL_261;
  assign _EVAL_151 = _EVAL_70 < plusarg_reader_out;
  assign _EVAL_48 = _EVAL_150 & _EVAL_119;
  assign _EVAL_241 = _EVAL_73 ? _EVAL_175 : 2'h0;
  assign _EVAL_206 = _EVAL_94 | _EVAL_4;
  assign _EVAL_24 = _EVAL_5 & _EVAL_178;
  assign _EVAL_146 = _EVAL_110 | _EVAL_4;
  assign _EVAL_183 = {_EVAL_88,_EVAL_99,_EVAL_125,_EVAL_226};
  assign _EVAL_268 = $signed(_EVAL_184) & -10'sh80;
  assign _EVAL_189 = _EVAL_217 - 1'h1;
  assign _EVAL_82 = _EVAL_5 & _EVAL_84;
  assign _EVAL_213 = _EVAL_167 | _EVAL_4;
  assign _EVAL_128 = _EVAL_1[0];
  assign _EVAL_255 = ~_EVAL_217;
  assign _EVAL_21 = ~_EVAL_72;
  assign _EVAL_198 = _EVAL_180 | _EVAL_187;
  assign _EVAL_244 = _EVAL_8 & _EVAL_161;
  assign _EVAL_103 = ~_EVAL_206;
  assign _EVAL_153 = _EVAL_199 | _EVAL_4;
  assign _EVAL_228 = _EVAL_104 | _EVAL_4;
  assign _EVAL_15 = _EVAL_8 & _EVAL_169;
  assign _EVAL_184 = {1'b0,$signed(_EVAL_131)};
  assign _EVAL_99 = _EVAL_157 | _EVAL_221;
  assign _EVAL_40 = $signed(_EVAL_67) == 10'sh0;
  assign _EVAL_235 = {1'b0,$signed(_EVAL_80)};
  assign _EVAL_67 = _EVAL_118;
  assign _EVAL_20 = _EVAL_112 & _EVAL_17;
  assign _EVAL_34 = _EVAL_97 | _EVAL_216;
  assign _EVAL_96 = ~_EVAL_147;
  assign _EVAL_110 = _EVAL_155 & _EVAL_195;
  assign _EVAL_66 = _EVAL_223 & _EVAL_18;
  assign _EVAL_84 = _EVAL_12 == 3'h5;
  assign _EVAL_111 = _EVAL_3 ^ 9'h60;
  assign _EVAL_22 = _EVAL_202;
  assign _EVAL_145 = _EVAL_5 & _EVAL_63;
  assign _EVAL_237 = _EVAL_30 >> _EVAL_10;
  assign _EVAL_53 = _EVAL != 3'h0;
  assign _EVAL_46 = _EVAL_12 == 3'h1;
  assign _EVAL_35 = _EVAL_5 & _EVAL_37;
  assign _EVAL_176 = {1'b0,$signed(_EVAL_3)};
  assign _EVAL_190 = _EVAL_185 | _EVAL_4;
  assign _EVAL_192 = $signed(_EVAL_194) & -10'shc;
  assign _EVAL_107 = _EVAL_11 >= 2'h2;
  assign _EVAL_130 = _EVAL_152 | _EVAL_4;
  assign _EVAL_114 = _EVAL_3 & _EVAL_238;
  assign _EVAL_243 = _EVAL_3[1];
  assign _EVAL_179 = |_EVAL_30;
  assign _EVAL_105 = _EVAL_2 == 3'h2;
  assign _EVAL_41 = _EVAL_258 | _EVAL_4;
  assign _EVAL_220 = _EVAL_28[0];
  assign _EVAL_230 = ~_EVAL_237;
  assign _EVAL_157 = _EVAL_97 | _EVAL_170;
  assign _EVAL_137 = _EVAL_107 | _EVAL_4;
  assign _EVAL_119 = ~_EVAL_144;
  assign _EVAL_210 = _EVAL_106 & _EVAL_267;
  assign _EVAL_122 = _EVAL_2 == 3'h3;
  assign _EVAL_64 = ~_EVAL_213;
  assign _EVAL_261 = _EVAL_25 & _EVAL_210;
  assign _EVAL_170 = _EVAL_257 & _EVAL_243;
  assign _EVAL_100 = ~_EVAL_162;
  assign _EVAL_113 = $signed(_EVAL_232) & -10'sh8;
  assign _EVAL_150 = _EVAL_7 & _EVAL_5;
  assign _EVAL_54 = _EVAL_16 ? _EVAL_31 : 2'h0;
  assign _EVAL_227 = _EVAL_168 | _EVAL_30;
  assign _EVAL_200 = _EVAL_2 == 3'h7;
  assign _EVAL_205 = _EVAL_208;
  assign _EVAL_38 = ~_EVAL_183;
  assign _EVAL_60 = ~_EVAL_228;
  assign _EVAL_168 = _EVAL_54[0];
  assign _EVAL_59 = _EVAL_12 == 3'h0;
  assign _EVAL_127 = ~_EVAL_41;
  assign _EVAL_253 = _EVAL == 3'h0;
  assign _EVAL_63 = ~_EVAL_119;
  assign _EVAL_77 = _EVAL_8 & _EVAL_105;
  assign _EVAL_72 = _EVAL_95 | _EVAL_4;
  assign _EVAL_112 = _EVAL_9 & _EVAL_8;
  assign _EVAL_258 = _EVAL_69 == 4'h0;
  assign _EVAL_101 = ~_EVAL_201;
  assign _EVAL_69 = _EVAL_13 & _EVAL_38;
  assign _EVAL_49 = _EVAL_251 | _EVAL_4;
  assign _EVAL_87 = _EVAL_268;
  assign _EVAL_158 = ~_EVAL_75;
  assign _EVAL_104 = _EVAL_1 == _EVAL_231;
  assign _EVAL_265 = _EVAL_144 - 1'h1;
  assign _EVAL_238 = {{7'd0}, _EVAL_158};
  assign _EVAL_147 = _EVAL_116 | _EVAL_4;
  assign _EVAL_141 = _EVAL_236 & _EVAL_199;
  assign _EVAL_52 = 2'h1 << _EVAL_128;
  assign _EVAL_250 = _EVAL == _EVAL_39;
  assign _EVAL_165 = _EVAL_5 & _EVAL_59;
  assign _EVAL_252 = _EVAL_2 == _EVAL_159;
  assign _EVAL_106 = ~_EVAL_243;
  assign _EVAL_207 = _EVAL_5 & _EVAL_262;
  assign _EVAL_121 = _EVAL_8 & _EVAL_254;
  assign _EVAL_102 = _EVAL_189[0];
  assign _EVAL_167 = _EVAL_3 == _EVAL_266;
  assign _EVAL_257 = _EVAL_55[1];
  assign _EVAL_155 = _EVAL_1 <= 2'h2;
  assign _EVAL_116 = _EVAL_0 == _EVAL_247;
  assign _EVAL_182 = _EVAL_12 <= 3'h6;
  assign _EVAL_174 = ~_EVAL_17;
  assign _EVAL_120 = ~_EVAL_267;
  assign _EVAL_126 = _EVAL_241[0];
  assign _EVAL_260 = _EVAL_156 | _EVAL_4;
  assign _EVAL_138 = _EVAL_141 | _EVAL_4;
  assign _EVAL_233 = _EVAL_248 | _EVAL_4;
  assign _EVAL_80 = _EVAL_3 ^ 9'h100;
  assign _EVAL_152 = _EVAL <= 3'h4;
  assign _EVAL_178 = _EVAL_12 == 3'h4;
  assign _EVAL_78 = ~_EVAL_259;
  assign _EVAL_160 = ~_EVAL_146;
  assign _EVAL_248 = _EVAL_227 >> _EVAL_0;
  assign _EVAL_140 = ~_EVAL_153;
  assign _EVAL_88 = _EVAL_157 | _EVAL_269;
  assign _EVAL_201 = _EVAL_253 | _EVAL_4;
  assign _EVAL_79 = ~_EVAL_137;
  assign _EVAL_131 = _EVAL_3 ^ 9'h80;
  assign _EVAL_76 = _EVAL_186 | _EVAL_4;
  assign _EVAL_194 = {1'b0,$signed(_EVAL_136)};
  assign _EVAL_216 = _EVAL_257 & _EVAL_106;
  assign _EVAL_132 = _EVAL_53 | _EVAL_4;
  assign _EVAL_32 = ~_EVAL_225;
  assign _EVAL_23 = $signed(_EVAL_87) == 10'sh0;
  assign _EVAL_256 = ~_EVAL_260;
  assign _EVAL_187 = $signed(_EVAL_117) == 10'sh0;
  assign _EVAL_177 = $signed(_EVAL_22) == 10'sh0;
  assign _EVAL_81 = _EVAL_250 | _EVAL_4;
  assign _EVAL_242 = ~_EVAL_123;
  assign _EVAL_175 = 2'h1 << _EVAL_0;
  assign _EVAL_91 = _EVAL_50 | _EVAL_4;
  assign _EVAL_93 = _EVAL_8 & _EVAL_174;
  assign _EVAL_55 = _EVAL_52 | 2'h1;
  assign _EVAL_161 = _EVAL_2 == 3'h4;
  assign _EVAL_196 = ~_EVAL_233;
  assign _EVAL_98 = ~_EVAL_4;
  assign _EVAL_26 = ~_EVAL_188;
  assign _EVAL_180 = _EVAL_177 | _EVAL_164;
  assign _EVAL_156 = ~_EVAL_0;
  always @(posedge _EVAL_14) begin
    if (_EVAL_4) begin
      _EVAL_30 <= 1'h0;
    end else begin
      _EVAL_30 <= _EVAL_66;
    end
    if (_EVAL_20) begin
      _EVAL_39 <= _EVAL;
    end
    if (_EVAL_4) begin
      _EVAL_70 <= 32'h0;
    end else if (_EVAL_197) begin
      _EVAL_70 <= 32'h0;
    end else begin
      _EVAL_70 <= _EVAL_129;
    end
    if (_EVAL_20) begin
      _EVAL_90 <= _EVAL_10;
    end
    if (_EVAL_4) begin
      _EVAL_92 <= 1'h0;
    end else if (_EVAL_112) begin
      if (_EVAL_108) begin
        _EVAL_92 <= 1'h0;
      end else begin
        _EVAL_92 <= _EVAL_263;
      end
    end
    if (_EVAL_4) begin
      _EVAL_109 <= 1'h0;
    end else if (_EVAL_112) begin
      if (_EVAL_17) begin
        _EVAL_109 <= 1'h0;
      end else begin
        _EVAL_109 <= _EVAL_220;
      end
    end
    if (_EVAL_48) begin
      _EVAL_135 <= _EVAL_12;
    end
    if (_EVAL_48) begin
      _EVAL_139 <= _EVAL_11;
    end
    if (_EVAL_4) begin
      _EVAL_144 <= 1'h0;
    end else if (_EVAL_150) begin
      if (_EVAL_119) begin
        _EVAL_144 <= 1'h0;
      end else begin
        _EVAL_144 <= _EVAL_68;
      end
    end
    if (_EVAL_20) begin
      _EVAL_159 <= _EVAL_2;
    end
    if (_EVAL_4) begin
      _EVAL_217 <= 1'h0;
    end else if (_EVAL_150) begin
      if (_EVAL_255) begin
        _EVAL_217 <= 1'h0;
      end else begin
        _EVAL_217 <= _EVAL_102;
      end
    end
    if (_EVAL_20) begin
      _EVAL_231 <= _EVAL_1;
    end
    if (_EVAL_48) begin
      _EVAL_247 <= _EVAL_0;
    end
    if (_EVAL_20) begin
      _EVAL_266 <= _EVAL_3;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a3121cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e83e3f69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c01120d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f1285e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3d05814)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6aaed6b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9e99a98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(523fa17b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fc6928c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d916047)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78991ada)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c4a7604)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e22b064a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3bdd7647)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(957b4780)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5701a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29df2a49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(faa08f1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(996e986)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3d1eca4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5499541)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff78af1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b5c9a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4f149dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c708182)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4fbe13d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(143d0d44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(466dbc06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f227a14b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_264) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bc0c1ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ded843e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f034a360)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_264) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b79a95c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd28019)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5a42e07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f4f18ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c927a38d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea09dde)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbdc1545)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf9fc3be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fd621b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(459e585b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dacd4855)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3179c9ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68489021)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15cbe659)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e02e2ed6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_5 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(241ad14f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c8c68be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd96bdf2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(613227a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ced1e0fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb7ea9df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3726a8d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f3bbe9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50ca9c6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89bc555d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(618c8de8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(270bce56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a60b5028)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(459e585b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(975bb474)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2f05e74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62055722)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c80e23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a39b7af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(daa674d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(218359c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d587d93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_256) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8c68e33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ac7eee1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7706982)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78cb089a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d25b2bc5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bac70c09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_30 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_39 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_70 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_90 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_92 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_109 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_135 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_139 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_144 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_159 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_217 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_231 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_247 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_266 = _RAND_13[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
