//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_46(
  input         _EVAL,
  output [2:0]  _EVAL_0,
  output        _EVAL_1,
  output [3:0]  _EVAL_2,
  output        _EVAL_3,
  output [11:0] _EVAL_4,
  input  [2:0]  _EVAL_5,
  output [4:0]  _EVAL_6,
  output        _EVAL_7,
  output [3:0]  _EVAL_8,
  input  [4:0]  _EVAL_9,
  input         _EVAL_10,
  output [2:0]  _EVAL_11,
  output [31:0] _EVAL_12,
  output [14:0] _EVAL_13,
  input  [4:0]  _EVAL_14,
  input  [1:0]  _EVAL_15,
  input  [2:0]  _EVAL_16,
  input  [31:0] _EVAL_17,
  output        _EVAL_18,
  input         _EVAL_19,
  input         _EVAL_20,
  output [31:0] _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23,
  input  [31:0] _EVAL_24,
  output        _EVAL_25,
  output        _EVAL_26,
  output [3:0]  _EVAL_27,
  output [1:0]  _EVAL_28,
  input         _EVAL_29,
  output [4:0]  _EVAL_30,
  output        _EVAL_31,
  input  [4:0]  _EVAL_32,
  input         _EVAL_33,
  output [2:0]  _EVAL_34,
  input         _EVAL_35,
  input  [1:0]  _EVAL_36,
  input         _EVAL_37,
  input         _EVAL_38,
  output [2:0]  _EVAL_39,
  output        _EVAL_40,
  input         _EVAL_41,
  output [25:0] _EVAL_42,
  output [3:0]  _EVAL_43,
  input         _EVAL_44,
  input         _EVAL_45,
  output [2:0]  _EVAL_46,
  output [2:0]  _EVAL_47,
  input         _EVAL_48,
  output [3:0]  _EVAL_49,
  output        _EVAL_50,
  output [2:0]  _EVAL_51,
  output        _EVAL_52,
  input  [31:0] _EVAL_53,
  output        _EVAL_54,
  output        _EVAL_55,
  output [2:0]  _EVAL_56,
  output [2:0]  _EVAL_57,
  output        _EVAL_58,
  output [2:0]  _EVAL_59,
  output        _EVAL_60,
  output        _EVAL_61,
  output [2:0]  _EVAL_62,
  output [3:0]  _EVAL_63,
  output [3:0]  _EVAL_64,
  input  [31:0] _EVAL_65,
  output        _EVAL_66,
  output        _EVAL_67,
  input         _EVAL_68,
  input  [2:0]  _EVAL_69,
  output        _EVAL_70,
  input         _EVAL_71,
  input  [4:0]  _EVAL_72,
  output [27:0] _EVAL_73,
  input  [31:0] _EVAL_74,
  input         _EVAL_75,
  input         _EVAL_76,
  input  [31:0] _EVAL_77,
  input  [2:0]  _EVAL_78,
  input  [2:0]  _EVAL_79,
  output        _EVAL_80,
  input  [4:0]  _EVAL_81,
  input         _EVAL_82,
  input  [2:0]  _EVAL_83,
  input         _EVAL_84,
  output        _EVAL_85,
  input         _EVAL_86,
  output [31:0] _EVAL_87,
  output        _EVAL_88,
  input  [2:0]  _EVAL_89,
  output        _EVAL_90,
  output [31:0] _EVAL_91,
  output [2:0]  _EVAL_92,
  output [4:0]  _EVAL_93,
  output [2:0]  _EVAL_94,
  output [2:0]  _EVAL_95,
  input  [2:0]  _EVAL_96,
  input         _EVAL_97,
  output        _EVAL_98,
  input  [31:0] _EVAL_99,
  input         _EVAL_100,
  output [2:0]  _EVAL_101,
  input  [2:0]  _EVAL_102,
  output        _EVAL_103,
  input  [4:0]  _EVAL_104,
  input  [31:0] _EVAL_105,
  input  [2:0]  _EVAL_106,
  input  [2:0]  _EVAL_107,
  output [3:0]  _EVAL_108,
  output        _EVAL_109,
  output [4:0]  _EVAL_110,
  input  [2:0]  _EVAL_111,
  input  [31:0] _EVAL_112,
  input  [3:0]  _EVAL_113,
  output [3:0]  _EVAL_114,
  output [2:0]  _EVAL_115,
  output [4:0]  _EVAL_116,
  output [2:0]  _EVAL_117,
  input  [2:0]  _EVAL_118,
  output [4:0]  _EVAL_119,
  output        _EVAL_120,
  output [2:0]  _EVAL_121,
  output        _EVAL_122,
  input  [2:0]  _EVAL_123,
  output [4:0]  _EVAL_124,
  input         _EVAL_125,
  output [13:0] _EVAL_126,
  input  [2:0]  _EVAL_127,
  input         _EVAL_128,
  output [29:0] _EVAL_129,
  input  [3:0]  _EVAL_130,
  input  [4:0]  _EVAL_131,
  input         _EVAL_132,
  output        _EVAL_133,
  output [2:0]  _EVAL_134,
  input  [3:0]  _EVAL_135,
  output [2:0]  _EVAL_136,
  output [4:0]  _EVAL_137,
  output [31:0] _EVAL_138,
  output [31:0] _EVAL_139,
  output        _EVAL_140,
  input  [4:0]  _EVAL_141,
  output [2:0]  _EVAL_142,
  input         _EVAL_143,
  output [31:0] _EVAL_144,
  output [31:0] _EVAL_145,
  input         _EVAL_146
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_147;
  wire [3:0] _EVAL_148;
  wire  _EVAL_149;
  wire [6:0] _EVAL_150;
  wire [6:0] _EVAL_151;
  wire [5:0] _EVAL_152;
  wire [32:0] _EVAL_153;
  wire [20:0] _EVAL_154;
  wire  _EVAL_155;
  wire [31:0] _EVAL_156;
  wire [32:0] _EVAL_157;
  wire [32:0] _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  reg [6:0] _EVAL_164;
  wire [6:0] _EVAL_165;
  wire [13:0] _EVAL_167;
  wire  _EVAL_168;
  wire [5:0] _EVAL_169;
  wire [3:0] _EVAL_170;
  wire [13:0] _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_174;
  wire [32:0] _EVAL_175;
  wire [2:0] _EVAL_176;
  wire  _EVAL_178;
  wire [3:0] _EVAL_179;
  wire [13:0] _EVAL_180;
  wire [31:0] _EVAL_181;
  wire  _EVAL_183;
  wire [4:0] _EVAL_184;
  wire [5:0] _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire [3:0] _EVAL_188;
  wire [4:0] _EVAL_189;
  reg  _EVAL_191;
  wire [2:0] _EVAL_192;
  wire [32:0] _EVAL_193;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_199;
  wire [5:0] _EVAL_200;
  wire [5:0] _EVAL_201;
  wire [22:0] _EVAL_202;
  wire [5:0] _EVAL_203;
  wire [32:0] _EVAL_204;
  wire [4:0] _EVAL_205;
  wire [13:0] _EVAL_206;
  wire [3:0] _EVAL_207;
  wire [20:0] _EVAL_208;
  wire [31:0] _EVAL_209;
  wire [6:0] _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire [4:0] _EVAL_215;
  wire [6:0] _EVAL_216;
  wire  _EVAL_218;
  wire  _EVAL_219;
  reg  _EVAL_221;
  wire [31:0] _EVAL_222;
  wire [3:0] _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire [3:0] _EVAL_226;
  wire  _EVAL_227;
  wire [3:0] _EVAL_228;
  wire  _EVAL_229;
  reg [5:0] _EVAL_231;
  wire [3:0] _EVAL_232;
  wire  _EVAL_233;
  wire [3:0] _EVAL_234;
  reg  _EVAL_236;
  wire [5:0] _EVAL_237;
  wire [3:0] _EVAL_238;
  wire [20:0] _EVAL_239;
  wire [31:0] _EVAL_240;
  wire [3:0] _EVAL_241;
  wire [13:0] _EVAL_242;
  wire [5:0] _EVAL_243;
  wire  _EVAL_244;
  wire [32:0] _EVAL_246;
  wire [3:0] _EVAL_247;
  wire [4:0] _EVAL_248;
  wire [31:0] _EVAL_249;
  wire [31:0] _EVAL_250;
  wire [4:0] _EVAL_251;
  wire [3:0] _EVAL_252;
  wire [32:0] _EVAL_253;
  wire [4:0] _EVAL_254;
  wire [2:0] _EVAL_257;
  wire  _EVAL_258;
  wire [31:0] _EVAL_259;
  wire [10:0] _EVAL_260;
  wire [32:0] _EVAL_261;
  wire  _EVAL_262;
  wire [3:0] _EVAL_263;
  wire [11:0] _EVAL_265;
  wire [1:0] _EVAL_266;
  wire [32:0] _EVAL_267;
  wire [2:0] _EVAL_268;
  wire [2:0] _EVAL_269;
  wire [3:0] _EVAL_270;
  wire [7:0] _EVAL_271;
  wire [2:0] _EVAL_274;
  wire  _EVAL_275;
  wire [2:0] _EVAL_276;
  wire [20:0] _EVAL_277;
  wire [5:0] _EVAL_278;
  wire  _EVAL_279;
  wire [1:0] _EVAL_280;
  wire [3:0] _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire [3:0] _EVAL_284;
  wire [31:0] _EVAL_285;
  wire [5:0] _EVAL_286;
  wire [3:0] _EVAL_287;
  wire [32:0] _EVAL_288;
  wire [3:0] _EVAL_289;
  wire [6:0] _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire [6:0] _EVAL_293;
  wire [5:0] _EVAL_294;
  wire [2:0] _EVAL_295;
  wire [5:0] _EVAL_296;
  wire  _EVAL_297;
  wire [8:0] _EVAL_298;
  wire [3:0] _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_302;
  wire  _EVAL_303;
  wire [3:0] _EVAL_304;
  wire [5:0] _EVAL_305;
  wire [32:0] _EVAL_306;
  wire [5:0] _EVAL_307;
  wire  _EVAL_308;
  wire [2:0] _EVAL_309;
  wire [32:0] _EVAL_310;
  wire [3:0] _EVAL_311;
  wire [3:0] _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_314;
  wire [5:0] _EVAL_316;
  wire [6:0] _EVAL_318;
  wire [6:0] _EVAL_319;
  wire [5:0] _EVAL_320;
  wire  _EVAL_321;
  wire  _EVAL_322;
  wire  _EVAL_323;
  wire [4:0] _EVAL_326;
  wire [31:0] _EVAL_327;
  wire [32:0] _EVAL_328;
  wire  _EVAL_330;
  wire  _EVAL_332;
  wire  _EVAL_333;
  wire  _EVAL_334;
  wire [31:0] _EVAL_335;
  wire  _EVAL_336;
  wire  _EVAL_337;
  wire  _EVAL_338;
  wire  _EVAL_339;
  wire [13:0] _EVAL_340;
  wire [6:0] _EVAL_341;
  wire  _EVAL_342;
  wire [32:0] _EVAL_343;
  wire [5:0] _EVAL_344;
  wire [32:0] _EVAL_345;
  wire [2:0] _EVAL_346;
  wire  _EVAL_347;
  wire  _EVAL_348;
  wire [3:0] _EVAL_351;
  wire  _EVAL_352;
  wire  _EVAL_353;
  wire [7:0] _EVAL_354;
  wire [9:0] _EVAL_355;
  wire [4:0] _EVAL_356;
  wire [2:0] _EVAL_357;
  wire  _EVAL_358;
  wire [4:0] _EVAL_359;
  wire [3:0] _EVAL_360;
  wire [3:0] _EVAL_361;
  wire  _EVAL_362;
  wire  _EVAL_364;
  wire [3:0] _EVAL_365;
  wire [31:0] _EVAL_366;
  wire  _EVAL_367;
  wire  _EVAL_368;
  wire [5:0] _EVAL_369;
  reg  _EVAL_370;
  wire [4:0] _EVAL_371;
  wire [32:0] _EVAL_372;
  wire [3:0] _EVAL_373;
  wire [2:0] _EVAL_374;
  wire  _EVAL_375;
  wire  _EVAL_377;
  wire  _EVAL_378;
  wire  _EVAL_379;
  wire [31:0] _EVAL_380;
  wire [32:0] _EVAL_381;
  wire [6:0] _EVAL_385;
  wire [31:0] _EVAL_386;
  wire [32:0] _EVAL_387;
  wire [5:0] _EVAL_388;
  wire [13:0] _EVAL_389;
  wire [31:0] _EVAL_390;
  wire [5:0] _EVAL_391;
  wire [7:0] _EVAL_392;
  reg  _EVAL_393;
  wire [32:0] _EVAL_394;
  wire [5:0] _EVAL_395;
  wire [3:0] _EVAL_396;
  wire [5:0] _EVAL_397;
  wire  _EVAL_398;
  wire [31:0] _EVAL_399;
  wire [3:0] _EVAL_400;
  wire [32:0] _EVAL_401;
  wire [5:0] _EVAL_402;
  wire  _EVAL_403;
  wire [12:0] _EVAL_404;
  wire [3:0] _EVAL_405;
  wire [13:0] _EVAL_407;
  wire [5:0] _EVAL_408;
  wire [3:0] _EVAL_409;
  wire [6:0] _EVAL_410;
  wire [13:0] _EVAL_411;
  wire [5:0] _EVAL_412;
  wire [32:0] _EVAL_414;
  wire  _EVAL_416;
  wire [5:0] _EVAL_418;
  wire  _EVAL_419;
  wire  _EVAL_421;
  wire [5:0] _EVAL_422;
  wire  _EVAL_424;
  wire  _EVAL_426;
  wire  _EVAL_427;
  wire  _EVAL_428;
  wire [6:0] _EVAL_429;
  wire [31:0] _EVAL_430;
  wire  _EVAL_431;
  wire [13:0] _EVAL_432;
  wire  _EVAL_433;
  wire [20:0] _EVAL_434;
  wire [3:0] _EVAL_435;
  wire  _EVAL_437;
  reg  _EVAL_438;
  wire [32:0] _EVAL_439;
  wire [5:0] _EVAL_440;
  wire [20:0] _EVAL_441;
  wire [31:0] _EVAL_442;
  wire [5:0] _EVAL_443;
  wire  _EVAL_444;
  wire [31:0] _EVAL_445;
  wire [4:0] _EVAL_446;
  wire [6:0] _EVAL_447;
  wire  _EVAL_448;
  wire  _EVAL_449;
  wire [3:0] _EVAL_450;
  wire [6:0] _EVAL_451;
  wire [32:0] _EVAL_452;
  wire  _EVAL_453;
  wire  _EVAL_454;
  wire [12:0] _EVAL_455;
  wire [3:0] _EVAL_456;
  reg  _EVAL_457;
  assign _EVAL_212 = _EVAL_199 & _EVAL_37;
  assign _EVAL_34 = _EVAL_83;
  assign _EVAL_185 = _EVAL_392[7:2];
  assign _EVAL_238 = _EVAL_361 | _EVAL_311;
  assign _EVAL_356 = _EVAL_446 | _EVAL_251;
  assign _EVAL_320 = {{5'd0}, _EVAL_282};
  assign _EVAL_181 = _EVAL_250 | _EVAL_335;
  assign _EVAL_430 = _EVAL_292 ? _EVAL_105 : 32'h0;
  assign _EVAL_398 = _EVAL_172 ? _EVAL_362 : _EVAL_236;
  assign _EVAL_2 = _EVAL_247 | _EVAL_289;
  assign _EVAL_80 = _EVAL_33 & _EVAL_419;
  assign _EVAL_379 = _EVAL_433 & _EVAL_75;
  assign _EVAL_294 = {{2'd0}, _EVAL_435};
  assign _EVAL_339 = _EVAL_172 ? _EVAL_227 : _EVAL_370;
  assign _EVAL_243 = ~_EVAL_391;
  assign _EVAL_25 = _EVAL_33 & _EVAL_375;
  assign _EVAL_27 = _EVAL_135;
  assign _EVAL_433 = _EVAL_429[6];
  assign _EVAL_222 = _EVAL_53 ^ 32'h2000000;
  assign _EVAL_374 = _EVAL_276 | _EVAL_346;
  assign _EVAL_26 = _EVAL_33 & _EVAL_183;
  assign _EVAL_40 = _EVAL_19 & _EVAL_449;
  assign _EVAL_196 = _EVAL_236 & _EVAL_29;
  assign _EVAL_375 = _EVAL_172 ? _EVAL_302 : _EVAL_393;
  assign _EVAL_229 = _EVAL_172 ? _EVAL_212 : _EVAL_191;
  assign _EVAL_435 = _EVAL_279 ? _EVAL_270 : 4'h0;
  assign _EVAL_395 = _EVAL_277[5:0];
  assign _EVAL_148 = _EVAL_159 ? _EVAL_241 : 4'h0;
  assign _EVAL_296 = _EVAL_239[5:0];
  assign _EVAL_57 = _EVAL_113[2:0];
  assign _EVAL_302 = _EVAL_429[0];
  assign _EVAL_386 = _EVAL_53 ^ 32'h2000;
  assign _EVAL_242 = {{4'd0}, _EVAL_355};
  assign _EVAL_51 = _EVAL_79;
  assign _EVAL_136 = _EVAL_113[2:0];
  assign _EVAL_122 = _EVAL_33 & _EVAL_336;
  assign _EVAL_115 = _EVAL_83;
  assign _EVAL_234 = _EVAL_292 ? _EVAL_130 : 4'h0;
  assign _EVAL_431 = _EVAL_332 | _EVAL_161;
  assign _EVAL_193 = $signed(_EVAL_343) & 33'shab004000;
  assign _EVAL_6 = _EVAL_14;
  assign _EVAL_199 = _EVAL_429[4];
  assign _EVAL_427 = _EVAL_225 | _EVAL_162;
  assign _EVAL_108 = _EVAL_113;
  assign _EVAL_318 = _EVAL_385 & _EVAL_447;
  assign _EVAL_354 = _EVAL_202[7:0];
  assign _EVAL_410 = ~_EVAL_164;
  assign _EVAL_340 = _EVAL_171 | _EVAL_407;
  assign _EVAL_95 = _EVAL_83;
  assign _EVAL_151 = _EVAL_271[6:0];
  assign _EVAL_157 = {1'b0,$signed(_EVAL_53)};
  assign _EVAL_439 = _EVAL_381;
  assign _EVAL_286 = _EVAL_316 | _EVAL_443;
  assign _EVAL_450 = {{1'd0}, _EVAL_127};
  assign _EVAL_434 = 21'h3f << _EVAL_405;
  assign _EVAL_405 = {{1'd0}, _EVAL_89};
  assign _EVAL_308 = $signed(_EVAL_158) == 33'sh0;
  assign _EVAL_178 = _EVAL_172 & _EVAL_33;
  assign _EVAL_293 = _EVAL_290 | _EVAL_341;
  assign _EVAL_192 = _EVAL_368 ? _EVAL_16 : 3'h0;
  assign _EVAL_60 = _EVAL_100;
  assign _EVAL_394 = _EVAL_253;
  assign _EVAL_145 = _EVAL_112;
  assign _EVAL_281 = _EVAL_339 ? _EVAL_287 : 4'h0;
  assign _EVAL_11 = _EVAL_113[2:0];
  assign _EVAL_327 = _EVAL_53 ^ 32'h20000000;
  assign _EVAL_455 = _EVAL_389[13:1];
  assign _EVAL_73 = _EVAL_53[27:0];
  assign _EVAL_101 = _EVAL_113[2:0];
  assign _EVAL_239 = 21'h3f << _EVAL_223;
  assign _EVAL_226 = _EVAL_243[5:2];
  assign _EVAL_207 = _EVAL_360 | _EVAL_232;
  assign _EVAL_451 = _EVAL_165 | _EVAL_151;
  assign _EVAL_276 = _EVAL_309 | _EVAL_269;
  assign _EVAL_309 = _EVAL_176 | _EVAL_268;
  assign _EVAL_345 = _EVAL_401;
  assign _EVAL_114 = _EVAL_135;
  assign _EVAL_278 = _EVAL_155 ? _EVAL_307 : 6'h0;
  assign _EVAL_47 = _EVAL_83;
  assign _EVAL_359 = _EVAL_353 ? _EVAL_104 : 5'h0;
  assign _EVAL_253 = $signed(_EVAL_387) & 33'shab006000;
  assign _EVAL_120 = _EVAL_19 & _EVAL_308;
  assign _EVAL_213 = _EVAL_172 ? _EVAL_168 : _EVAL_370;
  assign _EVAL_170 = _EVAL_333 ? _EVAL_188 : 4'h0;
  assign _EVAL_444 = _EVAL_197 | _EVAL_367;
  assign _EVAL_275 = $signed(_EVAL_306) == 33'sh0;
  assign _EVAL_208 = 21'h3f << _EVAL_409;
  assign _EVAL_316 = _EVAL_402 | _EVAL_201;
  assign _EVAL_169 = _EVAL_150[5:0];
  assign _EVAL_355 = _EVAL_180[13:4];
  assign _EVAL_88 = _EVAL_313 | _EVAL_347;
  assign _EVAL_422 = {{2'd0}, _EVAL_263};
  assign _EVAL_437 = _EVAL_292 & _EVAL;
  assign _EVAL_49 = _EVAL_135;
  assign _EVAL_426 = _EVAL_221 & _EVAL_45;
  assign _EVAL_119 = _EVAL_14;
  assign _EVAL_452 = $signed(_EVAL_157) & 33'shab006000;
  assign _EVAL_400 = _EVAL_368 ? _EVAL_373 : 4'h0;
  assign _EVAL_165 = _EVAL_429 & _EVAL_216;
  assign _EVAL_447 = _EVAL_340[6:0];
  assign _EVAL_176 = _EVAL_292 ? _EVAL_123 : 3'h0;
  assign _EVAL_367 = _EVAL_322 & _EVAL_20;
  assign _EVAL_210 = _EVAL_298[6:0];
  assign _EVAL_274 = _EVAL_257 | _EVAL_192;
  assign _EVAL_43 = _EVAL_135;
  assign _EVAL_224 = _EVAL_275 & _EVAL_10;
  assign _EVAL_133 = _EVAL_100;
  assign _EVAL_21 = _EVAL_112;
  assign _EVAL_416 = _EVAL_429[2];
  assign _EVAL_290 = _EVAL_451 | _EVAL_210;
  assign _EVAL_252 = _EVAL_227 ? _EVAL_148 : 4'h0;
  assign _EVAL_209 = _EVAL_53 ^ 32'h4000;
  assign _EVAL_402 = _EVAL_412 | _EVAL_422;
  assign _EVAL_172 = _EVAL_231 == 6'h0;
  assign _EVAL_91 = _EVAL_112;
  assign _EVAL_411 = {_EVAL_319,_EVAL_75,_EVAL_146,_EVAL_37,_EVAL_45,_EVAL_29,_EVAL_143,_EVAL_132};
  assign _EVAL_137 = _EVAL_14;
  assign _EVAL_259 = _EVAL_53 ^ 32'h1000000;
  assign _EVAL_216 = {_EVAL_75,_EVAL_146,_EVAL_37,_EVAL_45,_EVAL_29,_EVAL_143,_EVAL_132};
  assign _EVAL_257 = _EVAL_374 | _EVAL_295;
  assign _EVAL_396 = _EVAL_388[5:2];
  assign _EVAL_266 = _EVAL_292 ? _EVAL_36 : 2'h0;
  assign _EVAL_365 = _EVAL_233 ? _EVAL_351 : 4'h0;
  assign _EVAL_50 = _EVAL_19 & _EVAL_322;
  assign _EVAL_305 = ~_EVAL_418;
  assign _EVAL_389 = _EVAL_180 | _EVAL_242;
  assign _EVAL_456 = _EVAL_200[5:2];
  assign _EVAL_258 = _EVAL_300 | _EVAL_421;
  assign _EVAL_289 = _EVAL_211 ? _EVAL_450 : 4'h0;
  assign _EVAL_319 = _EVAL_216 & _EVAL_410;
  assign _EVAL_28 = _EVAL_266 | _EVAL_280;
  assign _EVAL_443 = {{2'd0}, _EVAL_299};
  assign _EVAL_110 = _EVAL_184 | _EVAL_205;
  assign _EVAL_251 = _EVAL_229 ? _EVAL_141 : 5'h0;
  assign _EVAL_303 = _EVAL_195 & _EVAL_41;
  assign _EVAL_442 = _EVAL_339 ? _EVAL_65 : 32'h0;
  assign _EVAL_233 = _EVAL_111[0];
  assign _EVAL_408 = _EVAL_441[5:0];
  assign _EVAL_61 = _EVAL_100;
  assign _EVAL_161 = _EVAL_378 & _EVAL_35;
  assign _EVAL_267 = {1'b0,$signed(_EVAL_390)};
  assign _EVAL_70 = _EVAL_437 | _EVAL_428;
  assign _EVAL_385 = _EVAL_340[13:7];
  assign _EVAL_150 = _EVAL_231 - _EVAL_320;
  assign _EVAL_328 = {1'b0,$signed(_EVAL_209)};
  assign _EVAL_381 = $signed(_EVAL_328) & 33'shab006000;
  assign _EVAL_432 = {{1'd0}, _EVAL_404};
  assign _EVAL_277 = 21'h3f << _EVAL_287;
  assign _EVAL_64 = _EVAL_135;
  assign _EVAL_92 = _EVAL_83;
  assign _EVAL_7 = _EVAL_19 & _EVAL_275;
  assign _EVAL_90 = _EVAL_33 & _EVAL_358;
  assign _EVAL_121 = _EVAL_79;
  assign _EVAL_156 = _EVAL_430 | _EVAL_442;
  assign _EVAL_87 = _EVAL_112;
  assign _EVAL_12 = _EVAL_112;
  assign _EVAL_269 = _EVAL_398 ? _EVAL_5 : 3'h0;
  assign _EVAL_63 = _EVAL_135;
  assign _EVAL_409 = {{1'd0}, _EVAL_107};
  assign _EVAL_429 = ~_EVAL_318;
  assign _EVAL_392 = ~_EVAL_354;
  assign _EVAL_387 = {1'b0,$signed(_EVAL_327)};
  assign _EVAL_346 = _EVAL_353 ? _EVAL_78 : 3'h0;
  assign _EVAL_202 = 23'hff << _EVAL_130;
  assign _EVAL_153 = _EVAL_414;
  assign _EVAL_323 = _EVAL_449 & _EVAL_86;
  assign _EVAL_138 = _EVAL_53;
  assign _EVAL_341 = _EVAL_260[6:0];
  assign _EVAL_219 = _EVAL_342 | _EVAL_426;
  assign _EVAL_344 = {{2'd0}, _EVAL_252};
  assign _EVAL_445 = _EVAL_156 | _EVAL_399;
  assign _EVAL_8 = _EVAL_135;
  assign _EVAL_246 = $signed(_EVAL_372) & 33'shab000000;
  assign _EVAL_454 = _EVAL_368 & _EVAL_71;
  assign _EVAL_397 = ~_EVAL_408;
  assign _EVAL_330 = _EVAL_5[0];
  assign _EVAL_241 = _EVAL_152[5:2];
  assign _EVAL_268 = _EVAL_339 ? _EVAL_96 : 3'h0;
  assign _EVAL_195 = $signed(_EVAL_394) == 33'sh0;
  assign _EVAL_321 = _EVAL_244 | _EVAL_45;
  assign _EVAL_3 = _EVAL_33 & _EVAL_213;
  assign _EVAL_271 = {_EVAL_165, 1'h0};
  assign _EVAL_13 = _EVAL_53[14:0];
  assign _EVAL_183 = _EVAL_172 ? _EVAL_453 : _EVAL_438;
  assign _EVAL_42 = _EVAL_53[25:0];
  assign _EVAL_361 = _EVAL_234 | _EVAL_281;
  assign _EVAL_168 = _EVAL_429[1];
  assign _EVAL_54 = _EVAL_160 | _EVAL_323;
  assign _EVAL_66 = _EVAL_84;
  assign _EVAL_18 = _EVAL_19 & _EVAL_378;
  assign _EVAL_184 = _EVAL_356 | _EVAL_215;
  assign _EVAL_404 = _EVAL_411[13:1];
  assign _EVAL_428 = _EVAL_368 & _EVAL_38;
  assign _EVAL_287 = {{1'd0}, _EVAL_102};
  assign _EVAL_283 = _EVAL_429[3];
  assign _EVAL_201 = {{2'd0}, _EVAL_170};
  assign _EVAL_117 = _EVAL_83;
  assign _EVAL_407 = {_EVAL_164, 7'h0};
  assign _EVAL_227 = _EVAL_168 & _EVAL_143;
  assign _EVAL_248 = _EVAL_254 | _EVAL_371;
  assign _EVAL_155 = _EVAL_302 & _EVAL_132;
  assign _EVAL_250 = _EVAL_240 | _EVAL_366;
  assign _EVAL_149 = _EVAL_457 & _EVAL_75;
  assign _EVAL_31 = _EVAL_23;
  assign _EVAL_62 = _EVAL_79;
  assign _EVAL_139 = _EVAL_112;
  assign _EVAL_335 = _EVAL_368 ? _EVAL_99 : 32'h0;
  assign _EVAL_215 = _EVAL_368 ? _EVAL_32 : 5'h0;
  assign _EVAL_357 = _EVAL_211 ? _EVAL_106 : 3'h0;
  assign _EVAL_265 = _EVAL_206[13:2];
  assign _EVAL_142 = _EVAL_113[2:0];
  assign _EVAL_163 = _EVAL_78[0];
  assign _EVAL_448 = _EVAL_172 ? _EVAL_283 : _EVAL_221;
  assign _EVAL_152 = ~_EVAL_395;
  assign _EVAL_225 = _EVAL_393 & _EVAL_132;
  assign _EVAL_94 = _EVAL_79;
  assign _EVAL_93 = _EVAL_14;
  assign _EVAL_1 = _EVAL_364 | _EVAL_454;
  assign _EVAL_228 = _EVAL_362 ? _EVAL_284 : 4'h0;
  assign _EVAL_158 = _EVAL_452;
  assign _EVAL_372 = {1'b0,$signed(_EVAL_285)};
  assign _EVAL_362 = _EVAL_416 & _EVAL_29;
  assign _EVAL_322 = _EVAL_147 | _EVAL_314;
  assign _EVAL_187 = _EVAL_16[0];
  assign _EVAL_126 = _EVAL_53[13:0];
  assign _EVAL_247 = _EVAL_207 | _EVAL_400;
  assign _EVAL_254 = _EVAL_292 ? _EVAL_131 : 5'h0;
  assign _EVAL_85 = _EVAL_19 & _EVAL_195;
  assign _EVAL_205 = _EVAL_211 ? _EVAL_81 : 5'h0;
  assign _EVAL_414 = $signed(_EVAL_267) & 33'shab004000;
  assign _EVAL_307 = _EVAL_174 ? _EVAL_185 : 6'h0;
  assign _EVAL_180 = _EVAL_206 | _EVAL_167;
  assign _EVAL_240 = _EVAL_445 | _EVAL_380;
  assign _EVAL_160 = _EVAL_444 | _EVAL_303;
  assign _EVAL_300 = _EVAL_219 | _EVAL_218;
  assign _EVAL_342 = _EVAL_427 | _EVAL_196;
  assign _EVAL_292 = _EVAL_172 ? _EVAL_155 : _EVAL_393;
  assign _EVAL_154 = 21'h3f << _EVAL_450;
  assign _EVAL_378 = $signed(_EVAL_345) == 33'sh0;
  assign _EVAL_306 = _EVAL_175;
  assign _EVAL_59 = _EVAL_79;
  assign _EVAL_314 = $signed(_EVAL_153) == 33'sh0;
  assign _EVAL_223 = {{1'd0}, _EVAL_118};
  assign _EVAL_403 = _EVAL_172 ? _EVAL_291 : _EVAL_262;
  assign _EVAL_377 = _EVAL_178 & _EVAL_297;
  assign _EVAL_261 = {1'b0,$signed(_EVAL_386)};
  assign _EVAL_304 = _EVAL_424 ? _EVAL_396 : 4'h0;
  assign _EVAL_312 = _EVAL_397[5:2];
  assign _EVAL_311 = _EVAL_398 ? _EVAL_409 : 4'h0;
  assign _EVAL_369 = {{2'd0}, _EVAL_228};
  assign _EVAL_204 = _EVAL_246;
  assign _EVAL_424 = _EVAL_106[0];
  assign _EVAL_147 = $signed(_EVAL_288) == 33'sh0;
  assign _EVAL_4 = _EVAL_53[11:0];
  assign _EVAL_284 = _EVAL_330 ? _EVAL_226 : 4'h0;
  assign _EVAL_171 = {{1'd0}, _EVAL_455};
  assign _EVAL_282 = _EVAL_33 & _EVAL_403;
  assign _EVAL_244 = _EVAL_334 | _EVAL_29;
  assign _EVAL_441 = 21'h3f << _EVAL_373;
  assign _EVAL_288 = _EVAL_193;
  assign _EVAL_188 = _EVAL_187 ? _EVAL_312 : 4'h0;
  assign _EVAL_52 = _EVAL_172 ? _EVAL_291 : _EVAL_262;
  assign _EVAL_140 = _EVAL_33 & _EVAL_448;
  assign _EVAL_421 = _EVAL_438 & _EVAL_146;
  assign _EVAL_67 = _EVAL_48;
  assign _EVAL_358 = _EVAL_172 ? _EVAL_416 : _EVAL_236;
  assign _EVAL_116 = _EVAL_14;
  assign _EVAL_159 = _EVAL_96[0];
  assign _EVAL_347 = _EVAL_368 & _EVAL_76;
  assign _EVAL_401 = $signed(_EVAL_310) & 33'shab000000;
  assign _EVAL_380 = _EVAL_353 ? _EVAL_24 : 32'h0;
  assign _EVAL_364 = _EVAL_292 & _EVAL_128;
  assign _EVAL_56 = _EVAL_83;
  assign _EVAL_162 = _EVAL_370 & _EVAL_143;
  assign _EVAL_129 = _EVAL_53[29:0];
  assign _EVAL_262 = _EVAL_258 | _EVAL_149;
  assign _EVAL_371 = _EVAL_339 ? _EVAL_72 : 5'h0;
  assign _EVAL_103 = _EVAL_44;
  assign _EVAL_453 = _EVAL_429[5];
  assign _EVAL_440 = _EVAL_203 | _EVAL_369;
  assign _EVAL_360 = _EVAL_238 | _EVAL_179;
  assign _EVAL_179 = _EVAL_353 ? _EVAL_223 : 4'h0;
  assign _EVAL_39 = _EVAL_113[2:0];
  assign _EVAL_30 = _EVAL_14;
  assign _EVAL_263 = _EVAL_212 ? _EVAL_365 : 4'h0;
  assign _EVAL_206 = _EVAL_411 | _EVAL_432;
  assign _EVAL_412 = _EVAL_440 | _EVAL_294;
  assign _EVAL_351 = _EVAL_305[5:2];
  assign _EVAL_343 = {1'b0,$signed(_EVAL_259)};
  assign _EVAL_295 = _EVAL_229 ? _EVAL_111 : 3'h0;
  assign _EVAL_186 = $signed(_EVAL_204) == 33'sh0;
  assign _EVAL_297 = |_EVAL_216;
  assign _EVAL_310 = {1'b0,$signed(_EVAL_222)};
  assign _EVAL_232 = _EVAL_229 ? _EVAL_405 : 4'h0;
  assign _EVAL_109 = _EVAL_100;
  assign _EVAL_298 = {_EVAL_451, 2'h0};
  assign _EVAL_368 = _EVAL_172 ? _EVAL_333 : _EVAL_438;
  assign _EVAL_332 = _EVAL_224 | _EVAL_348;
  assign _EVAL_203 = _EVAL_278 | _EVAL_344;
  assign _EVAL_390 = _EVAL_53 ^ 32'h80000000;
  assign _EVAL_449 = $signed(_EVAL_439) == 33'sh0;
  assign _EVAL_399 = _EVAL_398 ? _EVAL_77 : 32'h0;
  assign _EVAL_419 = _EVAL_172 ? _EVAL_199 : _EVAL_191;
  assign _EVAL_291 = _EVAL_337 | _EVAL_75;
  assign _EVAL_353 = _EVAL_172 ? _EVAL_279 : _EVAL_221;
  assign _EVAL_352 = _EVAL_308 & _EVAL_125;
  assign _EVAL_98 = _EVAL_100;
  assign _EVAL_167 = {{2'd0}, _EVAL_265};
  assign _EVAL_134 = _EVAL_79;
  assign _EVAL_285 = _EVAL_53 ^ 32'h8000000;
  assign _EVAL_174 = _EVAL_123[0];
  assign _EVAL_446 = _EVAL_189 | _EVAL_359;
  assign _EVAL_348 = _EVAL_186 & _EVAL_97;
  assign _EVAL_46 = _EVAL_79;
  assign _EVAL_144 = _EVAL_181 | _EVAL_249;
  assign _EVAL_211 = _EVAL_172 ? _EVAL_379 : _EVAL_457;
  assign _EVAL_391 = _EVAL_208[5:0];
  assign _EVAL_313 = _EVAL_292 & _EVAL_82;
  assign _EVAL_373 = {{1'd0}, _EVAL_69};
  assign _EVAL_336 = _EVAL_172 ? _EVAL_433 : _EVAL_457;
  assign _EVAL_299 = _EVAL_379 ? _EVAL_304 : 4'h0;
  assign _EVAL_197 = _EVAL_431 | _EVAL_352;
  assign _EVAL_334 = _EVAL_132 | _EVAL_143;
  assign _EVAL_175 = $signed(_EVAL_261) & 33'shab006000;
  assign _EVAL_326 = _EVAL_398 ? _EVAL_9 : 5'h0;
  assign _EVAL_249 = _EVAL_211 ? _EVAL_74 : 32'h0;
  assign _EVAL_338 = _EVAL_321 | _EVAL_37;
  assign _EVAL_388 = ~_EVAL_237;
  assign _EVAL_337 = _EVAL_338 | _EVAL_146;
  assign _EVAL_0 = _EVAL_274 | _EVAL_357;
  assign _EVAL_58 = _EVAL_100;
  assign _EVAL_55 = _EVAL_19 & _EVAL_186;
  assign _EVAL_218 = _EVAL_191 & _EVAL_37;
  assign _EVAL_279 = _EVAL_283 & _EVAL_45;
  assign _EVAL_280 = _EVAL_368 ? _EVAL_15 : 2'h0;
  assign _EVAL_237 = _EVAL_154[5:0];
  assign _EVAL_270 = _EVAL_163 ? _EVAL_456 : 4'h0;
  assign _EVAL_200 = ~_EVAL_296;
  assign _EVAL_124 = _EVAL_14;
  assign _EVAL_333 = _EVAL_453 & _EVAL_146;
  assign _EVAL_366 = _EVAL_229 ? _EVAL_17 : 32'h0;
  assign _EVAL_189 = _EVAL_248 | _EVAL_326;
  assign _EVAL_418 = _EVAL_434[5:0];
  assign _EVAL_260 = {_EVAL_290, 4'h0};
  always @(posedge _EVAL_22) begin
    if (_EVAL_68) begin
      _EVAL_164 <= 7'h7f;
    end else if (_EVAL_377) begin
      _EVAL_164 <= _EVAL_293;
    end
    if (_EVAL_68) begin
      _EVAL_191 <= 1'h0;
    end else if (_EVAL_172) begin
      _EVAL_191 <= _EVAL_212;
    end
    if (_EVAL_68) begin
      _EVAL_221 <= 1'h0;
    end else if (_EVAL_172) begin
      _EVAL_221 <= _EVAL_279;
    end
    if (_EVAL_68) begin
      _EVAL_231 <= 6'h0;
    end else if (_EVAL_178) begin
      _EVAL_231 <= _EVAL_286;
    end else begin
      _EVAL_231 <= _EVAL_169;
    end
    if (_EVAL_68) begin
      _EVAL_236 <= 1'h0;
    end else if (_EVAL_172) begin
      _EVAL_236 <= _EVAL_362;
    end
    if (_EVAL_68) begin
      _EVAL_370 <= 1'h0;
    end else if (_EVAL_172) begin
      _EVAL_370 <= _EVAL_227;
    end
    if (_EVAL_68) begin
      _EVAL_393 <= 1'h0;
    end else if (_EVAL_172) begin
      _EVAL_393 <= _EVAL_155;
    end
    if (_EVAL_68) begin
      _EVAL_438 <= 1'h0;
    end else if (_EVAL_172) begin
      _EVAL_438 <= _EVAL_333;
    end
    if (_EVAL_68) begin
      _EVAL_457 <= 1'h0;
    end else if (_EVAL_172) begin
      _EVAL_457 <= _EVAL_379;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_164 = _RAND_0[6:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_191 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_221 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_231 = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_236 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_370 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_393 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_438 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_457 = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
