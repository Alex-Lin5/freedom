//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
bind _EVAL_3 _EVAL_3_assert _EVAL_3_assert_0 (.*);
bind _EVAL_6 _EVAL_6_assert _EVAL_6_assert_0 (.*);
bind _EVAL_8 _EVAL_8_assert _EVAL_8_assert_0 (.*);
bind _EVAL_10 _EVAL_10_assert _EVAL_10_assert_0 (.*);
bind _EVAL_15 _EVAL_15_assert _EVAL_15_assert_0 (.*);
bind _EVAL_19 _EVAL_19_assert _EVAL_19_assert_0 (.*);
bind _EVAL_25 _EVAL_25_assert _EVAL_25_assert_0 (.*);
bind _EVAL_29 _EVAL_29_assert _EVAL_29_assert_0 (.*);
bind _EVAL_32 _EVAL_32_assert _EVAL_32_assert_0 (.*);
bind _EVAL_35 _EVAL_35_assert _EVAL_35_assert_0 (.*);
bind _EVAL_37 _EVAL_37_assert _EVAL_37_assert_0 (.*);
bind _EVAL_38 _EVAL_38_assert _EVAL_38_assert_0 (.*);
bind _EVAL_44 _EVAL_44_assert _EVAL_44_assert_0 (.*);
bind _EVAL_46 _EVAL_46_assert _EVAL_46_assert_0 (.*);
bind _EVAL_50 _EVAL_50_assert _EVAL_50_assert_0 (.*);
bind _EVAL_52 _EVAL_52_assert _EVAL_52_assert_0 (.*);
bind _EVAL_55 _EVAL_55_assert _EVAL_55_assert_0 (.*);
bind _EVAL_58 _EVAL_58_assert _EVAL_58_assert_0 (.*);
bind _EVAL_62 _EVAL_62_assert _EVAL_62_assert_0 (.*);
bind _EVAL_66 _EVAL_66_assert _EVAL_66_assert_0 (.*);
bind _EVAL_70 _EVAL_70_assert _EVAL_70_assert_0 (.*);
bind _EVAL_73 _EVAL_73_assert _EVAL_73_assert_0 (.*);
bind _EVAL_75 _EVAL_75_assert _EVAL_75_assert_0 (.*);
bind _EVAL_80 _EVAL_80_assert _EVAL_80_assert_0 (.*);
bind _EVAL_84 _EVAL_84_assert _EVAL_84_assert_0 (.*);
bind _EVAL_87 _EVAL_87_assert _EVAL_87_assert_0 (.*);
bind _EVAL_92 _EVAL_92_assert _EVAL_92_assert_0 (.*);
bind _EVAL_99 _EVAL_99_assert _EVAL_99_assert_0 (.*);
bind _EVAL_103 _EVAL_103_assert _EVAL_103_assert_0 (.*);
bind _EVAL_104 _EVAL_104_assert _EVAL_104_assert_0 (.*);
bind _EVAL_105 _EVAL_105_assert _EVAL_105_assert_0 (.*);
bind _EVAL_110 _EVAL_110_assert _EVAL_110_assert_0 (.*);
bind _EVAL_111 _EVAL_111_assert _EVAL_111_assert_0 (.*);
bind _EVAL_115 _EVAL_115_assert _EVAL_115_assert_0 (.*);
bind _EVAL_117 _EVAL_117_assert _EVAL_117_assert_0 (.*);
bind _EVAL_120 _EVAL_120_assert _EVAL_120_assert_0 (.*);
bind _EVAL_124 _EVAL_124_assert _EVAL_124_assert_0 (.*);
bind _EVAL_126 _EVAL_126_assert _EVAL_126_assert_0 (.*);
bind _EVAL_127 _EVAL_127_assert _EVAL_127_assert_0 (.*);
bind _EVAL_133 _EVAL_133_assert _EVAL_133_assert_0 (.*);
bind _EVAL_134 _EVAL_134_assert _EVAL_134_assert_0 (.*);
bind _EVAL_136 _EVAL_136_assert _EVAL_136_assert_0 (.*);
bind _EVAL_137 _EVAL_137_assert _EVAL_137_assert_0 (.*);
bind _EVAL_138 _EVAL_138_assert _EVAL_138_assert_0 (.*);
bind _EVAL_139 _EVAL_139_assert _EVAL_139_assert_0 (.*);
bind _EVAL_140 _EVAL_140_assert _EVAL_140_assert_0 (.*);
bind _EVAL_151 _EVAL_151_assert _EVAL_151_assert_0 (.*);
bind _EVAL_153 _EVAL_153_assert _EVAL_153_assert_0 (.*);
bind _EVAL_156 _EVAL_156_assert _EVAL_156_assert_0 (.*);
bind _EVAL_159 _EVAL_159_assert _EVAL_159_assert_0 (.*);
bind _EVAL_161 _EVAL_161_assert _EVAL_161_assert_0 (.*);
bind _EVAL_169 _EVAL_169_assert _EVAL_169_assert_0 (.*);
bind _EVAL_173 _EVAL_173_assert _EVAL_173_assert_0 (.*);
bind _EVAL_177 _EVAL_177_assert _EVAL_177_assert_0 (.*);
bind _EVAL_181 _EVAL_181_assert _EVAL_181_assert_0 (.*);
bind SiFive_TLTestIndicator SiFive_TLTestIndicator_assert SiFive_TLTestIndicator_assert_0 (.*);
bind _EVAL_197 _EVAL_197_assert _EVAL_197_assert_0 (.*);
bind _EVAL_198 _EVAL_198_assert _EVAL_198_assert_0 (.*);
bind _EVAL_199 _EVAL_199_assert _EVAL_199_assert_0 (.*);
bind _EVAL_200 _EVAL_200_assert _EVAL_200_assert_0 (.*);
bind _EVAL_201 _EVAL_201_assert _EVAL_201_assert_0 (.*);
bind _EVAL_203 _EVAL_203_assert _EVAL_203_assert_0 (.*);
bind _EVAL_204 _EVAL_204_assert _EVAL_204_assert_0 (.*);
bind SiFive_CoreIPSubsystem SiFive_CoreIPSubsystem_assert SiFive_CoreIPSubsystem_assert_0 (.*);