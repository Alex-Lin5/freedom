//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_24_assert(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input  [1:0]  _EVAL_3,
  input  [3:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input  [3:0]  _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  input  [31:0] _EVAL_14,
  input  [3:0]  _EVAL_15,
  input  [2:0]  _EVAL_16,
  input  [2:0]  _EVAL_17
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire [7:0] _EVAL_26;
  wire  _EVAL_27;
  wire [31:0] _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  reg [2:0] _EVAL_34;
  wire  _EVAL_35;
  wire [3:0] _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire [32:0] _EVAL_42;
  wire  _EVAL_43;
  wire [31:0] _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire [31:0] _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_61;
  wire  _EVAL_62;
  reg [3:0] _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire [5:0] _EVAL_67;
  wire [32:0] _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  reg  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  reg [5:0] _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire [32:0] _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_103;
  wire [6:0] _EVAL_104;
  wire [5:0] _EVAL_105;
  wire [32:0] _EVAL_106;
  wire [32:0] _EVAL_107;
  wire  _EVAL_108;
  wire [32:0] _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire [32:0] _EVAL_114;
  wire [31:0] _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire [6:0] _EVAL_121;
  wire  _EVAL_122;
  wire [6:0] _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire [3:0] _EVAL_130;
  wire  _EVAL_131;
  wire [1:0] _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire [1:0] _EVAL_136;
  wire [6:0] _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_141;
  wire [5:0] _EVAL_142;
  wire [1:0] _EVAL_144;
  wire [32:0] _EVAL_145;
  wire  _EVAL_146;
  wire [5:0] _EVAL_147;
  wire [32:0] _EVAL_148;
  wire  _EVAL_149;
  wire [32:0] _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire [3:0] _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  reg [3:0] _EVAL_160;
  wire  _EVAL_161;
  wire [3:0] _EVAL_162;
  wire [32:0] _EVAL_163;
  wire [32:0] _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire [22:0] _EVAL_170;
  wire [32:0] _EVAL_171;
  wire  _EVAL_172;
  wire [1:0] _EVAL_174;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire [31:0] _EVAL_180;
  wire  _EVAL_181;
  wire [32:0] _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  reg [5:0] _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire [7:0] _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_205;
  wire [32:0] _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire [31:0] _EVAL_210;
  reg  _EVAL_211;
  wire [31:0] _EVAL_212;
  wire  _EVAL_213;
  reg [1:0] _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  reg [31:0] _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire [32:0] _EVAL_245;
  wire  _EVAL_246;
  reg [5:0] _EVAL_247;
  reg [5:0] _EVAL_248;
  wire [32:0] _EVAL_249;
  wire  _EVAL_250;
  wire [5:0] _EVAL_251;
  wire [32:0] _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire [7:0] _EVAL_256;
  wire [5:0] _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire [32:0] _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  reg [31:0] _EVAL_263;
  wire [31:0] _EVAL_264;
  wire [32:0] _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  reg [2:0] _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire [32:0] _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire [32:0] _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire [31:0] _EVAL_292;
  wire  _EVAL_293;
  reg  _EVAL_294;
  wire  _EVAL_295;
  wire  _EVAL_296;
  wire  _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_302;
  reg [2:0] _EVAL_303;
  wire  _EVAL_304;
  wire [32:0] _EVAL_305;
  wire  _EVAL_306;
  wire [31:0] _EVAL_307;
  wire  _EVAL_308;
  wire  _EVAL_309;
  reg  _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire [7:0] _EVAL_314;
  wire  _EVAL_315;
  wire [32:0] _EVAL_316;
  wire  _EVAL_317;
  wire  _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_320;
  wire  _EVAL_321;
  wire  _EVAL_322;
  wire  _EVAL_323;
  wire [22:0] _EVAL_324;
  wire  _EVAL_325;
  wire  _EVAL_326;
  wire  _EVAL_327;
  wire  _EVAL_328;
  wire  _EVAL_329;
  wire [1:0] _EVAL_330;
  wire  _EVAL_331;
  wire  _EVAL_332;
  wire [32:0] _EVAL_333;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_30 = ~_EVAL_184;
  assign _EVAL_194 = _EVAL_16 == 3'h4;
  assign _EVAL_206 = _EVAL_148;
  assign _EVAL_135 = ~_EVAL_185;
  assign _EVAL_157 = _EVAL_215 & _EVAL_183;
  assign _EVAL_296 = _EVAL_301 & _EVAL_128;
  assign _EVAL_37 = _EVAL_241 < plusarg_reader_out;
  assign _EVAL_151 = {1'b0,$signed(_EVAL_28)};
  assign _EVAL_315 = _EVAL_97 | _EVAL_13;
  assign _EVAL_321 = _EVAL_14 == _EVAL_263;
  assign _EVAL_256 = ~_EVAL_26;
  assign _EVAL_212 = _EVAL_14 ^ 32'h40000000;
  assign _EVAL_35 = ~_EVAL_13;
  assign _EVAL_25 = ~_EVAL_81;
  assign _EVAL_301 = _EVAL_4 <= 4'hb;
  assign _EVAL_107 = {1'b0,$signed(_EVAL_44)};
  assign _EVAL_217 = _EVAL_215 & _EVAL_283;
  assign _EVAL_323 = _EVAL_73 | _EVAL_318;
  assign _EVAL_285 = ~_EVAL_2;
  assign _EVAL_131 = _EVAL_144[1];
  assign _EVAL_118 = ~_EVAL_279;
  assign _EVAL_196 = _EVAL_16 == 3'h6;
  assign _EVAL_245 = _EVAL_114;
  assign _EVAL_81 = _EVAL_285 | _EVAL_13;
  assign _EVAL_290 = _EVAL_327 & _EVAL_56;
  assign _EVAL_320 = _EVAL_4 == _EVAL_160;
  assign _EVAL_279 = _EVAL_261 | _EVAL_13;
  assign _EVAL_250 = _EVAL_132[0];
  assign _EVAL_120 = _EVAL_11 & _EVAL_226;
  assign _EVAL_293 = _EVAL_12 != 3'h0;
  assign _EVAL_210 = _EVAL_14 ^ 32'h2000000;
  assign _EVAL_275 = _EVAL_16 == 3'h3;
  assign _EVAL_98 = ~_EVAL_133;
  assign _EVAL_80 = _EVAL_11 & _EVAL_196;
  assign _EVAL_209 = _EVAL_103 | _EVAL_13;
  assign _EVAL_69 = _EVAL_17[0];
  assign _EVAL_286 = $signed(_EVAL_206) == 33'sh0;
  assign _EVAL_44 = _EVAL_14 ^ 32'h20000000;
  assign _EVAL_170 = 23'hff << _EVAL_4;
  assign _EVAL_58 = _EVAL_90 | _EVAL_13;
  assign _EVAL_189 = _EVAL_88 | _EVAL_13;
  assign _EVAL_40 = _EVAL_82 | _EVAL_149;
  assign _EVAL_197 = ~_EVAL_76;
  assign _EVAL_306 = _EVAL_300 & _EVAL_237;
  assign _EVAL_156 = _EVAL_219 | _EVAL_13;
  assign _EVAL_238 = _EVAL_65 | _EVAL_13;
  assign _EVAL_96 = _EVAL_79 | _EVAL_141;
  assign _EVAL_89 = _EVAL_6 & _EVAL_122;
  assign _EVAL_326 = _EVAL_205 | _EVAL_13;
  assign _EVAL_137 = _EVAL_247 - 6'h1;
  assign _EVAL_187 = ~_EVAL_189;
  assign _EVAL_65 = _EVAL_155 == 4'h0;
  assign _EVAL_314 = ~_EVAL_201;
  assign _EVAL_234 = _EVAL_167 | _EVAL_13;
  assign _EVAL_292 = _EVAL_14 & _EVAL_307;
  assign _EVAL_289 = ~_EVAL_242;
  assign _EVAL_31 = _EVAL_14[1];
  assign _EVAL_24 = |_EVAL_318;
  assign _EVAL_110 = _EVAL_6 & _EVAL_45;
  assign _EVAL_277 = ~_EVAL_322;
  assign _EVAL_332 = _EVAL_3 != 2'h2;
  assign _EVAL_32 = _EVAL_292 == 32'h0;
  assign _EVAL_145 = {1'b0,$signed(_EVAL_14)};
  assign _EVAL_225 = _EVAL_6 & _EVAL_124;
  assign _EVAL_152 = ~_EVAL_45;
  assign _EVAL_207 = ~_EVAL_83;
  assign _EVAL_226 = _EVAL_16 == 3'h0;
  assign _EVAL_242 = _EVAL_158 | _EVAL_13;
  assign _EVAL_49 = ~_EVAL_116;
  assign _EVAL_48 = _EVAL_66 | _EVAL_79;
  assign _EVAL_258 = _EVAL_297 | _EVAL_13;
  assign _EVAL_95 = {1'b0,$signed(_EVAL_212)};
  assign _EVAL_243 = ~_EVAL_315;
  assign _EVAL_121 = _EVAL_248 - 6'h1;
  assign _EVAL_153 = _EVAL_77 | _EVAL_13;
  assign _EVAL_174 = _EVAL_217 ? _EVAL_330 : 2'h0;
  assign _EVAL_284 = _EVAL_230 | _EVAL_199;
  assign _EVAL_23 = _EVAL_6 & _EVAL_138;
  assign _EVAL_28 = _EVAL_14 ^ 32'h80000000;
  assign _EVAL_240 = _EVAL_202 & _EVAL_152;
  assign _EVAL_72 = ~_EVAL_8;
  assign _EVAL_123 = _EVAL_193 - 6'h1;
  assign _EVAL_192 = ~_EVAL_302;
  assign _EVAL_36 = {_EVAL_223,_EVAL_284,_EVAL_40,_EVAL_312};
  assign _EVAL_159 = _EVAL_11 & _EVAL_288;
  assign _EVAL_195 = _EVAL_207 | _EVAL_13;
  assign _EVAL_218 = _EVAL_332 | _EVAL_13;
  assign _EVAL_75 = ~_EVAL_58;
  assign _EVAL_283 = _EVAL_84 == 6'h0;
  assign _EVAL_146 = _EVAL_318 != _EVAL_250;
  assign _EVAL_176 = _EVAL_59 | _EVAL_13;
  assign _EVAL_78 = _EVAL_327 & _EVAL_96;
  assign _EVAL_287 = $signed(_EVAL_95) & -33'sh2000;
  assign _EVAL_90 = _EVAL_12 == 3'h0;
  assign _EVAL_291 = ~_EVAL_86;
  assign _EVAL_255 = ~_EVAL_218;
  assign _EVAL_268 = _EVAL_72 | _EVAL_13;
  assign _EVAL_312 = _EVAL_82 | _EVAL_306;
  assign _EVAL_273 = ~_EVAL_99;
  assign _EVAL_318 = _EVAL_174[0];
  assign _EVAL_139 = ~_EVAL_20;
  assign _EVAL_29 = ~_EVAL_209;
  assign _EVAL_213 = _EVAL_93 | _EVAL_13;
  assign _EVAL_198 = _EVAL_216 | _EVAL_13;
  assign _EVAL_172 = _EVAL_16 == 3'h5;
  assign _EVAL_122 = _EVAL_17 == 3'h5;
  assign _EVAL_104 = _EVAL_84 - 6'h1;
  assign _EVAL_93 = _EVAL_4 >= 4'h2;
  assign _EVAL_181 = _EVAL_11 & _EVAL_275;
  assign _EVAL_64 = _EVAL_295 | _EVAL_13;
  assign _EVAL_39 = ~_EVAL_268;
  assign _EVAL_45 = _EVAL_17 == 3'h6;
  assign _EVAL_74 = |_EVAL_73;
  assign _EVAL_288 = _EVAL_16 == 3'h2;
  assign _EVAL_253 = _EVAL_11 & _EVAL_172;
  assign _EVAL_191 = ~_EVAL_24;
  assign _EVAL_325 = _EVAL_193 == 6'h0;
  assign _EVAL_164 = _EVAL_265;
  assign _EVAL_219 = _EVAL_12 <= 3'h2;
  assign _EVAL_166 = ~_EVAL_154;
  assign _EVAL_322 = _EVAL_190 | _EVAL_13;
  assign _EVAL_87 = _EVAL_31 & _EVAL_291;
  assign _EVAL_161 = _EVAL_188 | _EVAL_227;
  assign _EVAL_86 = _EVAL_14[0];
  assign _EVAL_105 = _EVAL_123[5:0];
  assign _EVAL_79 = $signed(_EVAL_106) == 33'sh0;
  assign _EVAL_91 = _EVAL_12 <= 3'h4;
  assign _EVAL_83 = _EVAL_73 >> _EVAL_0;
  assign _EVAL_55 = _EVAL_14 ^ 32'h1800000;
  assign _EVAL_57 = ~_EVAL_308;
  assign _EVAL_106 = _EVAL_274;
  assign _EVAL_265 = $signed(_EVAL_260) & -33'sh1000;
  assign _EVAL_330 = 2'h1 << _EVAL_0;
  assign _EVAL_85 = ~_EVAL_153;
  assign _EVAL_249 = _EVAL_252;
  assign _EVAL_130 = ~_EVAL_15;
  assign _EVAL_51 = _EVAL_4 <= 4'h8;
  assign _EVAL_165 = _EVAL_52 | _EVAL_13;
  assign _EVAL_99 = _EVAL_254 | _EVAL_13;
  assign _EVAL_108 = _EVAL_3 == _EVAL_214;
  assign _EVAL_27 = _EVAL_17 == 3'h1;
  assign _EVAL_333 = _EVAL_171;
  assign _EVAL_267 = ~_EVAL_331;
  assign _EVAL_269 = _EVAL_6 & _EVAL_27;
  assign _EVAL_304 = _EVAL_3 == 2'h0;
  assign _EVAL_20 = _EVAL_91 | _EVAL_13;
  assign _EVAL_112 = _EVAL_2 == _EVAL_294;
  assign _EVAL_260 = {1'b0,$signed(_EVAL_264)};
  assign _EVAL_228 = _EVAL_3 <= 2'h2;
  assign _EVAL_266 = _EVAL_177 | _EVAL_13;
  assign _EVAL_246 = ~_EVAL_31;
  assign _EVAL_38 = _EVAL_16[2];
  assign _EVAL_216 = _EVAL_262 | _EVAL_37;
  assign _EVAL_42 = {1'b0,$signed(_EVAL_55)};
  assign _EVAL_300 = _EVAL_144[0];
  assign _EVAL_274 = $signed(_EVAL_107) & -33'sh2000;
  assign _EVAL_222 = _EVAL_327 & _EVAL_161;
  assign _EVAL_88 = _EVAL_5 == _EVAL_211;
  assign _EVAL_59 = _EVAL_12 <= 3'h3;
  assign _EVAL_271 = _EVAL_108 | _EVAL_13;
  assign _EVAL_126 = ~_EVAL_234;
  assign _EVAL_155 = _EVAL_15 & _EVAL_162;
  assign _EVAL_313 = _EVAL_300 & _EVAL_281;
  assign _EVAL_257 = _EVAL_137[5:0];
  assign _EVAL_134 = ~_EVAL_282;
  assign _EVAL_149 = _EVAL_300 & _EVAL_129;
  assign _EVAL_70 = ~_EVAL_176;
  assign _EVAL_254 = _EVAL_54 | _EVAL_78;
  assign _EVAL_125 = ~_EVAL_1;
  assign _EVAL_208 = ~_EVAL_229;
  assign _EVAL_68 = $signed(_EVAL_109) & -33'sh400000;
  assign _EVAL_46 = _EVAL & _EVAL_6;
  assign _EVAL_163 = _EVAL_241 + 32'h1;
  assign _EVAL_328 = _EVAL_128 | _EVAL_13;
  assign _EVAL_272 = ~_EVAL_113;
  assign _EVAL_33 = _EVAL_317 | _EVAL_286;
  assign _EVAL_200 = ~_EVAL_326;
  assign _EVAL_169 = ~_EVAL_74;
  assign _EVAL_144 = _EVAL_136 | 2'h1;
  assign _EVAL_168 = $signed(_EVAL_333) == 33'sh0;
  assign _EVAL_113 = _EVAL_296 | _EVAL_13;
  assign _EVAL_282 = _EVAL_112 | _EVAL_13;
  assign _EVAL_186 = ~_EVAL_213;
  assign _EVAL_19 = _EVAL_11 & _EVAL_21;
  assign _EVAL_264 = _EVAL_14 ^ 32'h3000;
  assign _EVAL_205 = _EVAL_296 & _EVAL_309;
  assign _EVAL_47 = _EVAL_11 & _EVAL_329;
  assign _EVAL_231 = _EVAL_11 & _EVAL_194;
  assign _EVAL_239 = ~_EVAL_238;
  assign _EVAL_299 = plusarg_reader_out == 32'h0;
  assign _EVAL_236 = ~_EVAL_198;
  assign _EVAL_220 = $signed(_EVAL_249) == 33'sh0;
  assign _EVAL_94 = ~_EVAL_266;
  assign _EVAL_100 = _EVAL_215 | _EVAL_46;
  assign _EVAL_307 = {{24'd0}, _EVAL_314};
  assign _EVAL_66 = _EVAL_33 | _EVAL_179;
  assign _EVAL_251 = _EVAL_256[7:2];
  assign _EVAL_202 = _EVAL_46 & _EVAL_325;
  assign _EVAL_133 = _EVAL_244 | _EVAL_13;
  assign _EVAL_232 = ~_EVAL_38;
  assign _EVAL_117 = ~_EVAL_165;
  assign _EVAL_308 = _EVAL_178 | _EVAL_13;
  assign _EVAL_82 = _EVAL_93 | _EVAL_61;
  assign _EVAL_199 = _EVAL_300 & _EVAL_87;
  assign _EVAL_54 = _EVAL_51 & _EVAL_259;
  assign _EVAL_309 = _EVAL_54 | _EVAL_222;
  assign _EVAL_237 = _EVAL_246 & _EVAL_291;
  assign _EVAL_71 = _EVAL_131 & _EVAL_31;
  assign _EVAL_158 = _EVAL_17 == _EVAL_303;
  assign _EVAL_230 = _EVAL_93 | _EVAL_71;
  assign _EVAL_138 = _EVAL_17 == 3'h0;
  assign _EVAL_331 = _EVAL_125 | _EVAL_13;
  assign _EVAL_41 = ~_EVAL_156;
  assign _EVAL_136 = 2'h1 << _EVAL_276;
  assign _EVAL_182 = _EVAL_287;
  assign _EVAL_223 = _EVAL_230 | _EVAL_313;
  assign _EVAL_111 = ~_EVAL_328;
  assign _EVAL_76 = _EVAL_309 | _EVAL_13;
  assign _EVAL_167 = _EVAL_0 == _EVAL_311;
  assign _EVAL_227 = $signed(_EVAL_245) == 33'sh0;
  assign _EVAL_114 = $signed(_EVAL_151) & -33'sh4000;
  assign _EVAL_142 = _EVAL_104[5:0];
  assign _EVAL_261 = _EVAL_17 <= 3'h6;
  assign _EVAL_235 = _EVAL_46 & _EVAL_229;
  assign _EVAL_116 = _EVAL_278 | _EVAL_13;
  assign _EVAL_278 = _EVAL_12 <= 3'h1;
  assign _EVAL_132 = _EVAL_240 ? 2'h1 : 2'h0;
  assign _EVAL_185 = _EVAL_320 | _EVAL_13;
  assign _EVAL_22 = ~_EVAL_271;
  assign _EVAL_18 = ~_EVAL_101;
  assign _EVAL_148 = $signed(_EVAL_305) & -33'sh10000;
  assign _EVAL_179 = $signed(_EVAL_316) == 33'sh0;
  assign _EVAL_50 = _EVAL_323 & _EVAL_319;
  assign _EVAL_21 = ~_EVAL_183;
  assign _EVAL_43 = _EVAL_11 & _EVAL_203;
  assign _EVAL_183 = _EVAL_248 == 6'h0;
  assign _EVAL_324 = 23'hff << _EVAL_10;
  assign _EVAL_244 = _EVAL_318 | _EVAL_73;
  assign _EVAL_62 = _EVAL_293 | _EVAL_13;
  assign _EVAL_67 = _EVAL_121[5:0];
  assign _EVAL_203 = _EVAL_16 == 3'h1;
  assign _EVAL_101 = _EVAL_32 | _EVAL_13;
  assign _EVAL_188 = _EVAL_48 | _EVAL_141;
  assign _EVAL_147 = _EVAL_314[7:2];
  assign _EVAL_252 = $signed(_EVAL_145) & -33'sh5000;
  assign _EVAL_129 = _EVAL_246 & _EVAL_86;
  assign _EVAL_92 = ~_EVAL_62;
  assign _EVAL_177 = _EVAL_54 | _EVAL_290;
  assign _EVAL_316 = _EVAL_68;
  assign _EVAL_127 = _EVAL_6 & _EVAL_208;
  assign _EVAL_190 = _EVAL_12 == _EVAL_34;
  assign _EVAL_128 = ~_EVAL_0;
  assign _EVAL_297 = _EVAL_146 | _EVAL_191;
  assign _EVAL_97 = _EVAL_16 == _EVAL_270;
  assign _EVAL_229 = _EVAL_247 == 6'h0;
  assign _EVAL_276 = _EVAL_4[0];
  assign _EVAL_26 = _EVAL_324[7:0];
  assign _EVAL_141 = $signed(_EVAL_182) == 33'sh0;
  assign _EVAL_295 = _EVAL_10 >= 4'h2;
  assign _EVAL_302 = _EVAL_321 | _EVAL_13;
  assign _EVAL_259 = $signed(_EVAL_164) == 33'sh0;
  assign _EVAL_52 = _EVAL_15 == _EVAL_36;
  assign _EVAL_180 = _EVAL_14 ^ 32'hc000000;
  assign _EVAL_53 = _EVAL_6 & _EVAL_298;
  assign _EVAL_162 = ~_EVAL_36;
  assign _EVAL_305 = {1'b0,$signed(_EVAL_210)};
  assign _EVAL_327 = _EVAL_4 <= 4'h6;
  assign _EVAL_178 = _EVAL_285 | _EVAL_1;
  assign _EVAL_109 = {1'b0,$signed(_EVAL_180)};
  assign _EVAL_124 = _EVAL_17 == 3'h4;
  assign _EVAL_233 = ~_EVAL_195;
  assign _EVAL_329 = _EVAL_16 == 3'h7;
  assign _EVAL_184 = _EVAL_304 | _EVAL_13;
  assign _EVAL_154 = _EVAL_228 | _EVAL_13;
  assign _EVAL_115 = _EVAL_163[31:0];
  assign _EVAL_56 = _EVAL_66 | _EVAL_227;
  assign _EVAL_262 = _EVAL_169 | _EVAL_299;
  assign _EVAL_119 = ~_EVAL_258;
  assign _EVAL_224 = ~_EVAL_64;
  assign _EVAL_103 = _EVAL_130 == 4'h0;
  assign _EVAL_319 = ~_EVAL_250;
  assign _EVAL_171 = $signed(_EVAL_42) & -33'sh4000;
  assign _EVAL_215 = _EVAL_9 & _EVAL_11;
  assign _EVAL_61 = _EVAL_131 & _EVAL_246;
  assign _EVAL_201 = _EVAL_170[7:0];
  assign _EVAL_77 = _EVAL_10 == _EVAL_63;
  assign _EVAL_281 = _EVAL_31 & _EVAL_86;
  assign _EVAL_317 = _EVAL_220 | _EVAL_168;
  assign _EVAL_298 = _EVAL_17 == 3'h2;
  always @(posedge _EVAL_7) begin
    if (_EVAL_157) begin
      _EVAL_34 <= _EVAL_12;
    end
    if (_EVAL_235) begin
      _EVAL_63 <= _EVAL_10;
    end
    if (_EVAL_13) begin
      _EVAL_73 <= 1'h0;
    end else begin
      _EVAL_73 <= _EVAL_50;
    end
    if (_EVAL_13) begin
      _EVAL_84 <= 6'h0;
    end else if (_EVAL_215) begin
      if (_EVAL_283) begin
        if (_EVAL_232) begin
          _EVAL_84 <= _EVAL_147;
        end else begin
          _EVAL_84 <= 6'h0;
        end
      end else begin
        _EVAL_84 <= _EVAL_142;
      end
    end
    if (_EVAL_157) begin
      _EVAL_160 <= _EVAL_4;
    end
    if (_EVAL_13) begin
      _EVAL_193 <= 6'h0;
    end else if (_EVAL_46) begin
      if (_EVAL_325) begin
        if (_EVAL_69) begin
          _EVAL_193 <= _EVAL_251;
        end else begin
          _EVAL_193 <= 6'h0;
        end
      end else begin
        _EVAL_193 <= _EVAL_105;
      end
    end
    if (_EVAL_235) begin
      _EVAL_211 <= _EVAL_5;
    end
    if (_EVAL_235) begin
      _EVAL_214 <= _EVAL_3;
    end
    if (_EVAL_13) begin
      _EVAL_241 <= 32'h0;
    end else if (_EVAL_100) begin
      _EVAL_241 <= 32'h0;
    end else begin
      _EVAL_241 <= _EVAL_115;
    end
    if (_EVAL_13) begin
      _EVAL_247 <= 6'h0;
    end else if (_EVAL_46) begin
      if (_EVAL_229) begin
        if (_EVAL_69) begin
          _EVAL_247 <= _EVAL_251;
        end else begin
          _EVAL_247 <= 6'h0;
        end
      end else begin
        _EVAL_247 <= _EVAL_257;
      end
    end
    if (_EVAL_13) begin
      _EVAL_248 <= 6'h0;
    end else if (_EVAL_215) begin
      if (_EVAL_183) begin
        if (_EVAL_232) begin
          _EVAL_248 <= _EVAL_147;
        end else begin
          _EVAL_248 <= 6'h0;
        end
      end else begin
        _EVAL_248 <= _EVAL_67;
      end
    end
    if (_EVAL_157) begin
      _EVAL_263 <= _EVAL_14;
    end
    if (_EVAL_157) begin
      _EVAL_270 <= _EVAL_16;
    end
    if (_EVAL_235) begin
      _EVAL_294 <= _EVAL_2;
    end
    if (_EVAL_235) begin
      _EVAL_303 <= _EVAL_17;
    end
    if (_EVAL_157) begin
      _EVAL_311 <= _EVAL_0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_289) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb38aa00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b5a0f06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(714464bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9c30e49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_255) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32149494)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86a75040)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_49) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf44e2df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(721b0970)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_25) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98f444df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f79dbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6810a024)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0a80fcd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da99645f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa3beb73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ade29e72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6502ece9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_197) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8973ef18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f368e7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_289) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb76526e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f8ea883)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f988994)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d1d23a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0ebd37e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a78c67d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4cb1a4fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e92c8cf5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_273) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a5d5282)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18a4b0d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(712742a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_49) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d4d545c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9321952)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(196965b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74da1502)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5834e05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_139) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64315535)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12e60ff6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d50bdc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3f9c70e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f8ea0a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(594c31d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5335eefc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e374b611)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_224) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_255) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7305a98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b91eb5ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_255) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8cbae113)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28913d3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_239) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49a99fb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(672cca0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_272) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5adf5346)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4da24bb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(911ea7b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(803bfea5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_186) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c320226)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52a1b109)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_272) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72d98bda)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63502a1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37f92993)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e902205f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45354780)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d1b0c5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d34d115)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_273) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9eb8386d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6380074d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e96966)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2b62259)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_231 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c183b117)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(881ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19144137)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_224) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7e0dd1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb8610b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf631267)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_139) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d367052)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35aac0da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd37a181)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(678c28a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_255) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97fa6dbe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_239) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c748d81a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_25) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13ddc35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(faf1d23b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4da24bb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_253 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65fc6ac3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(311194)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(232e637a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab341295)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_186) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(631227c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e1399af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc5dd0f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_34 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_63 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_73 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_84 = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_160 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_193 = _RAND_5[5:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_211 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_214 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_241 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_247 = _RAND_9[5:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_248 = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_263 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_270 = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_294 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_303 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_311 = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
