//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_130(
  input         _EVAL,
  output        _EVAL_0,
  output [31:0] _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input  [3:0]  _EVAL_4,
  input         _EVAL_5,
  input  [31:0] _EVAL_6,
  output [4:0]  _EVAL_7,
  input  [4:0]  _EVAL_8,
  input  [31:0] _EVAL_9,
  input         _EVAL_10,
  output        _EVAL_11
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [95:0] _RAND_6;
  reg [63:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_12;
  wire [3:0] _EVAL_13;
  wire [15:0] _EVAL_14;
  wire [15:0] _EVAL_15;
  wire [3:0] _EVAL_16;
  wire [7:0] _EVAL_17;
  wire  _EVAL_18;
  wire [3:0] _EVAL_19;
  wire [3:0] _EVAL_20;
  wire [15:0] _EVAL_21;
  wire [7:0] _EVAL_22;
  reg  _EVAL_23;
  wire [3:0] _EVAL_24;
  wire  _EVAL_26;
  wire [1:0] _EVAL_27;
  wire [3:0] _EVAL_28;
  wire [31:0] _EVAL_30;
  wire [1:0] _EVAL_31;
  wire  _EVAL_32;
  wire [64:0] _EVAL_33;
  wire [31:0] _EVAL_34;
  wire [2:0] _EVAL_35;
  wire [1:0] _EVAL_36;
  wire [4:0] _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire [31:0] _EVAL_41;
  wire [32:0] _EVAL_42;
  wire [2:0] _EVAL_43;
  wire [3:0] _EVAL_44;
  wire [1:0] _EVAL_45;
  wire [3:0] _EVAL_46;
  wire [3:0] _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire [1:0] _EVAL_50;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire [1:0] _EVAL_54;
  wire  _EVAL_55;
  wire [1:0] _EVAL_56;
  wire [3:0] _EVAL_57;
  wire [1:0] _EVAL_58;
  wire  _EVAL_59;
  wire [1:0] _EVAL_60;
  reg  _EVAL_61;
  wire [15:0] _EVAL_62;
  wire [3:0] _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire [1:0] _EVAL_72;
  wire [2:0] _EVAL_73;
  wire [2:0] _EVAL_74;
  wire [2:0] _EVAL_75;
  wire [2:0] _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire [65:0] _EVAL_79;
  wire [7:0] _EVAL_80;
  wire [3:0] _EVAL_81;
  wire [2:0] _EVAL_82;
  reg  _EVAL_83;
  wire  _EVAL_84;
  wire [15:0] _EVAL_85;
  wire [5:0] _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire [2:0] _EVAL_91;
  reg [2:0] _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire [3:0] _EVAL_97;
  wire [15:0] _EVAL_98;
  wire  _EVAL_99;
  wire [15:0] _EVAL_100;
  wire  _EVAL_101;
  wire [7:0] _EVAL_102;
  wire  _EVAL_103;
  wire [1:0] _EVAL_104;
  wire [1:0] _EVAL_105;
  wire [2:0] _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire [2:0] _EVAL_111;
  reg [5:0] _EVAL_112;
  wire [2:0] _EVAL_113;
  wire  _EVAL_114;
  wire [31:0] _EVAL_116;
  wire [1:0] _EVAL_117;
  wire  _EVAL_118;
  wire [2:0] _EVAL_119;
  wire [1:0] _EVAL_120;
  wire [1:0] _EVAL_121;
  wire [1:0] _EVAL_122;
  wire [3:0] _EVAL_123;
  wire  _EVAL_124;
  wire [33:0] _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire [2:0] _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire [1:0] _EVAL_134;
  wire [3:0] _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire [1:0] _EVAL_138;
  wire [7:0] _EVAL_139;
  wire [5:0] _EVAL_140;
  wire [1:0] _EVAL_141;
  wire  _EVAL_142;
  wire [32:0] _EVAL_143;
  wire [4:0] _EVAL_144;
  wire [62:0] _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire [1:0] _EVAL_148;
  wire  _EVAL_149;
  wire [3:0] _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire [3:0] _EVAL_154;
  wire [1:0] _EVAL_155;
  wire [1:0] _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire [62:0] _EVAL_159;
  wire [15:0] _EVAL_160;
  wire [1:0] _EVAL_161;
  wire [3:0] _EVAL_162;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire [1:0] _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire [7:0] _EVAL_171;
  wire  _EVAL_173;
  wire [3:0] _EVAL_174;
  wire [6:0] _EVAL_175;
  wire [1:0] _EVAL_176;
  wire  _EVAL_177;
  wire [3:0] _EVAL_178;
  wire [1:0] _EVAL_179;
  wire  _EVAL_180;
  reg [4:0] _EVAL_181;
  wire [1:0] _EVAL_182;
  wire [1:0] _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire [1:0] _EVAL_186;
  reg [65:0] _EVAL_187;
  wire  _EVAL_188;
  wire [31:0] _EVAL_189;
  wire [1:0] _EVAL_190;
  wire [3:0] _EVAL_191;
  wire  _EVAL_192;
  wire [3:0] _EVAL_193;
  wire  _EVAL_194;
  wire [4:0] _EVAL_195;
  wire  _EVAL_196;
  wire [32:0] _EVAL_197;
  wire [1:0] _EVAL_198;
  wire [3:0] _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire [1:0] _EVAL_202;
  wire  _EVAL_203;
  wire [2:0] _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire [1:0] _EVAL_208;
  wire [7:0] _EVAL_209;
  wire [1:0] _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  reg [32:0] _EVAL_216;
  wire [32:0] _EVAL_217;
  wire [2:0] _EVAL_218;
  wire  _EVAL_219;
  wire [1:0] _EVAL_220;
  wire [7:0] _EVAL_221;
  wire [31:0] _EVAL_222;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire [1:0] _EVAL_226;
  wire  _EVAL_227;
  wire [31:0] _EVAL_228;
  wire [1:0] _EVAL_229;
  wire [3:0] _EVAL_230;
  wire  _EVAL_231;
  wire [2:0] _EVAL_232;
  wire  _EVAL_233;
  wire [31:0] _EVAL_234;
  wire [1:0] _EVAL_235;
  wire [1:0] _EVAL_236;
  wire [4:0] _EVAL_237;
  wire  _EVAL_238;
  wire [1:0] _EVAL_239;
  wire  _EVAL_240;
  wire [15:0] _EVAL_241;
  wire  _EVAL_242;
  wire [64:0] _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire [31:0] _EVAL_248;
  wire [15:0] _EVAL_249;
  wire  _EVAL_250;
  assign _EVAL_242 = _EVAL_44[2];
  assign _EVAL_221 = _EVAL_14[7:0];
  assign _EVAL_65 = _EVAL_24[1];
  assign _EVAL_162 = {_EVAL_196,_EVAL_119};
  assign _EVAL_174 = _EVAL_171[7:4];
  assign _EVAL_200 = _EVAL_238 & _EVAL_136;
  assign _EVAL_106 = {_EVAL_124,_EVAL_60};
  assign _EVAL_212 = _EVAL_131 | _EVAL_18;
  assign _EVAL_155 = _EVAL_225 ? 2'h2 : {{1'd0}, _EVAL_101};
  assign _EVAL_136 = ~_EVAL_96;
  assign _EVAL_45 = _EVAL_59 ? 2'h3 : _EVAL_31;
  assign _EVAL_239 = _EVAL_149 ? _EVAL_182 : _EVAL_202;
  assign _EVAL_75 = _EVAL_89 ? 3'h7 : _EVAL_43;
  assign _EVAL_111 = _EVAL_23 ? 3'h5 : 3'h7;
  assign _EVAL_72 = _EVAL_70 ? 2'h3 : _EVAL_229;
  assign _EVAL_117 = _EVAL_170 ? 2'h2 : {{1'd0}, _EVAL_180};
  assign _EVAL_31 = _EVAL_12 ? 2'h2 : {{1'd0}, _EVAL_65};
  assign _EVAL_49 = _EVAL_150 == 4'h2;
  assign _EVAL_43 = _EVAL_247 ? 3'h3 : _EVAL_92;
  assign _EVAL_58 = _EVAL_184 ? 2'h2 : {{1'd0}, _EVAL_94};
  assign _EVAL_154 = _EVAL_171[3:0];
  assign _EVAL_33 = _EVAL_52 ? {{2'd0}, _EVAL_145} : _EVAL_243;
  assign _EVAL_13 = _EVAL_80[7:4];
  assign _EVAL_203 = _EVAL_63[3];
  assign _EVAL_81 = _EVAL_139[3:0];
  assign _EVAL_217 = 32'h0 - _EVAL_248;
  assign _EVAL_249 = _EVAL_6[15:0];
  assign _EVAL_87 = _EVAL_97[1];
  assign _EVAL_237 = {_EVAL_38,_EVAL_123};
  assign _EVAL_234 = _EVAL_217[31:0];
  assign _EVAL_77 = _EVAL_132 | _EVAL_2;
  assign _EVAL_93 = _EVAL_20[1];
  assign _EVAL_148 = _EVAL_26 ? 2'h3 : _EVAL_236;
  assign _EVAL_219 = _EVAL_135[2];
  assign _EVAL_107 = _EVAL_178[3];
  assign _EVAL_137 = |_EVAL_174;
  assign _EVAL_14 = _EVAL_189[31:16];
  assign _EVAL_101 = _EVAL_174[1];
  assign _EVAL_73 = {_EVAL_137,_EVAL_120};
  assign _EVAL_165 = _EVAL_230[2];
  assign _EVAL_171 = _EVAL_15[15:8];
  assign _EVAL_11 = _EVAL_213 | _EVAL_153;
  assign _EVAL_128 = _EVAL_191[3];
  assign _EVAL_135 = _EVAL_22[3:0];
  assign _EVAL_35 = _EVAL_194 ? _EVAL_204 : _EVAL_113;
  assign _EVAL_18 = _EVAL_108 & _EVAL_95;
  assign _EVAL_152 = _EVAL_0 & _EVAL_3;
  assign _EVAL_213 = _EVAL_92 == 3'h6;
  assign _EVAL_193 = _EVAL_67 ? _EVAL_28 : _EVAL_16;
  assign _EVAL_123 = _EVAL_38 ? _EVAL_19 : _EVAL_162;
  assign _EVAL_243 = {_EVAL_41,_EVAL_189,_EVAL_207};
  assign _EVAL_129 = |_EVAL_44;
  assign _EVAL_98 = _EVAL_34[31:16];
  assign _EVAL_85 = _EVAL_9[31:16];
  assign _EVAL_227 = _EVAL_97[2];
  assign _EVAL_124 = |_EVAL_230;
  assign _EVAL_63 = _EVAL_221[3:0];
  assign _EVAL_202 = _EVAL_39 ? 2'h3 : _EVAL_117;
  assign _EVAL_102 = _EVAL_100[7:0];
  assign _EVAL_250 = _EVAL_191[2];
  assign _EVAL_57 = _EVAL_4 & 4'h1;
  assign _EVAL_156 = _EVAL_242 ? 2'h2 : {{1'd0}, _EVAL_177};
  assign _EVAL_30 = _EVAL_187[64:33];
  assign _EVAL_210 = _EVAL_64 ? 2'h2 : {{1'd0}, _EVAL_173};
  assign _EVAL_195 = {_EVAL_67,_EVAL_193};
  assign _EVAL_99 = _EVAL_20[2];
  assign _EVAL_147 = _EVAL_6[31];
  assign _EVAL_204 = {_EVAL_185,_EVAL_141};
  assign _EVAL_211 = |_EVAL_209;
  assign _EVAL_47 = _EVAL_17[3:0];
  assign _EVAL_178 = _EVAL_209[7:4];
  assign _EVAL_225 = _EVAL_174[2];
  assign _EVAL_205 = |_EVAL_17;
  assign _EVAL_142 = _EVAL_143[32];
  assign _EVAL_127 = _EVAL_230[1];
  assign _EVAL_82 = _EVAL_211 ? _EVAL_76 : _EVAL_91;
  assign _EVAL_131 = _EVAL_108 & _EVAL_147;
  assign _EVAL_44 = _EVAL_102[7:4];
  assign _EVAL_52 = _EVAL_200 & _EVAL_231;
  assign _EVAL_79 = _EVAL_78 ? {{34'd0}, _EVAL_234} : _EVAL_187;
  assign _EVAL_173 = _EVAL_46[1];
  assign _EVAL_12 = _EVAL_24[2];
  assign _EVAL_88 = _EVAL_13[3];
  assign _EVAL_71 = _EVAL_46[3];
  assign _EVAL_160 = _EVAL_248[31:16];
  assign _EVAL_42 = {_EVAL_18,_EVAL_85,_EVAL_241};
  assign _EVAL_130 = _EVAL_205 ? _EVAL_106 : _EVAL_218;
  assign _EVAL_0 = _EVAL_92 == 3'h0;
  assign _EVAL_146 = _EVAL_112 == 6'h20;
  assign _EVAL_145 = _EVAL_159 << _EVAL_144;
  assign _EVAL_240 = _EVAL_131 != _EVAL_18;
  assign _EVAL_138 = _EVAL_158 ? 2'h3 : _EVAL_156;
  assign _EVAL_197 = _EVAL_187[64:32];
  assign _EVAL_89 = _EVAL_92 == 3'h5;
  assign _EVAL_114 = _EVAL_154[2];
  assign _EVAL_16 = {_EVAL_205,_EVAL_130};
  assign _EVAL_238 = _EVAL_112 == 6'h0;
  assign _EVAL_182 = _EVAL_107 ? 2'h3 : _EVAL_54;
  assign _EVAL_170 = _EVAL_199[2];
  assign _EVAL_100 = _EVAL_34[15:0];
  assign _EVAL_80 = _EVAL_14[15:8];
  assign _EVAL_59 = _EVAL_24[3];
  assign _EVAL_20 = _EVAL_80[3:0];
  assign _EVAL_229 = _EVAL_227 ? 2'h2 : {{1'd0}, _EVAL_87};
  assign _EVAL_231 = _EVAL_144 >= 5'h1;
  assign _EVAL_235 = _EVAL_133 ? 2'h3 : _EVAL_122;
  assign _EVAL_90 = _EVAL_96 & _EVAL_188;
  assign _EVAL_122 = _EVAL_164 ? 2'h2 : {{1'd0}, _EVAL_233};
  assign _EVAL_19 = {_EVAL_194,_EVAL_35};
  assign _EVAL_158 = _EVAL_44[3];
  assign _EVAL_95 = _EVAL_9[31];
  assign _EVAL_48 = _EVAL_230[3];
  assign _EVAL_246 = |_EVAL_97;
  assign _EVAL_168 = _EVAL_219 ? 2'h2 : {{1'd0}, _EVAL_32};
  assign _EVAL_153 = _EVAL_92 == 3'h7;
  assign _EVAL_206 = |_EVAL_24;
  assign _EVAL_15 = _EVAL_189[15:0];
  assign _EVAL_104 = _EVAL_48 ? 2'h3 : _EVAL_183;
  assign _EVAL_177 = _EVAL_44[1];
  assign _EVAL_53 = _EVAL_178[2];
  assign _EVAL_133 = _EVAL_47[3];
  assign _EVAL_125 = _EVAL_197 - _EVAL_216;
  assign _EVAL_248 = _EVAL_83 ? _EVAL_30 : _EVAL_189;
  assign _EVAL_236 = _EVAL_114 ? 2'h2 : {{1'd0}, _EVAL_84};
  assign _EVAL_55 = _EVAL_92 == 3'h3;
  assign _EVAL_67 = |_EVAL_98;
  assign _EVAL_209 = _EVAL_98[15:8];
  assign _EVAL_199 = _EVAL_209[3:0];
  assign _EVAL_118 = _EVAL_81[3];
  assign _EVAL_84 = _EVAL_154[1];
  assign _EVAL_39 = _EVAL_199[3];
  assign _EVAL_149 = |_EVAL_178;
  assign _EVAL_22 = _EVAL_15[7:0];
  assign _EVAL_186 = _EVAL_71 ? 2'h3 : _EVAL_210;
  assign _EVAL_68 = _EVAL_89 ? 1'h0 : _EVAL_83;
  assign _EVAL_180 = _EVAL_199[1];
  assign _EVAL_103 = _EVAL_81[2];
  assign _EVAL_179 = _EVAL_103 ? 2'h2 : {{1'd0}, _EVAL_245};
  assign _EVAL_198 = _EVAL_203 ? 2'h3 : _EVAL_50;
  assign _EVAL_60 = _EVAL_124 ? _EVAL_104 : _EVAL_235;
  assign _EVAL_36 = _EVAL_129 ? _EVAL_138 : _EVAL_134;
  assign _EVAL_17 = _EVAL_100[15:8];
  assign _EVAL_76 = {_EVAL_149,_EVAL_239};
  assign _EVAL_21 = _EVAL_248[15:0];
  assign _EVAL_166 = _EVAL_63[2];
  assign _EVAL_119 = _EVAL_196 ? _EVAL_73 : _EVAL_232;
  assign _EVAL_26 = _EVAL_154[3];
  assign _EVAL_28 = {_EVAL_211,_EVAL_82};
  assign _EVAL_224 = _EVAL_20[3];
  assign _EVAL_54 = _EVAL_53 ? 2'h2 : {{1'd0}, _EVAL_151};
  assign _EVAL_37 = _EVAL_140[4:0];
  assign _EVAL_144 = ~_EVAL_37;
  assign _EVAL_245 = _EVAL_81[1];
  assign _EVAL_139 = _EVAL_98[7:0];
  assign _EVAL_140 = _EVAL_237 - _EVAL_195;
  assign _EVAL_32 = _EVAL_135[1];
  assign _EVAL_247 = _EVAL_92 == 3'h1;
  assign _EVAL_220 = _EVAL_224 ? 2'h3 : _EVAL_208;
  assign _EVAL_46 = _EVAL_221[7:4];
  assign _EVAL_189 = _EVAL_187[31:0];
  assign _EVAL_56 = _EVAL_118 ? 2'h3 : _EVAL_179;
  assign _EVAL_134 = _EVAL_128 ? 2'h3 : _EVAL_161;
  assign _EVAL_244 = |_EVAL_46;
  assign _EVAL_241 = _EVAL_9[15:0];
  assign _EVAL_176 = _EVAL_169 ? 2'h3 : _EVAL_168;
  assign _EVAL_34 = _EVAL_216[31:0];
  assign _EVAL_201 = _EVAL_216[31];
  assign _EVAL_232 = {_EVAL_246,_EVAL_190};
  assign _EVAL_207 = ~_EVAL_142;
  assign _EVAL_175 = _EVAL_112 + 6'h1;
  assign _EVAL_62 = _EVAL_6[31:16];
  assign _EVAL_159 = {{31'd0}, _EVAL_189};
  assign _EVAL_38 = |_EVAL_14;
  assign _EVAL_157 = _EVAL_191[1];
  assign _EVAL_64 = _EVAL_46[2];
  assign _EVAL_78 = _EVAL_187[31];
  assign _EVAL_185 = |_EVAL_13;
  assign _EVAL_143 = _EVAL_125[32:0];
  assign _EVAL_70 = _EVAL_97[3];
  assign _EVAL_120 = _EVAL_137 ? _EVAL_226 : _EVAL_148;
  assign _EVAL_41 = _EVAL_142 ? _EVAL_116 : _EVAL_222;
  assign _EVAL_121 = _EVAL_88 ? 2'h3 : _EVAL_58;
  assign _EVAL_222 = _EVAL_143[31:0];
  assign _EVAL_141 = _EVAL_185 ? _EVAL_121 : _EVAL_220;
  assign _EVAL_188 = ~_EVAL_61;
  assign _EVAL_94 = _EVAL_13[1];
  assign _EVAL_24 = _EVAL_139[7:4];
  assign _EVAL_161 = _EVAL_250 ? 2'h2 : {{1'd0}, _EVAL_157};
  assign _EVAL_116 = _EVAL_187[63:32];
  assign _EVAL_50 = _EVAL_166 ? 2'h2 : {{1'd0}, _EVAL_126};
  assign _EVAL_74 = _EVAL_146 ? _EVAL_111 : _EVAL_75;
  assign _EVAL_151 = _EVAL_178[1];
  assign _EVAL_150 = _EVAL_4 & 4'h2;
  assign _EVAL_97 = _EVAL_22[7:4];
  assign _EVAL_192 = _EVAL_174[3];
  assign _EVAL_108 = _EVAL_57 == 4'h0;
  assign _EVAL_105 = _EVAL_206 ? _EVAL_45 : _EVAL_56;
  assign _EVAL_228 = {_EVAL_62,_EVAL_249};
  assign _EVAL_96 = _EVAL_238 & _EVAL_207;
  assign _EVAL_126 = _EVAL_63[1];
  assign _EVAL_194 = |_EVAL_80;
  assign _EVAL_208 = _EVAL_99 ? 2'h2 : {{1'd0}, _EVAL_93};
  assign _EVAL_218 = {_EVAL_129,_EVAL_36};
  assign _EVAL_191 = _EVAL_102[3:0];
  assign _EVAL_196 = |_EVAL_171;
  assign _EVAL_169 = _EVAL_135[3];
  assign _EVAL_164 = _EVAL_47[2];
  assign _EVAL_91 = {_EVAL_206,_EVAL_105};
  assign _EVAL_7 = _EVAL_181;
  assign _EVAL_86 = _EVAL_175[5:0];
  assign _EVAL_230 = _EVAL_17[7:4];
  assign _EVAL_1 = {_EVAL_160,_EVAL_21};
  assign _EVAL_190 = _EVAL_246 ? _EVAL_72 : _EVAL_176;
  assign _EVAL_113 = {_EVAL_244,_EVAL_27};
  assign _EVAL_233 = _EVAL_47[1];
  assign _EVAL_226 = _EVAL_192 ? 2'h3 : _EVAL_155;
  assign _EVAL_132 = _EVAL_10 & _EVAL_11;
  assign _EVAL_183 = _EVAL_165 ? 2'h2 : {{1'd0}, _EVAL_127};
  assign _EVAL_184 = _EVAL_13[2];
  assign _EVAL_27 = _EVAL_244 ? _EVAL_186 : _EVAL_198;
  always @(posedge _EVAL) begin
    if (_EVAL_152) begin
      if (_EVAL_49) begin
        _EVAL_23 <= _EVAL_131;
      end else begin
        _EVAL_23 <= _EVAL_240;
      end
    end else if (_EVAL_55) begin
      if (_EVAL_90) begin
        _EVAL_23 <= 1'h0;
      end
    end
    if (_EVAL_152) begin
      _EVAL_61 <= _EVAL_49;
    end
    if (_EVAL_152) begin
      _EVAL_83 <= 1'h0;
    end else if (_EVAL_55) begin
      if (_EVAL_146) begin
        _EVAL_83 <= _EVAL_61;
      end else begin
        _EVAL_83 <= _EVAL_68;
      end
    end else begin
      _EVAL_83 <= _EVAL_68;
    end
    if (_EVAL_5) begin
      _EVAL_92 <= 3'h0;
    end else if (_EVAL_152) begin
      if (_EVAL_212) begin
        _EVAL_92 <= 3'h1;
      end else begin
        _EVAL_92 <= 3'h3;
      end
    end else if (_EVAL_77) begin
      _EVAL_92 <= 3'h0;
    end else if (_EVAL_55) begin
      _EVAL_92 <= _EVAL_74;
    end else begin
      _EVAL_92 <= _EVAL_75;
    end
    if (_EVAL_152) begin
      _EVAL_112 <= 6'h0;
    end else if (_EVAL_55) begin
      if (_EVAL_52) begin
        _EVAL_112 <= {{1'd0}, _EVAL_144};
      end else begin
        _EVAL_112 <= _EVAL_86;
      end
    end
    if (_EVAL_152) begin
      _EVAL_181 <= _EVAL_8;
    end
    if (_EVAL_152) begin
      _EVAL_187 <= {{34'd0}, _EVAL_228};
    end else if (_EVAL_55) begin
      _EVAL_187 <= {{1'd0}, _EVAL_33};
    end else if (_EVAL_89) begin
      _EVAL_187 <= {{34'd0}, _EVAL_234};
    end else if (_EVAL_247) begin
      _EVAL_187 <= _EVAL_79;
    end
    if (_EVAL_152) begin
      _EVAL_216 <= _EVAL_42;
    end else if (_EVAL_247) begin
      if (_EVAL_201) begin
        _EVAL_216 <= _EVAL_143;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_23 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_61 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_83 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_92 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_112 = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_181 = _RAND_5[4:0];
  _RAND_6 = {3{`RANDOM}};
  _EVAL_187 = _RAND_6[65:0];
  _RAND_7 = {2{`RANDOM}};
  _EVAL_216 = _RAND_7[32:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
