//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_158_assert(
  input        _EVAL,
  input        _EVAL_0,
  input        _EVAL_1,
  input        _EVAL_2,
  input        _EVAL_3,
  input  [8:0] _EVAL_4,
  input  [1:0] _EVAL_5,
  input        _EVAL_6,
  input  [2:0] _EVAL_7,
  input        _EVAL_8,
  input  [1:0] _EVAL_9,
  input        _EVAL_10,
  input  [2:0] _EVAL_11,
  input        _EVAL_12,
  input        _EVAL_13
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_14;
  wire  _EVAL_15;
  wire [1:0] _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire [9:0] _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire [1:0] _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire [31:0] _EVAL_36;
  reg [8:0] _EVAL_37;
  wire [9:0] _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire [31:0] plusarg_reader_out;
  wire [1:0] _EVAL_46;
  wire  _EVAL_47;
  wire [1:0] _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  reg [1:0] _EVAL_51;
  reg [1:0] _EVAL_52;
  wire  _EVAL_53;
  wire [9:0] _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire [9:0] _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire [9:0] _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire [9:0] _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  reg [31:0] _EVAL_82;
  wire [9:0] _EVAL_83;
  wire [8:0] _EVAL_84;
  reg [2:0] _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire [1:0] _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  reg  _EVAL_93;
  wire  _EVAL_94;
  wire [9:0] _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire [9:0] _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire [9:0] _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire [9:0] _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  reg  _EVAL_124;
  wire  _EVAL_125;
  wire [8:0] _EVAL_126;
  wire [8:0] _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire [9:0] _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire [1:0] _EVAL_137;
  wire  _EVAL_138;
  reg  _EVAL_139;
  reg [2:0] _EVAL_140;
  wire [32:0] _EVAL_141;
  wire  _EVAL_142;
  wire [9:0] _EVAL_143;
  wire  _EVAL_144;
  reg  _EVAL_145;
  wire [9:0] _EVAL_146;
  reg  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  reg  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire [8:0] _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire [9:0] _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire [9:0] _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  reg  _EVAL_178;
  wire  _EVAL_179;
  wire [9:0] _EVAL_180;
  wire [8:0] _EVAL_181;
  wire [9:0] _EVAL_182;
  wire  _EVAL_183;
  reg  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire [1:0] _EVAL_199;
  wire [8:0] _EVAL_200;
  wire  _EVAL_201;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_94 = ~_EVAL_178;
  assign _EVAL_24 = ~_EVAL_44;
  assign _EVAL_170 = _EVAL_96 & _EVAL_33;
  assign _EVAL_88 = _EVAL_111 | _EVAL_27;
  assign _EVAL_35 = _EVAL_105 | _EVAL_27;
  assign _EVAL_164 = _EVAL_7 == 3'h7;
  assign _EVAL_153 = ~_EVAL_97;
  assign _EVAL_23 = _EVAL_55 | _EVAL_27;
  assign _EVAL_47 = ~_EVAL_68;
  assign _EVAL_179 = _EVAL_195 | _EVAL_27;
  assign _EVAL_138 = _EVAL_98 | _EVAL_27;
  assign _EVAL_43 = _EVAL_82 < plusarg_reader_out;
  assign _EVAL_80 = ~_EVAL_20;
  assign _EVAL_78 = _EVAL_7 == 3'h6;
  assign _EVAL_150 = $signed(_EVAL_131) == 10'sh0;
  assign _EVAL_71 = _EVAL_2 & _EVAL_153;
  assign _EVAL_54 = $signed(_EVAL_180) & -10'sh40;
  assign _EVAL_115 = _EVAL_172 | _EVAL_150;
  assign _EVAL_73 = _EVAL & _EVAL_148;
  assign _EVAL_28 = ~_EVAL_15;
  assign _EVAL_129 = _EVAL_8 == _EVAL_124;
  assign _EVAL_176 = _EVAL_116 | _EVAL_27;
  assign _EVAL_53 = |_EVAL_147;
  assign _EVAL_133 = _EVAL_7 == 3'h4;
  assign _EVAL_75 = {1'b0,$signed(_EVAL_181)};
  assign _EVAL_17 = ~_EVAL_72;
  assign _EVAL_36 = _EVAL_141[31:0];
  assign _EVAL_20 = _EVAL_45 | _EVAL_27;
  assign _EVAL_174 = _EVAL_2 & _EVAL_164;
  assign _EVAL_155 = _EVAL_4 ^ 9'h44;
  assign _EVAL_201 = _EVAL_48[0];
  assign _EVAL_87 = ~_EVAL_186;
  assign _EVAL_72 = _EVAL_107 | _EVAL_27;
  assign _EVAL_50 = _EVAL_119 | _EVAL_27;
  assign _EVAL_103 = ~_EVAL_201;
  assign _EVAL_90 = _EVAL & _EVAL_106;
  assign _EVAL_69 = $signed(_EVAL_26) & -10'shc;
  assign _EVAL_100 = _EVAL_198 & _EVAL_94;
  assign _EVAL_116 = _EVAL_5 == _EVAL_51;
  assign _EVAL_61 = _EVAL_2 & _EVAL_187;
  assign _EVAL_162 = _EVAL_96 & _EVAL_97;
  assign _EVAL_101 = _EVAL_38;
  assign _EVAL_111 = _EVAL_60 >> _EVAL_0;
  assign _EVAL_148 = _EVAL_11 == 3'h2;
  assign _EVAL_168 = _EVAL_11 == 3'h1;
  assign _EVAL_198 = _EVAL_10 & _EVAL;
  assign _EVAL_191 = ~_EVAL_23;
  assign _EVAL_99 = _EVAL_89[0];
  assign _EVAL_127 = _EVAL_4 ^ 9'h100;
  assign _EVAL_195 = _EVAL_11 <= 3'h6;
  assign _EVAL_30 = ~_EVAL_151;
  assign _EVAL_196 = $signed(_EVAL_101) == 10'sh0;
  assign _EVAL_63 = _EVAL & _EVAL_65;
  assign _EVAL_34 = _EVAL_11 == 3'h4;
  assign _EVAL_83 = _EVAL_143;
  assign _EVAL_143 = $signed(_EVAL_113) & -10'sh8;
  assign _EVAL_130 = _EVAL_32[0];
  assign _EVAL_171 = $signed(_EVAL_79) == 10'sh0;
  assign _EVAL_22 = ~_EVAL_179;
  assign _EVAL_55 = _EVAL_12 == _EVAL_145;
  assign _EVAL_97 = ~_EVAL_93;
  assign _EVAL_21 = ~_EVAL_35;
  assign _EVAL_57 = $signed(_EVAL_83) == 10'sh0;
  assign _EVAL_156 = _EVAL_59 | _EVAL_27;
  assign _EVAL_159 = ~_EVAL_132;
  assign _EVAL_135 = _EVAL_2 & _EVAL_78;
  assign _EVAL_68 = _EVAL_197 | _EVAL_27;
  assign _EVAL_107 = _EVAL_0 == _EVAL_152;
  assign _EVAL_59 = ~_EVAL_8;
  assign _EVAL_144 = _EVAL_9 >= 2'h2;
  assign _EVAL_167 = _EVAL_2 & _EVAL_58;
  assign _EVAL_121 = _EVAL_11 == 3'h6;
  assign _EVAL_132 = _EVAL_134 | _EVAL_27;
  assign _EVAL_131 = _EVAL_169;
  assign _EVAL_41 = ~_EVAL_114;
  assign _EVAL_189 = ~_EVAL_121;
  assign _EVAL_81 = ~_EVAL_138;
  assign _EVAL_177 = _EVAL_144 | _EVAL_27;
  assign _EVAL_65 = ~_EVAL_94;
  assign _EVAL_86 = _EVAL_59 | _EVAL_6;
  assign _EVAL_128 = _EVAL_147 | _EVAL_190;
  assign _EVAL_39 = _EVAL_154 | _EVAL_27;
  assign _EVAL_79 = _EVAL_54;
  assign _EVAL_190 = _EVAL_137[0];
  assign _EVAL_192 = _EVAL_109 | _EVAL_27;
  assign _EVAL_95 = {1'b0,$signed(_EVAL_127)};
  assign _EVAL_98 = _EVAL_175 | _EVAL_43;
  assign _EVAL_56 = ~_EVAL_192;
  assign _EVAL_40 = _EVAL_96 | _EVAL_198;
  assign _EVAL_166 = _EVAL_198 & _EVAL_87;
  assign _EVAL_149 = _EVAL_9 == _EVAL_52;
  assign _EVAL_91 = _EVAL_199[0];
  assign _EVAL_89 = _EVAL_139 - 1'h1;
  assign _EVAL_123 = _EVAL_171 | _EVAL_31;
  assign _EVAL_199 = _EVAL_178 - 1'h1;
  assign _EVAL_46 = _EVAL_186 - 1'h1;
  assign _EVAL_193 = ~_EVAL_177;
  assign _EVAL_137 = _EVAL_170 ? 2'h1 : 2'h0;
  assign _EVAL_142 = ~_EVAL_27;
  assign _EVAL_58 = _EVAL_7 == 3'h1;
  assign _EVAL_74 = _EVAL_5 != 2'h2;
  assign _EVAL_112 = _EVAL_108 | _EVAL_27;
  assign _EVAL_105 = _EVAL_7 == _EVAL_140;
  assign _EVAL_187 = _EVAL_7 == 3'h3;
  assign _EVAL_77 = ~_EVAL_88;
  assign _EVAL_49 = _EVAL_7 == 3'h2;
  assign _EVAL_146 = _EVAL_69;
  assign _EVAL_62 = _EVAL_2 & _EVAL_104;
  assign _EVAL_32 = _EVAL_93 - 1'h1;
  assign _EVAL_38 = $signed(_EVAL_75) & -10'sh20;
  assign _EVAL_96 = _EVAL_3 & _EVAL_2;
  assign _EVAL_158 = _EVAL_4 == _EVAL_37;
  assign _EVAL_25 = _EVAL_2 & _EVAL_133;
  assign _EVAL_122 = ~_EVAL_50;
  assign _EVAL_169 = $signed(_EVAL_182) & -10'sh80;
  assign _EVAL_16 = 2'h1 << _EVAL_0;
  assign _EVAL_183 = ~_EVAL_165;
  assign _EVAL_66 = ~_EVAL_42;
  assign _EVAL_108 = _EVAL_200 == 9'h0;
  assign _EVAL_125 = _EVAL & _EVAL_168;
  assign _EVAL_19 = _EVAL_46[0];
  assign _EVAL_180 = {1'b0,$signed(_EVAL_4)};
  assign _EVAL_48 = _EVAL_173 ? _EVAL_16 : 2'h0;
  assign _EVAL_154 = ~_EVAL_147;
  assign _EVAL_163 = _EVAL_7 == 3'h5;
  assign _EVAL_117 = _EVAL_2 & _EVAL_163;
  assign _EVAL_104 = _EVAL_7 == 3'h0;
  assign _EVAL_84 = _EVAL_4 ^ 9'h58;
  assign _EVAL_70 = ~_EVAL_112;
  assign _EVAL_102 = _EVAL_123 | _EVAL_57;
  assign _EVAL_109 = ~_EVAL_6;
  assign _EVAL_151 = _EVAL_158 | _EVAL_27;
  assign _EVAL_194 = _EVAL & _EVAL_121;
  assign _EVAL_118 = _EVAL_160;
  assign _EVAL_136 = _EVAL_11 == 3'h5;
  assign _EVAL_126 = _EVAL_4 ^ 9'h80;
  assign _EVAL_197 = _EVAL_5 == 2'h0;
  assign _EVAL_188 = _EVAL & _EVAL_136;
  assign _EVAL_76 = _EVAL_2 & _EVAL_49;
  assign _EVAL_175 = _EVAL_67 | _EVAL_14;
  assign _EVAL_181 = _EVAL_4 ^ 9'h60;
  assign _EVAL_182 = {1'b0,$signed(_EVAL_126)};
  assign _EVAL_92 = _EVAL & _EVAL_34;
  assign _EVAL_172 = _EVAL_102 | _EVAL_196;
  assign _EVAL_15 = _EVAL_129 | _EVAL_27;
  assign _EVAL_114 = _EVAL_74 | _EVAL_27;
  assign _EVAL_27 = _EVAL_1;
  assign _EVAL_173 = _EVAL_166 & _EVAL_189;
  assign _EVAL_42 = _EVAL_86 | _EVAL_27;
  assign _EVAL_44 = _EVAL_161 | _EVAL_27;
  assign _EVAL_60 = _EVAL_190 | _EVAL_147;
  assign _EVAL_120 = $signed(_EVAL_118) == 10'sh0;
  assign _EVAL_31 = $signed(_EVAL_146) == 10'sh0;
  assign _EVAL_26 = {1'b0,$signed(_EVAL_155)};
  assign _EVAL_160 = $signed(_EVAL_95) & -10'sh100;
  assign _EVAL_141 = _EVAL_82 + 32'h1;
  assign _EVAL_18 = ~_EVAL_39;
  assign _EVAL_165 = _EVAL_149 | _EVAL_27;
  assign _EVAL_113 = {1'b0,$signed(_EVAL_84)};
  assign _EVAL_119 = _EVAL_5 <= 2'h2;
  assign _EVAL_161 = _EVAL_115 | _EVAL_120;
  assign _EVAL_67 = ~_EVAL_53;
  assign _EVAL_33 = ~_EVAL_139;
  assign _EVAL_106 = _EVAL_11 == 3'h0;
  assign _EVAL_157 = ~_EVAL_156;
  assign _EVAL_14 = plusarg_reader_out == 32'h0;
  assign _EVAL_64 = ~_EVAL_176;
  assign _EVAL_134 = _EVAL_11 == _EVAL_85;
  assign _EVAL_45 = ~_EVAL_0;
  assign _EVAL_200 = _EVAL_4 & 9'h3;
  always @(posedge _EVAL_13) begin
    if (_EVAL_162) begin
      _EVAL_37 <= _EVAL_4;
    end
    if (_EVAL_100) begin
      _EVAL_51 <= _EVAL_5;
    end
    if (_EVAL_100) begin
      _EVAL_52 <= _EVAL_9;
    end
    if (_EVAL_100) begin
      _EVAL_85 <= _EVAL_11;
    end
    if (_EVAL_100) begin
      _EVAL_124 <= _EVAL_8;
    end
    if (_EVAL_162) begin
      _EVAL_140 <= _EVAL_7;
    end
    if (_EVAL_100) begin
      _EVAL_145 <= _EVAL_12;
    end
    if (_EVAL_100) begin
      _EVAL_152 <= _EVAL_0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdb6227f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(def75916)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e71159ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_64) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_66) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af84117c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9d07e2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_64) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(991b6978)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(369edc37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74d3d1ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6c7c094)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45bc21c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f7f0979)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63371720)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d4a86dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44d027cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af44c3e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_157) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b2bf369)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8a60bd3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ab1379c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b855277d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_66) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(860821fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_66) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8f58bb4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7974ea06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8184a20e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d94e844)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bba0fad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(580e0eae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b2013cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_157) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c897384)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a357ca1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eff8ba10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54252c41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cc87288)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38372487)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de88dfcf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccab37b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8ba1183)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(803af8c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81b763be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_66) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_17) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3390c489)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac8286fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3240cdf6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6d37be2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(992bc55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3f7e3a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28632d50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40086447)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84f554a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_173 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab4c0607)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96940ede)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(811d57a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(93736cc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(accf47f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_135 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccab37b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a050b9b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f41724f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c43bee9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7e8f170)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4dfa7445)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a693fbe0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge _EVAL_13 or posedge _EVAL_1) begin
    if (_EVAL_1) begin
      _EVAL_82 <= 32'h0;
    end else if (_EVAL_40) begin
      _EVAL_82 <= 32'h0;
    end else begin
      _EVAL_82 <= _EVAL_36;
    end
  end
  always @(posedge _EVAL_13 or posedge _EVAL_1) begin
    if (_EVAL_1) begin
      _EVAL_93 <= 1'h0;
    end else if (_EVAL_96) begin
      if (_EVAL_97) begin
        _EVAL_93 <= 1'h0;
      end else begin
        _EVAL_93 <= _EVAL_130;
      end
    end
  end
  always @(posedge _EVAL_13 or posedge _EVAL_1) begin
    if (_EVAL_1) begin
      _EVAL_139 <= 1'h0;
    end else if (_EVAL_96) begin
      if (_EVAL_33) begin
        _EVAL_139 <= 1'h0;
      end else begin
        _EVAL_139 <= _EVAL_99;
      end
    end
  end
  always @(posedge _EVAL_13 or posedge _EVAL_1) begin
    if (_EVAL_1) begin
      _EVAL_147 <= 1'h0;
    end else begin
      _EVAL_147 <= _EVAL_128 & _EVAL_103;
    end
  end
  always @(posedge _EVAL_13 or posedge _EVAL_1) begin
    if (_EVAL_1) begin
      _EVAL_178 <= 1'h0;
    end else if (_EVAL_198) begin
      if (_EVAL_94) begin
        _EVAL_178 <= 1'h0;
      end else begin
        _EVAL_178 <= _EVAL_91;
      end
    end
  end
  always @(posedge _EVAL_13 or posedge _EVAL_1) begin
    if (_EVAL_1) begin
      _EVAL_186 <= 1'h0;
    end else if (_EVAL_198) begin
      if (_EVAL_87) begin
        _EVAL_186 <= 1'h0;
      end else begin
        _EVAL_186 <= _EVAL_19;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_37 = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_51 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_52 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_82 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_85 = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_93 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_124 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_139 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_140 = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_145 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_147 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_152 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_178 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_186 = _RAND_13[0:0];
`endif // RANDOMIZE_REG_INIT
  if (_EVAL_1) begin
    _EVAL_82 = 32'h0;
  end
  if (_EVAL_1) begin
    _EVAL_93 = 1'h0;
  end
  if (_EVAL_1) begin
    _EVAL_139 = 1'h0;
  end
  if (_EVAL_1) begin
    _EVAL_147 = 1'h0;
  end
  if (_EVAL_1) begin
    _EVAL_178 = 1'h0;
  end
  if (_EVAL_1) begin
    _EVAL_186 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
