//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_56_assert(
  input  [2:0]  _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [3:0]  _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input  [13:0] _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  input  [4:0]  _EVAL_8,
  input  [2:0]  _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input  [3:0]  _EVAL_13,
  input         _EVAL_14,
  input  [1:0]  _EVAL_15,
  input         _EVAL_16,
  input  [3:0]  _EVAL_17,
  input  [4:0]  _EVAL_18
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_19;
  wire [31:0] _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire [17:0] _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire [3:0] _EVAL_31;
  reg  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire [17:0] _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  reg [2:0] _EVAL_40;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire [3:0] _EVAL_53;
  wire  _EVAL_54;
  wire [13:0] _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  reg [5:0] _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire [1:0] _EVAL_72;
  wire [7:0] _EVAL_73;
  wire  _EVAL_74;
  wire [3:0] _EVAL_75;
  wire [1:0] _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire [17:0] _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire [17:0] _EVAL_90;
  wire [5:0] _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  reg [2:0] _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire [7:0] _EVAL_106;
  wire [5:0] _EVAL_107;
  wire [31:0] _EVAL_108;
  wire  _EVAL_109;
  reg [5:0] _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire [14:0] _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire [7:0] _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire [3:0] _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  reg [5:0] _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  reg [13:0] _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire [6:0] _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire [22:0] _EVAL_165;
  wire  _EVAL_166;
  wire [17:0] _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  reg [3:0] _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire [5:0] _EVAL_173;
  wire [31:0] _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_178;
  wire  _EVAL_179;
  reg  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  reg [17:0] _EVAL_186;
  wire  _EVAL_187;
  wire [17:0] _EVAL_188;
  wire [17:0] _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire [7:0] _EVAL_193;
  wire  _EVAL_194;
  wire [6:0] _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_198;
  wire [13:0] _EVAL_199;
  reg [2:0] _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  reg [3:0] _EVAL_205;
  wire [13:0] _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  reg [4:0] _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire [6:0] _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  reg [4:0] _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  reg [1:0] _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire [17:0] _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire [5:0] _EVAL_251;
  wire  _EVAL_252;
  wire [31:0] _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire [22:0] _EVAL_256;
  wire [1:0] _EVAL_257;
  wire  _EVAL_258;
  wire [14:0] _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire [31:0] _EVAL_265;
  wire [32:0] _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire [5:0] _EVAL_272;
  wire  _EVAL_274;
  reg [5:0] _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire [14:0] _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_294;
  wire  _EVAL_295;
  wire  _EVAL_296;
  wire  _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire [1:0] _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire [6:0] _EVAL_307;
  wire [2:0] _EVAL_308;
  wire [2:0] _EVAL_309;
  wire  _EVAL_310;
  wire  _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_317;
  reg [31:0] _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_320;
  wire  _EVAL_321;
  wire [5:0] _EVAL_322;
  wire  _EVAL_323;
  wire  _EVAL_324;
  wire  _EVAL_325;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_223 = _EVAL_313 | _EVAL_19;
  assign _EVAL_190 = _EVAL_6 == 3'h3;
  assign _EVAL_247 = ~_EVAL_176;
  assign _EVAL_321 = _EVAL_123 & _EVAL_296;
  assign _EVAL_211 = _EVAL_15 == 2'h0;
  assign _EVAL_176 = _EVAL_114 | _EVAL_12;
  assign _EVAL_63 = _EVAL_223 | _EVAL_38;
  assign _EVAL_144 = _EVAL_245 | _EVAL_12;
  assign _EVAL_214 = _EVAL_66 - 6'h1;
  assign _EVAL_309 = _EVAL_18[2:0];
  assign _EVAL_114 = _EVAL_51 | _EVAL_203;
  assign _EVAL_151 = ~_EVAL_241;
  assign _EVAL_59 = _EVAL_8 == 5'h11;
  assign _EVAL_168 = _EVAL <= 3'h2;
  assign _EVAL_71 = ~_EVAL_164;
  assign _EVAL_257 = _EVAL_8[4:3];
  assign _EVAL_204 = _EVAL_172 | _EVAL_12;
  assign _EVAL_130 = {_EVAL_239,_EVAL_109,_EVAL_81,_EVAL_22};
  assign _EVAL_270 = _EVAL_9 == 3'h6;
  assign _EVAL_252 = _EVAL_82 | _EVAL_12;
  assign _EVAL_232 = _EVAL_186 | _EVAL_85;
  assign _EVAL_173 = _EVAL_214[5:0];
  assign _EVAL_125 = _EVAL_264 | _EVAL_12;
  assign _EVAL_206 = _EVAL_5 & _EVAL_55;
  assign _EVAL_307 = _EVAL_275 - 6'h1;
  assign _EVAL_231 = _EVAL_121 | _EVAL_12;
  assign _EVAL_324 = _EVAL_15 == _EVAL_226;
  assign _EVAL_30 = _EVAL_316 & _EVAL_301;
  assign _EVAL_128 = ~_EVAL_142;
  assign _EVAL_277 = _EVAL_9[0];
  assign _EVAL_165 = 23'hff << _EVAL_2;
  assign _EVAL_268 = $signed(_EVAL_119) == 15'sh0;
  assign _EVAL_235 = _EVAL_306 & _EVAL_123;
  assign _EVAL_39 = ~_EVAL_61;
  assign _EVAL_137 = _EVAL_17 >= 4'h2;
  assign _EVAL_241 = _EVAL_104 | _EVAL_12;
  assign _EVAL_299 = _EVAL_287 | _EVAL_12;
  assign _EVAL_221 = _EVAL_2 == _EVAL_205;
  assign _EVAL_178 = _EVAL_211 | _EVAL_12;
  assign _EVAL_100 = _EVAL_6 == 3'h1;
  assign _EVAL_33 = _EVAL_9 == 3'h1;
  assign _EVAL_124 = _EVAL_75 == 4'h0;
  assign _EVAL_44 = 4'h6 == _EVAL_17;
  assign _EVAL_118 = _EVAL_137 | _EVAL_235;
  assign _EVAL_133 = _EVAL_18 == 5'h11;
  assign _EVAL_107 = _EVAL_127[7:2];
  assign _EVAL_228 = _EVAL_157 | _EVAL_12;
  assign _EVAL_35 = _EVAL_186 >> _EVAL_18;
  assign _EVAL_293 = ~_EVAL_156;
  assign _EVAL_185 = _EVAL_5 == _EVAL_150;
  assign _EVAL_143 = _EVAL_9 == 3'h0;
  assign _EVAL_316 = ~_EVAL_123;
  assign _EVAL_102 = _EVAL_136 & _EVAL_19;
  assign _EVAL_300 = ~_EVAL_289;
  assign _EVAL_95 = _EVAL_17[0];
  assign _EVAL_193 = _EVAL_165[7:0];
  assign _EVAL_250 = _EVAL_17 <= 4'hb;
  assign _EVAL_202 = _EVAL_137 | _EVAL_12;
  assign _EVAL_308 = _EVAL_8[2:0];
  assign _EVAL_36 = ~_EVAL_131;
  assign _EVAL_126 = _EVAL_137 | _EVAL_34;
  assign _EVAL_311 = _EVAL_250 & _EVAL_216;
  assign _EVAL_77 = |_EVAL_186;
  assign _EVAL_79 = _EVAL_50 | _EVAL_105;
  assign _EVAL_19 = _EVAL_285 & _EVAL_224;
  assign _EVAL_152 = _EVAL_257 == 2'h0;
  assign _EVAL_53 = ~_EVAL_130;
  assign _EVAL_319 = ~_EVAL_144;
  assign _EVAL_297 = _EVAL_318 < plusarg_reader_out;
  assign _EVAL_115 = _EVAL_67 | _EVAL_12;
  assign _EVAL_97 = _EVAL_183 | _EVAL_12;
  assign _EVAL_306 = _EVAL_302[1];
  assign _EVAL_162 = _EVAL_314 | _EVAL_12;
  assign _EVAL_29 = _EVAL_6[2];
  assign _EVAL_70 = ~_EVAL_231;
  assign _EVAL_237 = ~_EVAL_97;
  assign _EVAL_136 = 4'h2 == _EVAL_17;
  assign _EVAL_169 = _EVAL_141 == 6'h0;
  assign _EVAL_157 = _EVAL <= 3'h3;
  assign _EVAL_27 = _EVAL_85 | _EVAL_186;
  assign _EVAL_272 = _EVAL_106[7:2];
  assign _EVAL_142 = _EVAL_111 | _EVAL_12;
  assign _EVAL_264 = _EVAL != 3'h0;
  assign _EVAL_201 = ~_EVAL_178;
  assign _EVAL_154 = ~_EVAL_11;
  assign _EVAL_127 = ~_EVAL_193;
  assign _EVAL_290 = _EVAL <= 3'h1;
  assign _EVAL_25 = _EVAL_4 & _EVAL_143;
  assign _EVAL_294 = _EVAL_167[0];
  assign _EVAL_90 = _EVAL_232 & _EVAL_188;
  assign _EVAL_50 = _EVAL_85 != _EVAL_189;
  assign _EVAL_166 = _EVAL_6 == 3'h6;
  assign _EVAL_48 = _EVAL_275 == 6'h0;
  assign _EVAL_111 = _EVAL_243 | _EVAL_68;
  assign _EVAL_167 = _EVAL_27 >> _EVAL_8;
  assign _EVAL_96 = _EVAL_262 & _EVAL_268;
  assign _EVAL_87 = _EVAL_227 & _EVAL_69;
  assign _EVAL_161 = ~_EVAL_1;
  assign _EVAL_189 = _EVAL_265[17:0];
  assign _EVAL_298 = _EVAL_6 == _EVAL_103;
  assign _EVAL_145 = _EVAL_17 <= 4'h8;
  assign _EVAL_288 = _EVAL_16 & _EVAL_190;
  assign _EVAL_62 = _EVAL_4 & _EVAL_33;
  assign _EVAL_312 = ~_EVAL_135;
  assign _EVAL_73 = _EVAL_256[7:0];
  assign _EVAL_233 = _EVAL_21 | _EVAL_12;
  assign _EVAL_43 = _EVAL_153 | _EVAL_12;
  assign _EVAL_134 = ~_EVAL_77;
  assign _EVAL_147 = _EVAL_152 & _EVAL_283;
  assign _EVAL_159 = ~_EVAL_146;
  assign _EVAL_238 = ~_EVAL_58;
  assign _EVAL_51 = _EVAL_179 | _EVAL_147;
  assign _EVAL_251 = _EVAL_160[5:0];
  assign _EVAL_20 = 32'h1 << _EVAL_8;
  assign _EVAL_85 = _EVAL_108[17:0];
  assign _EVAL_313 = _EVAL_133 | _EVAL_216;
  assign _EVAL_242 = ~_EVAL_233;
  assign _EVAL_203 = _EVAL_8 == 5'h8;
  assign _EVAL_67 = ~_EVAL_14;
  assign _EVAL_131 = _EVAL_112 | _EVAL_12;
  assign _EVAL_195 = _EVAL_110 - 6'h1;
  assign _EVAL_175 = _EVAL_16 & _EVAL_258;
  assign _EVAL_112 = _EVAL == _EVAL_200;
  assign _EVAL_72 = 2'h1 << _EVAL_95;
  assign _EVAL_116 = ~_EVAL_12;
  assign _EVAL_254 = ~_EVAL_252;
  assign _EVAL_213 = ~_EVAL_202;
  assign _EVAL_207 = _EVAL == 3'h0;
  assign _EVAL_296 = ~_EVAL_301;
  assign _EVAL_260 = ~_EVAL_192;
  assign _EVAL_69 = ~_EVAL_270;
  assign _EVAL_158 = ~_EVAL_249;
  assign _EVAL_263 = _EVAL_8 == 5'h10;
  assign _EVAL_179 = _EVAL_59 | _EVAL_263;
  assign _EVAL_135 = _EVAL_230 | _EVAL_12;
  assign _EVAL_129 = _EVAL_4 & _EVAL_98;
  assign _EVAL_172 = _EVAL_18 == _EVAL_217;
  assign _EVAL_262 = _EVAL_17 <= 4'h2;
  assign _EVAL_224 = _EVAL_309 <= 3'h6;
  assign _EVAL_234 = _EVAL_194 | _EVAL_12;
  assign _EVAL_248 = _EVAL_316 & _EVAL_296;
  assign _EVAL_245 = _EVAL_8 == _EVAL_210;
  assign _EVAL_106 = ~_EVAL_73;
  assign _EVAL_26 = _EVAL_6 == 3'h4;
  assign _EVAL_38 = _EVAL_18 == 5'h8;
  assign _EVAL_284 = _EVAL <= 3'h4;
  assign _EVAL_60 = ~_EVAL_228;
  assign _EVAL_317 = _EVAL_145 & _EVAL_268;
  assign _EVAL_104 = _EVAL_206 == 14'h0;
  assign _EVAL_88 = ~_EVAL_139;
  assign _EVAL_218 = ~_EVAL_271;
  assign _EVAL_49 = _EVAL_6 == 3'h0;
  assign _EVAL_101 = _EVAL_185 | _EVAL_12;
  assign _EVAL_105 = ~_EVAL_24;
  assign _EVAL_139 = _EVAL_246 | _EVAL_12;
  assign _EVAL_45 = _EVAL_37 & _EVAL_321;
  assign _EVAL_295 = _EVAL_28 | _EVAL_12;
  assign _EVAL_187 = ~_EVAL_48;
  assign _EVAL_209 = _EVAL_35[0];
  assign _EVAL_99 = ~_EVAL_94;
  assign _EVAL_322 = _EVAL_195[5:0];
  assign _EVAL_184 = _EVAL_37 & _EVAL_30;
  assign _EVAL_315 = _EVAL_16 & _EVAL_100;
  assign _EVAL_305 = _EVAL_4 & _EVAL_255;
  assign _EVAL_98 = _EVAL_9 == 3'h4;
  assign _EVAL_24 = |_EVAL_85;
  assign _EVAL_196 = _EVAL_168 | _EVAL_12;
  assign _EVAL_289 = _EVAL_207 | _EVAL_12;
  assign _EVAL_109 = _EVAL_118 | _EVAL_45;
  assign _EVAL_215 = ~_EVAL_125;
  assign _EVAL_155 = ~_EVAL_101;
  assign _EVAL_227 = _EVAL_320 & _EVAL_169;
  assign _EVAL_188 = ~_EVAL_189;
  assign _EVAL_194 = _EVAL_2 >= 4'h2;
  assign _EVAL_47 = ~_EVAL_274;
  assign _EVAL_92 = _EVAL_307[5:0];
  assign _EVAL_64 = _EVAL_16 & _EVAL_171;
  assign _EVAL_239 = _EVAL_118 | _EVAL_222;
  assign _EVAL_58 = _EVAL_66 == 6'h0;
  assign _EVAL_120 = ~_EVAL_295;
  assign _EVAL_255 = _EVAL_9 == 3'h5;
  assign _EVAL_54 = _EVAL_276 | _EVAL_320;
  assign _EVAL_42 = _EVAL_16 & _EVAL_49;
  assign _EVAL_93 = _EVAL_4 & _EVAL_270;
  assign _EVAL_75 = ~_EVAL_13;
  assign _EVAL_108 = _EVAL_323 ? _EVAL_174 : 32'h0;
  assign _EVAL_301 = _EVAL_5[0];
  assign _EVAL_274 = _EVAL_154 | _EVAL_12;
  assign _EVAL_119 = _EVAL_281;
  assign _EVAL_222 = _EVAL_37 & _EVAL_113;
  assign _EVAL_220 = plusarg_reader_out == 32'h0;
  assign _EVAL_304 = ~_EVAL_196;
  assign _EVAL_163 = _EVAL_320 & _EVAL_48;
  assign _EVAL_208 = _EVAL_16 & _EVAL_26;
  assign _EVAL_276 = _EVAL_3 & _EVAL_16;
  assign _EVAL_259 = {1'b0,$signed(_EVAL_199)};
  assign _EVAL_267 = _EVAL_4 & _EVAL_187;
  assign _EVAL_291 = _EVAL_317 | _EVAL_12;
  assign _EVAL_84 = _EVAL_16 & _EVAL_166;
  assign _EVAL_113 = _EVAL_123 & _EVAL_301;
  assign _EVAL_283 = _EVAL_308 <= 3'h6;
  assign _EVAL_156 = _EVAL_290 | _EVAL_12;
  assign _EVAL_34 = _EVAL_306 & _EVAL_316;
  assign _EVAL_80 = _EVAL_11 == _EVAL_32;
  assign _EVAL_153 = _EVAL_17 == _EVAL_170;
  assign _EVAL_281 = $signed(_EVAL_259) & -15'sh1000;
  assign _EVAL_55 = {{6'd0}, _EVAL_106};
  assign _EVAL_244 = _EVAL_124 | _EVAL_12;
  assign _EVAL_286 = ~_EVAL_204;
  assign _EVAL_74 = _EVAL_9 == 3'h2;
  assign _EVAL_117 = _EVAL_134 | _EVAL_220;
  assign _EVAL_253 = _EVAL_266[31:0];
  assign _EVAL_52 = _EVAL_37 & _EVAL_248;
  assign _EVAL_68 = _EVAL_44 & _EVAL_38;
  assign _EVAL_78 = _EVAL_16 & _EVAL_238;
  assign _EVAL_132 = _EVAL_262 & _EVAL_46;
  assign _EVAL_37 = _EVAL_302[0];
  assign _EVAL_249 = _EVAL_298 | _EVAL_12;
  assign _EVAL_310 = ~_EVAL_278;
  assign _EVAL_325 = _EVAL_31 == 4'h0;
  assign _EVAL_287 = _EVAL_13 == _EVAL_130;
  assign _EVAL_46 = _EVAL_133 | _EVAL_19;
  assign _EVAL_82 = _EVAL_102 & _EVAL_96;
  assign _EVAL_61 = _EVAL_284 | _EVAL_12;
  assign _EVAL_191 = ~_EVAL_291;
  assign _EVAL_146 = _EVAL_198 | _EVAL_12;
  assign _EVAL_140 = _EVAL_221 | _EVAL_12;
  assign _EVAL_229 = _EVAL_9 <= 3'h6;
  assign _EVAL_199 = _EVAL_5 ^ 14'h3000;
  assign _EVAL_83 = ~_EVAL_234;
  assign _EVAL_183 = _EVAL_15 != 2'h2;
  assign _EVAL_243 = _EVAL_132 | _EVAL_311;
  assign _EVAL_192 = _EVAL_324 | _EVAL_12;
  assign _EVAL_81 = _EVAL_126 | _EVAL_184;
  assign _EVAL_28 = _EVAL_10 == _EVAL_180;
  assign _EVAL_285 = _EVAL_76 == 2'h0;
  assign _EVAL_121 = ~_EVAL_209;
  assign _EVAL_198 = _EVAL_154 | _EVAL_1;
  assign _EVAL_94 = _EVAL_79 | _EVAL_12;
  assign _EVAL_269 = _EVAL_276 & _EVAL_58;
  assign _EVAL_230 = _EVAL_243 & _EVAL_317;
  assign _EVAL_278 = _EVAL_325 | _EVAL_12;
  assign _EVAL_261 = ~_EVAL_115;
  assign _EVAL_256 = 23'hff << _EVAL_17;
  assign _EVAL_171 = _EVAL_6 == 3'h7;
  assign _EVAL_323 = _EVAL_276 & _EVAL_303;
  assign _EVAL_160 = _EVAL_141 - 6'h1;
  assign _EVAL_266 = _EVAL_318 + 32'h1;
  assign _EVAL_282 = ~_EVAL_43;
  assign _EVAL_31 = _EVAL_13 & _EVAL_53;
  assign _EVAL_164 = _EVAL_229 | _EVAL_12;
  assign _EVAL_57 = ~_EVAL_29;
  assign _EVAL_56 = ~_EVAL_122;
  assign _EVAL_86 = _EVAL_16 & _EVAL_279;
  assign _EVAL_314 = _EVAL_117 | _EVAL_297;
  assign _EVAL_271 = _EVAL_161 | _EVAL_12;
  assign _EVAL_265 = _EVAL_87 ? _EVAL_20 : 32'h0;
  assign _EVAL_246 = _EVAL_15 <= 2'h2;
  assign _EVAL_240 = _EVAL_63 | _EVAL_12;
  assign _EVAL_302 = _EVAL_72 | 2'h1;
  assign _EVAL_320 = _EVAL_7 & _EVAL_4;
  assign _EVAL_303 = _EVAL_110 == 6'h0;
  assign _EVAL_292 = ~_EVAL_299;
  assign _EVAL_174 = 32'h1 << _EVAL_18;
  assign _EVAL_22 = _EVAL_126 | _EVAL_52;
  assign _EVAL_236 = ~_EVAL_244;
  assign _EVAL_216 = _EVAL_18 == 5'h10;
  assign _EVAL_212 = ~_EVAL_162;
  assign _EVAL_123 = _EVAL_5[1];
  assign _EVAL_279 = _EVAL_6 == 3'h2;
  assign _EVAL_138 = ~_EVAL_65;
  assign _EVAL_122 = _EVAL_80 | _EVAL_12;
  assign _EVAL_182 = ~_EVAL_240;
  assign _EVAL_21 = _EVAL_9 == _EVAL_40;
  assign _EVAL_76 = _EVAL_18[4:3];
  assign _EVAL_258 = _EVAL_6 == 3'h5;
  assign _EVAL_89 = _EVAL_4 & _EVAL_74;
  assign _EVAL_65 = _EVAL_294 | _EVAL_12;
  assign _EVAL_181 = ~_EVAL_140;
  always @(posedge _EVAL_0) begin
    if (_EVAL_163) begin
      _EVAL_32 <= _EVAL_11;
    end
    if (_EVAL_163) begin
      _EVAL_40 <= _EVAL_9;
    end
    if (_EVAL_12) begin
      _EVAL_66 <= 6'h0;
    end else if (_EVAL_276) begin
      if (_EVAL_58) begin
        if (_EVAL_57) begin
          _EVAL_66 <= _EVAL_272;
        end else begin
          _EVAL_66 <= 6'h0;
        end
      end else begin
        _EVAL_66 <= _EVAL_173;
      end
    end
    if (_EVAL_269) begin
      _EVAL_103 <= _EVAL_6;
    end
    if (_EVAL_12) begin
      _EVAL_110 <= 6'h0;
    end else if (_EVAL_276) begin
      if (_EVAL_303) begin
        if (_EVAL_57) begin
          _EVAL_110 <= _EVAL_272;
        end else begin
          _EVAL_110 <= 6'h0;
        end
      end else begin
        _EVAL_110 <= _EVAL_322;
      end
    end
    if (_EVAL_12) begin
      _EVAL_141 <= 6'h0;
    end else if (_EVAL_320) begin
      if (_EVAL_169) begin
        if (_EVAL_277) begin
          _EVAL_141 <= _EVAL_107;
        end else begin
          _EVAL_141 <= 6'h0;
        end
      end else begin
        _EVAL_141 <= _EVAL_251;
      end
    end
    if (_EVAL_269) begin
      _EVAL_150 <= _EVAL_5;
    end
    if (_EVAL_269) begin
      _EVAL_170 <= _EVAL_17;
    end
    if (_EVAL_163) begin
      _EVAL_180 <= _EVAL_10;
    end
    if (_EVAL_12) begin
      _EVAL_186 <= 18'h0;
    end else begin
      _EVAL_186 <= _EVAL_90;
    end
    if (_EVAL_269) begin
      _EVAL_200 <= _EVAL;
    end
    if (_EVAL_163) begin
      _EVAL_205 <= _EVAL_2;
    end
    if (_EVAL_163) begin
      _EVAL_210 <= _EVAL_8;
    end
    if (_EVAL_269) begin
      _EVAL_217 <= _EVAL_18;
    end
    if (_EVAL_163) begin
      _EVAL_226 <= _EVAL_15;
    end
    if (_EVAL_12) begin
      _EVAL_275 <= 6'h0;
    end else if (_EVAL_320) begin
      if (_EVAL_48) begin
        if (_EVAL_277) begin
          _EVAL_275 <= _EVAL_107;
        end else begin
          _EVAL_275 <= 6'h0;
        end
      end else begin
        _EVAL_275 <= _EVAL_92;
      end
    end
    if (_EVAL_12) begin
      _EVAL_318 <= 32'h0;
    end else if (_EVAL_54) begin
      _EVAL_318 <= 32'h0;
    end else begin
      _EVAL_318 <= _EVAL_253;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_293) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65fe7531)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d9c7a0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_304) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b23c97de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_305 & _EVAL_237) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bf484e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3fe56e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_304) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a2ae11c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5740e4e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(155d3ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(832e05c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0f6cb4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_292) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_292) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_292) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(683b308e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75c149c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_300) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce34ed74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_300) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef1584cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e98ad5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b50e53b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84fc106d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7b82ab4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9fd49a4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_305 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_304) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c67ba299)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_215) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef951629)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(875c2874)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9fcbc2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_310) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fe95341)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eac11f99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a06f583b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab601b39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bcdf0fb3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_237) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(269553af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3ffd589)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_300) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_310) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb16a104)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbc33868)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9c67044)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa8d4e3c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(511c59d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43093589)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_319) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9fd49a4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ec8ea3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26020a73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94b487d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_300) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3cd2de7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71d291f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb5496e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c553881f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_300) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3abf49f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_305 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b212432c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5972b9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3cc23a99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_292) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd28f759)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_305 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bd6106c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5714e903)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_300) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_305 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c5f20b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e2b6dbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a847c8a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_319) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b81d709)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_305 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f93583f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_237) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b201a5e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4f1920b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff7556e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a46c7a7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8be212)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_305 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfd13e56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbc22a12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_305 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c8dcd65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ab80a0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d71a6edd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49398eb2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_215) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d257590)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db64023d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_305 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_305 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b66eb75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cc71201)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42acc934)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91656769)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a341809a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6375235)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad6c3171)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_89 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_267 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eabbc38a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(334d48f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_304) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80fc8412)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_305 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(862b7c51)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_305 & _EVAL_237) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8fcd005f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2dd72362)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_282) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bd92c35)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7afd0998)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f13921)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61023f88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f75d8ce3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_293) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_292) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_4 & _EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55171513)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a307e21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae5367ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15117a6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b74cc88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5596d63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2c5dfd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_32 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_40 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_66 = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_103 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_110 = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_141 = _RAND_5[5:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_150 = _RAND_6[13:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_170 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_180 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_186 = _RAND_9[17:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_200 = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_205 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_210 = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_217 = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_226 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_275 = _RAND_15[5:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_318 = _RAND_16[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
