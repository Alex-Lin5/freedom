//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_93(
  output        _EVAL,
  input  [2:0]  _EVAL_0,
  input  [3:0]  _EVAL_1,
  output [1:0]  _EVAL_2,
  output [31:0] _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  output [2:0]  _EVAL_7,
  output        _EVAL_8,
  output        _EVAL_9,
  output [31:0] _EVAL_10,
  output        _EVAL_11,
  output [14:0] _EVAL_12,
  output [2:0]  _EVAL_13,
  output [4:0]  _EVAL_14,
  input  [14:0] _EVAL_15,
  input         _EVAL_16,
  output [9:0]  _EVAL_17,
  input         _EVAL_18,
  input  [4:0]  _EVAL_19,
  input  [2:0]  _EVAL_20,
  input  [2:0]  _EVAL_21,
  output [3:0]  _EVAL_22,
  input         _EVAL_23,
  input  [31:0] _EVAL_24,
  input  [9:0]  _EVAL_25,
  output [2:0]  _EVAL_26,
  input  [31:0] _EVAL_27,
  input  [2:0]  _EVAL_28,
  input         _EVAL_29,
  output [2:0]  _EVAL_30,
  input  [1:0]  _EVAL_31,
  output        _EVAL_32
);
  wire [2:0] _EVAL_33;
  wire [14:0] _EVAL_34;
  wire  _EVAL_35;
  wire [31:0] _EVAL_36;
  wire [4:0] _EVAL_37;
  wire [2:0] _EVAL_38;
  wire [31:0] _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire [14:0] _EVAL_42;
  wire [4:0] _EVAL_43;
  wire [2:0] _EVAL_44;
  wire  _EVAL_45;
  wire [4:0] _EVAL_46;
  wire [2:0] _EVAL_47;
  wire [2:0] _EVAL_48;
  wire  fragmenter__EVAL;
  wire [2:0] fragmenter__EVAL_0;
  wire  fragmenter__EVAL_1;
  wire  fragmenter__EVAL_2;
  wire [2:0] fragmenter__EVAL_3;
  wire [1:0] fragmenter__EVAL_4;
  wire [9:0] fragmenter__EVAL_5;
  wire [9:0] fragmenter__EVAL_6;
  wire [2:0] fragmenter__EVAL_7;
  wire  fragmenter__EVAL_8;
  wire [2:0] fragmenter__EVAL_9;
  wire [31:0] fragmenter__EVAL_10;
  wire  fragmenter__EVAL_11;
  wire [4:0] fragmenter__EVAL_12;
  wire [1:0] fragmenter__EVAL_13;
  wire [3:0] fragmenter__EVAL_14;
  wire [2:0] fragmenter__EVAL_15;
  wire  fragmenter__EVAL_16;
  wire  fragmenter__EVAL_17;
  wire  fragmenter__EVAL_18;
  wire [3:0] fragmenter__EVAL_19;
  wire [31:0] fragmenter__EVAL_20;
  wire [14:0] fragmenter__EVAL_21;
  wire [2:0] fragmenter__EVAL_22;
  wire [31:0] fragmenter__EVAL_23;
  wire [2:0] fragmenter__EVAL_24;
  wire [31:0] fragmenter__EVAL_25;
  wire  fragmenter__EVAL_26;
  wire  fragmenter__EVAL_27;
  wire [2:0] fragmenter__EVAL_28;
  wire [4:0] fragmenter__EVAL_29;
  wire  fragmenter__EVAL_30;
  wire  fragmenter__EVAL_31;
  wire [14:0] fragmenter__EVAL_32;
  wire [3:0] _EVAL_49;
  wire  _EVAL_50;
  wire [31:0] _EVAL_51;
  wire  _EVAL_52;
  wire [2:0] _EVAL_53;
  wire [2:0] _EVAL_54;
  wire [4:0] _EVAL_55;
  wire  _EVAL_56;
  wire [31:0] _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire [2:0] _EVAL_60;
  wire [2:0] _EVAL_61;
  wire  _EVAL_62;
  wire [3:0] _EVAL_63;
  wire [2:0] _EVAL_64;
  _EVAL_92 fragmenter (
    ._EVAL(fragmenter__EVAL),
    ._EVAL_0(fragmenter__EVAL_0),
    ._EVAL_1(fragmenter__EVAL_1),
    ._EVAL_2(fragmenter__EVAL_2),
    ._EVAL_3(fragmenter__EVAL_3),
    ._EVAL_4(fragmenter__EVAL_4),
    ._EVAL_5(fragmenter__EVAL_5),
    ._EVAL_6(fragmenter__EVAL_6),
    ._EVAL_7(fragmenter__EVAL_7),
    ._EVAL_8(fragmenter__EVAL_8),
    ._EVAL_9(fragmenter__EVAL_9),
    ._EVAL_10(fragmenter__EVAL_10),
    ._EVAL_11(fragmenter__EVAL_11),
    ._EVAL_12(fragmenter__EVAL_12),
    ._EVAL_13(fragmenter__EVAL_13),
    ._EVAL_14(fragmenter__EVAL_14),
    ._EVAL_15(fragmenter__EVAL_15),
    ._EVAL_16(fragmenter__EVAL_16),
    ._EVAL_17(fragmenter__EVAL_17),
    ._EVAL_18(fragmenter__EVAL_18),
    ._EVAL_19(fragmenter__EVAL_19),
    ._EVAL_20(fragmenter__EVAL_20),
    ._EVAL_21(fragmenter__EVAL_21),
    ._EVAL_22(fragmenter__EVAL_22),
    ._EVAL_23(fragmenter__EVAL_23),
    ._EVAL_24(fragmenter__EVAL_24),
    ._EVAL_25(fragmenter__EVAL_25),
    ._EVAL_26(fragmenter__EVAL_26),
    ._EVAL_27(fragmenter__EVAL_27),
    ._EVAL_28(fragmenter__EVAL_28),
    ._EVAL_29(fragmenter__EVAL_29),
    ._EVAL_30(fragmenter__EVAL_30),
    ._EVAL_31(fragmenter__EVAL_31),
    ._EVAL_32(fragmenter__EVAL_32)
  );
  assign fragmenter__EVAL_8 = _EVAL_5;
  assign _EVAL_40 = _EVAL_56;
  assign _EVAL_59 = _EVAL_16;
  assign _EVAL_8 = _EVAL_45;
  assign fragmenter__EVAL_10 = _EVAL_57;
  assign _EVAL_58 = fragmenter__EVAL_1;
  assign _EVAL_35 = _EVAL_62;
  assign _EVAL_50 = fragmenter__EVAL;
  assign _EVAL_3 = fragmenter__EVAL_20;
  assign _EVAL_61 = _EVAL_64;
  assign fragmenter__EVAL_27 = _EVAL_29;
  assign fragmenter__EVAL_21 = _EVAL_42;
  assign _EVAL_63 = _EVAL_1;
  assign fragmenter__EVAL_11 = _EVAL_35;
  assign _EVAL_32 = fragmenter__EVAL_17;
  assign fragmenter__EVAL_9 = _EVAL_47;
  assign _EVAL_34 = _EVAL_15;
  assign _EVAL_45 = _EVAL_58;
  assign _EVAL_56 = _EVAL_18;
  assign _EVAL_54 = _EVAL_21;
  assign fragmenter__EVAL_14 = _EVAL_49;
  assign fragmenter__EVAL_2 = _EVAL_40;
  assign fragmenter__EVAL_4 = _EVAL_31;
  assign _EVAL = fragmenter__EVAL_31;
  assign _EVAL_2 = fragmenter__EVAL_13;
  assign _EVAL_13 = _EVAL_44;
  assign _EVAL_64 = _EVAL_0;
  assign _EVAL_22 = fragmenter__EVAL_19;
  assign _EVAL_53 = _EVAL_33;
  assign _EVAL_38 = _EVAL_54;
  assign _EVAL_42 = _EVAL_34;
  assign _EVAL_49 = _EVAL_63;
  assign _EVAL_57 = _EVAL_51;
  assign _EVAL_55 = _EVAL_19;
  assign fragmenter__EVAL_28 = _EVAL_61;
  assign _EVAL_43 = _EVAL_37;
  assign _EVAL_36 = fragmenter__EVAL_23;
  assign _EVAL_47 = _EVAL_60;
  assign _EVAL_14 = _EVAL_43;
  assign _EVAL_11 = _EVAL_41;
  assign _EVAL_10 = _EVAL_39;
  assign _EVAL_39 = _EVAL_36;
  assign _EVAL_33 = fragmenter__EVAL_3;
  assign _EVAL_30 = fragmenter__EVAL_22;
  assign _EVAL_48 = fragmenter__EVAL_24;
  assign fragmenter__EVAL_16 = _EVAL_6;
  assign fragmenter__EVAL_25 = _EVAL_27;
  assign _EVAL_44 = _EVAL_48;
  assign fragmenter__EVAL_0 = _EVAL_28;
  assign fragmenter__EVAL_12 = _EVAL_46;
  assign _EVAL_7 = _EVAL_53;
  assign fragmenter__EVAL_26 = _EVAL_23;
  assign _EVAL_37 = fragmenter__EVAL_29;
  assign _EVAL_62 = _EVAL_4;
  assign _EVAL_26 = fragmenter__EVAL_7;
  assign _EVAL_51 = _EVAL_24;
  assign fragmenter__EVAL_15 = _EVAL_38;
  assign fragmenter__EVAL_30 = _EVAL_52;
  assign _EVAL_46 = _EVAL_55;
  assign _EVAL_9 = fragmenter__EVAL_18;
  assign _EVAL_52 = _EVAL_59;
  assign fragmenter__EVAL_6 = _EVAL_25;
  assign _EVAL_41 = _EVAL_50;
  assign _EVAL_17 = fragmenter__EVAL_5;
  assign _EVAL_60 = _EVAL_20;
  assign _EVAL_12 = fragmenter__EVAL_32;
endmodule
