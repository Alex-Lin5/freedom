//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_76(
  input         _EVAL,
  input         _EVAL_0,
  output [4:0]  _EVAL_1,
  input  [2:0]  _EVAL_2,
  input  [4:0]  _EVAL_3,
  output [2:0]  _EVAL_4,
  output [2:0]  _EVAL_5,
  output [3:0]  _EVAL_6,
  input  [2:0]  _EVAL_7,
  input  [4:0]  _EVAL_8,
  input  [2:0]  _EVAL_9,
  output [2:0]  _EVAL_10,
  output [1:0]  _EVAL_11,
  output [2:0]  _EVAL_12,
  input  [3:0]  _EVAL_13,
  input  [31:0] _EVAL_14,
  input  [2:0]  _EVAL_15,
  input         _EVAL_16,
  output        _EVAL_17,
  input  [31:0] _EVAL_18,
  input         _EVAL_19,
  input  [31:0] _EVAL_20,
  output [4:0]  _EVAL_21,
  input  [31:0] _EVAL_22,
  output [31:0] _EVAL_23,
  output [4:0]  _EVAL_24,
  output        _EVAL_25,
  output [31:0] _EVAL_26,
  output [1:0]  _EVAL_27,
  output [31:0] _EVAL_28,
  output [31:0] _EVAL_29,
  input  [2:0]  _EVAL_30,
  output [2:0]  _EVAL_31,
  output        _EVAL_32,
  output [2:0]  _EVAL_33,
  input         _EVAL_34,
  input  [2:0]  _EVAL_35,
  input  [1:0]  _EVAL_36,
  output [2:0]  _EVAL_37,
  input  [4:0]  _EVAL_38,
  input  [1:0]  _EVAL_39,
  input  [2:0]  _EVAL_40,
  output [31:0] _EVAL_41,
  output [2:0]  _EVAL_42,
  input         _EVAL_43,
  output        _EVAL_44,
  output [3:0]  _EVAL_45
);
  wire  bundleIn_0_d_sink__EVAL;
  wire [1:0] bundleIn_0_d_sink__EVAL_0;
  wire [2:0] bundleIn_0_d_sink__EVAL_1;
  wire [2:0] bundleIn_0_d_sink__EVAL_2;
  wire [2:0] bundleIn_0_d_sink__EVAL_3;
  wire  bundleIn_0_d_sink__EVAL_4;
  wire  bundleIn_0_d_sink__EVAL_5;
  wire [31:0] bundleIn_0_d_sink__EVAL_6;
  wire [31:0] bundleIn_0_d_sink__EVAL_7;
  wire  bundleIn_0_d_sink__EVAL_8;
  wire [1:0] bundleIn_0_d_sink__EVAL_9;
  wire  bundleIn_0_d_sink__EVAL_10;
  wire [4:0] bundleIn_0_d_sink__EVAL_11;
  wire [2:0] bundleIn_0_d_sink__EVAL_12;
  wire [2:0] bundleIn_0_d_sink__EVAL_13;
  wire [31:0] bundleIn_0_d_sink__EVAL_14;
  wire [2:0] bundleIn_0_d_sink__EVAL_15;
  wire [4:0] bundleIn_0_d_sink__EVAL_16;
  wire [4:0] bundleIn_0_d_sink__EVAL_17;
  wire  bundleIn_0_d_sink__EVAL_18;
  wire [31:0] bundleOut_0_a_source__EVAL;
  wire [31:0] bundleOut_0_a_source__EVAL_0;
  wire [2:0] bundleOut_0_a_source__EVAL_1;
  wire [3:0] bundleOut_0_a_source__EVAL_2;
  wire [31:0] bundleOut_0_a_source__EVAL_3;
  wire [3:0] bundleOut_0_a_source__EVAL_4;
  wire [2:0] bundleOut_0_a_source__EVAL_5;
  wire [2:0] bundleOut_0_a_source__EVAL_6;
  wire [2:0] bundleOut_0_a_source__EVAL_7;
  wire [31:0] bundleOut_0_a_source__EVAL_8;
  wire [1:0] bundleOut_0_a_source__EVAL_9;
  wire [4:0] bundleOut_0_a_source__EVAL_10;
  wire [2:0] bundleOut_0_a_source__EVAL_11;
  wire  bundleOut_0_a_source__EVAL_12;
  wire  bundleOut_0_a_source__EVAL_13;
  wire [2:0] bundleOut_0_a_source__EVAL_14;
  wire [4:0] bundleOut_0_a_source__EVAL_15;
  wire [2:0] bundleOut_0_a_source__EVAL_16;
  wire [1:0] bundleOut_0_a_source__EVAL_17;
  wire  bundleOut_0_a_source__EVAL_18;
  wire [31:0] bundleOut_0_a_source__EVAL_19;
  wire  bundleOut_0_a_source__EVAL_20;
  wire  bundleOut_0_a_source__EVAL_21;
  wire [4:0] bundleOut_0_a_source__EVAL_22;
  wire  bundleOut_0_a_source__EVAL_23;
  wire [31:0] bundleOut_0_a_source__EVAL_24;
  wire [3:0] bundleOut_0_a_source__EVAL_25;
  wire [2:0] bundleOut_0_a_source__EVAL_26;
  wire [2:0] bundleOut_0_a_source__EVAL_27;
  _EVAL_75 bundleIn_0_d_sink (
    ._EVAL(bundleIn_0_d_sink__EVAL),
    ._EVAL_0(bundleIn_0_d_sink__EVAL_0),
    ._EVAL_1(bundleIn_0_d_sink__EVAL_1),
    ._EVAL_2(bundleIn_0_d_sink__EVAL_2),
    ._EVAL_3(bundleIn_0_d_sink__EVAL_3),
    ._EVAL_4(bundleIn_0_d_sink__EVAL_4),
    ._EVAL_5(bundleIn_0_d_sink__EVAL_5),
    ._EVAL_6(bundleIn_0_d_sink__EVAL_6),
    ._EVAL_7(bundleIn_0_d_sink__EVAL_7),
    ._EVAL_8(bundleIn_0_d_sink__EVAL_8),
    ._EVAL_9(bundleIn_0_d_sink__EVAL_9),
    ._EVAL_10(bundleIn_0_d_sink__EVAL_10),
    ._EVAL_11(bundleIn_0_d_sink__EVAL_11),
    ._EVAL_12(bundleIn_0_d_sink__EVAL_12),
    ._EVAL_13(bundleIn_0_d_sink__EVAL_13),
    ._EVAL_14(bundleIn_0_d_sink__EVAL_14),
    ._EVAL_15(bundleIn_0_d_sink__EVAL_15),
    ._EVAL_16(bundleIn_0_d_sink__EVAL_16),
    ._EVAL_17(bundleIn_0_d_sink__EVAL_17),
    ._EVAL_18(bundleIn_0_d_sink__EVAL_18)
  );
  _EVAL_73 bundleOut_0_a_source (
    ._EVAL(bundleOut_0_a_source__EVAL),
    ._EVAL_0(bundleOut_0_a_source__EVAL_0),
    ._EVAL_1(bundleOut_0_a_source__EVAL_1),
    ._EVAL_2(bundleOut_0_a_source__EVAL_2),
    ._EVAL_3(bundleOut_0_a_source__EVAL_3),
    ._EVAL_4(bundleOut_0_a_source__EVAL_4),
    ._EVAL_5(bundleOut_0_a_source__EVAL_5),
    ._EVAL_6(bundleOut_0_a_source__EVAL_6),
    ._EVAL_7(bundleOut_0_a_source__EVAL_7),
    ._EVAL_8(bundleOut_0_a_source__EVAL_8),
    ._EVAL_9(bundleOut_0_a_source__EVAL_9),
    ._EVAL_10(bundleOut_0_a_source__EVAL_10),
    ._EVAL_11(bundleOut_0_a_source__EVAL_11),
    ._EVAL_12(bundleOut_0_a_source__EVAL_12),
    ._EVAL_13(bundleOut_0_a_source__EVAL_13),
    ._EVAL_14(bundleOut_0_a_source__EVAL_14),
    ._EVAL_15(bundleOut_0_a_source__EVAL_15),
    ._EVAL_16(bundleOut_0_a_source__EVAL_16),
    ._EVAL_17(bundleOut_0_a_source__EVAL_17),
    ._EVAL_18(bundleOut_0_a_source__EVAL_18),
    ._EVAL_19(bundleOut_0_a_source__EVAL_19),
    ._EVAL_20(bundleOut_0_a_source__EVAL_20),
    ._EVAL_21(bundleOut_0_a_source__EVAL_21),
    ._EVAL_22(bundleOut_0_a_source__EVAL_22),
    ._EVAL_23(bundleOut_0_a_source__EVAL_23),
    ._EVAL_24(bundleOut_0_a_source__EVAL_24),
    ._EVAL_25(bundleOut_0_a_source__EVAL_25),
    ._EVAL_26(bundleOut_0_a_source__EVAL_26),
    ._EVAL_27(bundleOut_0_a_source__EVAL_27)
  );
  assign bundleIn_0_d_sink__EVAL_13 = _EVAL_40;
  assign _EVAL_29 = bundleOut_0_a_source__EVAL_0;
  assign bundleOut_0_a_source__EVAL_22 = _EVAL_38;
  assign _EVAL_33 = bundleIn_0_d_sink__EVAL_2;
  assign bundleIn_0_d_sink__EVAL_14 = _EVAL_20;
  assign _EVAL_41 = bundleIn_0_d_sink__EVAL_7;
  assign bundleIn_0_d_sink__EVAL_18 = _EVAL_0;
  assign _EVAL_5 = bundleIn_0_d_sink__EVAL_1;
  assign _EVAL_27 = bundleOut_0_a_source__EVAL_9;
  assign _EVAL_28 = bundleOut_0_a_source__EVAL_3;
  assign bundleIn_0_d_sink__EVAL_15 = _EVAL_30;
  assign bundleOut_0_a_source__EVAL_12 = _EVAL;
  assign _EVAL_42 = bundleOut_0_a_source__EVAL_11;
  assign _EVAL_24 = bundleOut_0_a_source__EVAL_15;
  assign bundleOut_0_a_source__EVAL_18 = _EVAL_43;
  assign _EVAL_4 = bundleOut_0_a_source__EVAL_7;
  assign _EVAL_21 = bundleOut_0_a_source__EVAL_10;
  assign _EVAL_31 = bundleOut_0_a_source__EVAL_26;
  assign _EVAL_37 = bundleOut_0_a_source__EVAL_1;
  assign _EVAL_6 = bundleOut_0_a_source__EVAL_25;
  assign bundleOut_0_a_source__EVAL_6 = _EVAL_35;
  assign bundleOut_0_a_source__EVAL_4 = _EVAL_13;
  assign _EVAL_1 = bundleIn_0_d_sink__EVAL_11;
  assign bundleIn_0_d_sink__EVAL_12 = _EVAL_2;
  assign bundleIn_0_d_sink__EVAL_8 = _EVAL_43;
  assign _EVAL_12 = bundleOut_0_a_source__EVAL_14;
  assign bundleOut_0_a_source__EVAL_13 = _EVAL_19;
  assign bundleOut_0_a_source__EVAL_16 = _EVAL_9;
  assign bundleOut_0_a_source__EVAL_27 = _EVAL_15;
  assign bundleIn_0_d_sink__EVAL_17 = _EVAL_8;
  assign bundleOut_0_a_source__EVAL_8 = _EVAL_22;
  assign _EVAL_45 = bundleOut_0_a_source__EVAL_2;
  assign bundleIn_0_d_sink__EVAL = _EVAL;
  assign _EVAL_11 = bundleIn_0_d_sink__EVAL_0;
  assign _EVAL_23 = bundleOut_0_a_source__EVAL_19;
  assign _EVAL_32 = bundleOut_0_a_source__EVAL_20;
  assign bundleIn_0_d_sink__EVAL_9 = _EVAL_39;
  assign bundleOut_0_a_source__EVAL = _EVAL_18;
  assign bundleIn_0_d_sink__EVAL_6 = _EVAL_14;
  assign bundleIn_0_d_sink__EVAL_3 = _EVAL_7;
  assign _EVAL_17 = bundleIn_0_d_sink__EVAL_10;
  assign bundleIn_0_d_sink__EVAL_5 = _EVAL_16;
  assign bundleOut_0_a_source__EVAL_21 = _EVAL_34;
  assign bundleOut_0_a_source__EVAL_17 = _EVAL_36;
  assign _EVAL_25 = bundleIn_0_d_sink__EVAL_4;
  assign _EVAL_44 = bundleOut_0_a_source__EVAL_23;
  assign _EVAL_26 = bundleOut_0_a_source__EVAL_24;
  assign _EVAL_10 = bundleOut_0_a_source__EVAL_5;
  assign bundleIn_0_d_sink__EVAL_16 = _EVAL_3;
endmodule
