//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_37(
  output [2:0]  _EVAL,
  input         _EVAL_0,
  input  [2:0]  _EVAL_1,
  input         _EVAL_2,
  output        _EVAL_3,
  output        _EVAL_4,
  input  [3:0]  _EVAL_5,
  input  [1:0]  _EVAL_6,
  output [3:0]  _EVAL_7,
  output        _EVAL_8,
  input  [3:0]  _EVAL_9,
  output [31:0] _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  output        _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  output [31:0] _EVAL_16,
  input  [3:0]  _EVAL_17,
  output        _EVAL_18,
  input         _EVAL_19,
  input         _EVAL_20,
  output        _EVAL_21,
  input         _EVAL_22,
  input  [31:0] _EVAL_23,
  input         _EVAL_24,
  input  [31:0] _EVAL_25,
  output [31:0] _EVAL_26,
  output        _EVAL_27,
  input         _EVAL_28,
  input         _EVAL_29,
  input         _EVAL_30,
  input         _EVAL_31,
  output        _EVAL_32,
  input  [31:0] _EVAL_33,
  output        _EVAL_34,
  output [3:0]  _EVAL_35,
  input         _EVAL_36,
  output        _EVAL_37
);
  assign _EVAL_16 = _EVAL_23;
  assign _EVAL_21 = _EVAL_36;
  assign _EVAL_27 = _EVAL_20;
  assign _EVAL_35 = _EVAL_17;
  assign _EVAL_13 = _EVAL_22;
  assign _EVAL_10 = _EVAL_25;
  assign _EVAL_7 = _EVAL_9;
  assign _EVAL_26 = _EVAL_33;
  assign _EVAL_3 = _EVAL_29;
  assign _EVAL_18 = _EVAL_2;
  assign _EVAL_4 = _EVAL_14;
  assign _EVAL = _EVAL_1;
  assign _EVAL_32 = _EVAL_30;
  assign _EVAL_8 = _EVAL_28;
  assign _EVAL_34 = _EVAL_24;
  assign _EVAL_37 = _EVAL_31;
endmodule
