//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_81_assert(
  input  [1:0]  _EVAL,
  input  [2:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  input  [1:0]  _EVAL_4,
  input         _EVAL_5,
  input  [9:0]  _EVAL_6,
  input         _EVAL_7,
  input  [9:0]  _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input  [1:0]  _EVAL_11,
  input  [29:0] _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input  [3:0]  _EVAL_16,
  input         _EVAL_17,
  input  [2:0]  _EVAL_18
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [575:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire [1023:0] _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire [1:0] _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire [1:0] _EVAL_31;
  wire [1:0] _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire [575:0] _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  reg [2:0] _EVAL_56;
  wire [3:0] _EVAL_57;
  wire [1:0] _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  reg  _EVAL_62;
  wire  _EVAL_63;
  reg  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  reg  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire [575:0] _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire [1023:0] _EVAL_77;
  reg [575:0] _EVAL_78;
  wire  _EVAL_79;
  wire [575:0] _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  reg [31:0] _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  reg [1:0] _EVAL_96;
  wire [32:0] _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  reg  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire [575:0] _EVAL_112;
  wire  _EVAL_113;
  wire [1023:0] _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  reg [29:0] _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire [3:0] _EVAL_126;
  wire  _EVAL_127;
  reg [9:0] _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire [30:0] _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_136;
  reg [2:0] _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire [30:0] _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire [575:0] _EVAL_143;
  wire  _EVAL_144;
  reg [1:0] _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire [1:0] _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire [3:0] _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire [1:0] _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire [29:0] _EVAL_169;
  wire  _EVAL_170;
  wire [1023:0] _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire [31:0] plusarg_reader_out;
  reg [9:0] _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire [29:0] _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  reg [2:0] _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  reg  _EVAL_193;
  wire [575:0] _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_199;
  wire [1:0] _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_206;
  wire  _EVAL_207;
  reg  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  reg [1:0] _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire [575:0] _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire [29:0] _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire [31:0] _EVAL_232;
  wire [3:0] _EVAL_233;
  wire  _EVAL_234;
  wire [1:0] _EVAL_235;
  wire [30:0] _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire [575:0] _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_262;
  wire [4:0] _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_245 = ~_EVAL_162;
  assign _EVAL_31 = _EVAL_69 - 1'h1;
  assign _EVAL_29 = _EVAL >= 2'h2;
  assign _EVAL_36 = _EVAL_204 | _EVAL_14;
  assign _EVAL_214 = ~_EVAL_252;
  assign _EVAL_44 = _EVAL_91 | _EVAL_14;
  assign _EVAL_224 = _EVAL_12 & _EVAL_169;
  assign _EVAL_256 = _EVAL_226 | _EVAL_14;
  assign _EVAL_74 = _EVAL_191 | _EVAL_130;
  assign _EVAL_114 = 1024'h1 << _EVAL_8;
  assign _EVAL_154 = _EVAL_16 & _EVAL_57;
  assign _EVAL_139 = _EVAL_0 == 3'h6;
  assign _EVAL_152 = _EVAL_52 | _EVAL_14;
  assign _EVAL_173 = $signed(_EVAL_140) == 31'sh0;
  assign _EVAL_263 = 5'h3 << _EVAL_4;
  assign _EVAL_100 = _EVAL_8 == _EVAL_128;
  assign _EVAL_150 = _EVAL_9 & _EVAL_219;
  assign _EVAL_215 = _EVAL_87 < plusarg_reader_out;
  assign _EVAL_88 = _EVAL_4 <= 2'h2;
  assign _EVAL_138 = _EVAL_4 >= 2'h2;
  assign _EVAL_174 = _EVAL_11 != 2'h2;
  assign _EVAL_161 = _EVAL_28 & _EVAL_94;
  assign _EVAL_199 = _EVAL_243 | _EVAL_14;
  assign _EVAL_22 = ~_EVAL_238;
  assign _EVAL_34 = _EVAL_32[0];
  assign _EVAL_155 = _EVAL_233 == 4'h0;
  assign _EVAL_77 = _EVAL_113 ? _EVAL_114 : 1024'h0;
  assign _EVAL_116 = ~_EVAL_172;
  assign _EVAL_151 = _EVAL_1 & _EVAL_229;
  assign _EVAL_177 = _EVAL_103 & _EVAL_22;
  assign _EVAL_131 = _EVAL_224 == 30'h0;
  assign _EVAL_244 = ~_EVAL_115;
  assign _EVAL_92 = _EVAL_8 <= 10'h23f;
  assign _EVAL_169 = {{28'd0}, _EVAL_235};
  assign _EVAL_182 = _EVAL_9 & _EVAL_123;
  assign _EVAL_39 = _EVAL_138 | _EVAL_146;
  assign _EVAL_94 = ~_EVAL_64;
  assign _EVAL_168 = _EVAL_187 | _EVAL_14;
  assign _EVAL_274 = _EVAL_3 == 3'h6;
  assign _EVAL_204 = _EVAL_4 == _EVAL_96;
  assign _EVAL_192 = ~_EVAL_199;
  assign _EVAL_35 = _EVAL_112 & _EVAL_241;
  assign _EVAL_210 = ~_EVAL_2;
  assign _EVAL_134 = _EVAL_237 | _EVAL_14;
  assign _EVAL_113 = _EVAL_260 & _EVAL_186;
  assign _EVAL_188 = _EVAL_11 == 2'h0;
  assign _EVAL_73 = _EVAL_195 >> _EVAL_8;
  assign _EVAL_268 = _EVAL_28 | _EVAL_221;
  assign _EVAL_50 = _EVAL_227 & _EVAL_103;
  assign _EVAL_68 = _EVAL_159 | _EVAL_14;
  assign _EVAL_98 = ~_EVAL_44;
  assign _EVAL_46 = _EVAL_39 | _EVAL_67;
  assign _EVAL_183 = _EVAL_12 ^ 30'h20000000;
  assign _EVAL_202 = ~_EVAL_13;
  assign _EVAL_216 = _EVAL_0 == 3'h1;
  assign _EVAL_33 = _EVAL_6 == _EVAL_175;
  assign _EVAL_93 = _EVAL_9 & _EVAL_185;
  assign _EVAL_28 = _EVAL_15 & _EVAL_9;
  assign _EVAL_89 = ~_EVAL_158;
  assign _EVAL_103 = ~_EVAL_222;
  assign _EVAL_184 = _EVAL_88 & _EVAL_173;
  assign _EVAL_233 = ~_EVAL_16;
  assign _EVAL_212 = _EVAL_117 | _EVAL_14;
  assign _EVAL_255 = ~_EVAL_79;
  assign _EVAL_228 = _EVAL_206 | _EVAL_14;
  assign _EVAL_106 = _EVAL_39 | _EVAL_51;
  assign _EVAL_142 = ~_EVAL_109;
  assign _EVAL_82 = _EVAL_24 | _EVAL_14;
  assign _EVAL_191 = ~_EVAL_76;
  assign _EVAL_136 = _EVAL_9 & _EVAL_38;
  assign _EVAL_276 = _EVAL_1 & _EVAL_245;
  assign _EVAL_230 = _EVAL_34 & _EVAL_95;
  assign _EVAL_181 = _EVAL_29 | _EVAL_14;
  assign _EVAL_65 = _EVAL == _EVAL_145;
  assign _EVAL_115 = _EVAL_25 | _EVAL_14;
  assign _EVAL_60 = _EVAL_18 <= 3'h4;
  assign _EVAL_23 = _EVAL_178 ? _EVAL_171 : 1024'h0;
  assign _EVAL_144 = ~_EVAL_147;
  assign _EVAL_278 = _EVAL_100 | _EVAL_14;
  assign _EVAL_176 = _EVAL_3 == 3'h0;
  assign _EVAL_266 = _EVAL_154 == 4'h0;
  assign _EVAL_55 = ~_EVAL_42;
  assign _EVAL_248 = _EVAL_163[0];
  assign _EVAL_226 = _EVAL_18 != 3'h0;
  assign _EVAL_231 = _EVAL_138 | _EVAL_50;
  assign _EVAL_147 = _EVAL_174 | _EVAL_14;
  assign _EVAL_51 = _EVAL_34 & _EVAL_207;
  assign _EVAL_159 = _EVAL_74 | _EVAL_215;
  assign _EVAL_253 = ~_EVAL_141;
  assign _EVAL_75 = ~_EVAL_47;
  assign _EVAL_236 = $signed(_EVAL_133) & -31'sh2000;
  assign _EVAL_124 = ~_EVAL_119;
  assign _EVAL_70 = ~_EVAL_129;
  assign _EVAL_97 = _EVAL_87 + 32'h1;
  assign _EVAL_203 = _EVAL_9 & _EVAL_251;
  assign _EVAL_26 = _EVAL_62 - 1'h1;
  assign _EVAL_81 = ~_EVAL_228;
  assign _EVAL_133 = {1'b0,$signed(_EVAL_183)};
  assign _EVAL_52 = _EVAL_18 == 3'h0;
  assign _EVAL_54 = ~_EVAL_37;
  assign _EVAL_41 = _EVAL_1 & _EVAL_105;
  assign _EVAL_227 = _EVAL_32[1];
  assign _EVAL_126 = {_EVAL_106,_EVAL_46,_EVAL_179,_EVAL_270};
  assign _EVAL_247 = ~_EVAL_72;
  assign _EVAL_207 = _EVAL_222 & _EVAL_238;
  assign _EVAL_101 = ~_EVAL_14;
  assign _EVAL_249 = _EVAL_18 <= 3'h2;
  assign _EVAL_149 = _EVAL_65 | _EVAL_14;
  assign _EVAL_260 = _EVAL_221 & _EVAL_156;
  assign _EVAL_275 = ~_EVAL_36;
  assign _EVAL_110 = ~_EVAL_149;
  assign _EVAL_277 = _EVAL_1 & _EVAL_157;
  assign _EVAL_79 = _EVAL_155 | _EVAL_14;
  assign _EVAL_246 = ~_EVAL_212;
  assign _EVAL_273 = _EVAL_0 == 3'h5;
  assign _EVAL_72 = _EVAL_257 | _EVAL_14;
  assign _EVAL_180 = ~_EVAL_104;
  assign _EVAL_129 = _EVAL_164 | _EVAL_14;
  assign _EVAL_38 = _EVAL_0 == 3'h4;
  assign _EVAL_32 = _EVAL_148 | 2'h1;
  assign _EVAL_221 = _EVAL_17 & _EVAL_1;
  assign _EVAL_85 = _EVAL_202 | _EVAL_14;
  assign _EVAL_57 = ~_EVAL_126;
  assign _EVAL_109 = _EVAL_138 | _EVAL_14;
  assign _EVAL_127 = ~_EVAL_99;
  assign _EVAL_240 = ~_EVAL_102;
  assign _EVAL_121 = ~_EVAL_68;
  assign _EVAL_123 = ~_EVAL_94;
  assign _EVAL_170 = ~_EVAL_209;
  assign _EVAL_125 = ~_EVAL_165;
  assign _EVAL_118 = ~_EVAL_168;
  assign _EVAL_164 = _EVAL_11 == _EVAL_211;
  assign _EVAL_59 = _EVAL_3 == _EVAL_190;
  assign _EVAL_102 = _EVAL_218[0];
  assign _EVAL_217 = ~_EVAL_108;
  assign _EVAL_25 = ~_EVAL_7;
  assign _EVAL_37 = _EVAL_188 | _EVAL_14;
  assign _EVAL_201 = _EVAL_26[0];
  assign _EVAL_148 = 2'h1 << _EVAL_120;
  assign _EVAL_80 = _EVAL_23[575:0];
  assign _EVAL_104 = |_EVAL_80;
  assign _EVAL_99 = _EVAL_213 | _EVAL_14;
  assign _EVAL_262 = _EVAL_9 & _EVAL_216;
  assign _EVAL_167 = _EVAL_267 | _EVAL_14;
  assign _EVAL_90 = _EVAL_1 & _EVAL_274;
  assign _EVAL_43 = ~_EVAL_196;
  assign _EVAL_235 = ~_EVAL_58;
  assign _EVAL_258 = _EVAL_3 == 3'h1;
  assign _EVAL_234 = _EVAL_5 == _EVAL_193;
  assign _EVAL_250 = ~_EVAL_82;
  assign _EVAL_189 = ~_EVAL_85;
  assign _EVAL_162 = ~_EVAL_69;
  assign _EVAL_218 = _EVAL_78 >> _EVAL_6;
  assign _EVAL_84 = _EVAL_0 == 3'h3;
  assign _EVAL_71 = ~_EVAL_152;
  assign _EVAL_83 = _EVAL_1 & _EVAL_258;
  assign _EVAL_48 = _EVAL_9 & _EVAL_139;
  assign _EVAL_156 = ~_EVAL_208;
  assign _EVAL_223 = ~_EVAL_134;
  assign _EVAL_30 = ~_EVAL_167;
  assign _EVAL_272 = _EVAL_80 != _EVAL_143;
  assign _EVAL_178 = _EVAL_28 & _EVAL_63;
  assign _EVAL_24 = _EVAL_18 == _EVAL_56;
  assign _EVAL_157 = _EVAL_3 == 3'h5;
  assign _EVAL_219 = _EVAL_0 == 3'h7;
  assign _EVAL_172 = _EVAL_59 | _EVAL_14;
  assign _EVAL_200 = _EVAL_64 - 1'h1;
  assign _EVAL_187 = _EVAL_91 & _EVAL_184;
  assign _EVAL_86 = _EVAL_266 | _EVAL_14;
  assign _EVAL_271 = _EVAL_9 & _EVAL_273;
  assign _EVAL_196 = _EVAL_92 | _EVAL_14;
  assign _EVAL_251 = _EVAL_0 == 3'h0;
  assign _EVAL_20 = ~_EVAL_264;
  assign _EVAL_146 = _EVAL_227 & _EVAL_222;
  assign _EVAL_91 = _EVAL_6 <= 10'h23f;
  assign _EVAL_232 = _EVAL_97[31:0];
  assign _EVAL_111 = _EVAL_18 <= 3'h1;
  assign _EVAL_63 = ~_EVAL_62;
  assign _EVAL_213 = _EVAL_7 == _EVAL_107;
  assign _EVAL_40 = _EVAL_12 == _EVAL_122;
  assign _EVAL_153 = _EVAL_111 | _EVAL_14;
  assign _EVAL_270 = _EVAL_231 | _EVAL_66;
  assign _EVAL_120 = _EVAL_4[0];
  assign _EVAL_186 = ~_EVAL_274;
  assign _EVAL_45 = ~_EVAL_153;
  assign _EVAL_171 = 1024'h1 << _EVAL_6;
  assign _EVAL_243 = _EVAL_11 <= 2'h2;
  assign _EVAL_47 = _EVAL_166 | _EVAL_14;
  assign _EVAL_132 = _EVAL_3 <= 3'h6;
  assign _EVAL_267 = _EVAL_272 | _EVAL_180;
  assign _EVAL_163 = _EVAL_208 - 1'h1;
  assign _EVAL_119 = _EVAL_40 | _EVAL_14;
  assign _EVAL_27 = _EVAL_31[0];
  assign _EVAL_140 = _EVAL_236;
  assign _EVAL_67 = _EVAL_34 & _EVAL_254;
  assign _EVAL_239 = _EVAL_9 & _EVAL_84;
  assign _EVAL_143 = _EVAL_77[575:0];
  assign _EVAL_130 = plusarg_reader_out == 32'h0;
  assign _EVAL_105 = _EVAL_3 == 3'h4;
  assign _EVAL_237 = _EVAL_25 | _EVAL_13;
  assign _EVAL_206 = _EVAL_16 == _EVAL_126;
  assign _EVAL_257 = _EVAL_18 <= 3'h3;
  assign _EVAL_158 = _EVAL_240 | _EVAL_14;
  assign _EVAL_254 = _EVAL_222 & _EVAL_22;
  assign _EVAL_95 = _EVAL_103 & _EVAL_238;
  assign _EVAL_76 = |_EVAL_78;
  assign _EVAL_49 = _EVAL_131 | _EVAL_14;
  assign _EVAL_53 = ~_EVAL_278;
  assign _EVAL_222 = _EVAL_12[1];
  assign _EVAL_66 = _EVAL_34 & _EVAL_177;
  assign _EVAL_241 = ~_EVAL_143;
  assign _EVAL_179 = _EVAL_231 | _EVAL_230;
  assign _EVAL_141 = _EVAL_184 | _EVAL_14;
  assign _EVAL_252 = _EVAL_234 | _EVAL_14;
  assign _EVAL_42 = _EVAL_132 | _EVAL_14;
  assign _EVAL_195 = _EVAL_80 | _EVAL_78;
  assign _EVAL_259 = _EVAL_221 & _EVAL_162;
  assign _EVAL_209 = _EVAL_249 | _EVAL_14;
  assign _EVAL_112 = _EVAL_78 | _EVAL_80;
  assign _EVAL_117 = _EVAL_0 == _EVAL_137;
  assign _EVAL_58 = _EVAL_263[1:0];
  assign _EVAL_19 = _EVAL_1 & _EVAL_176;
  assign _EVAL_220 = ~_EVAL_256;
  assign _EVAL_185 = _EVAL_0 == 3'h2;
  assign _EVAL_21 = ~_EVAL_181;
  assign _EVAL_242 = _EVAL_200[0];
  assign _EVAL_225 = ~_EVAL_86;
  assign _EVAL_264 = _EVAL_60 | _EVAL_14;
  assign _EVAL_160 = ~_EVAL_49;
  assign _EVAL_166 = _EVAL_73[0];
  assign _EVAL_165 = _EVAL_210 | _EVAL_14;
  assign _EVAL_238 = _EVAL_12[0];
  assign _EVAL_108 = _EVAL_33 | _EVAL_14;
  assign _EVAL_229 = _EVAL_3 == 3'h2;
  always @(posedge _EVAL_10) begin
    if (_EVAL_161) begin
      _EVAL_56 <= _EVAL_18;
    end
    if (_EVAL_14) begin
      _EVAL_62 <= 1'h0;
    end else if (_EVAL_28) begin
      if (_EVAL_63) begin
        _EVAL_62 <= 1'h0;
      end else begin
        _EVAL_62 <= _EVAL_201;
      end
    end
    if (_EVAL_14) begin
      _EVAL_64 <= 1'h0;
    end else if (_EVAL_28) begin
      if (_EVAL_94) begin
        _EVAL_64 <= 1'h0;
      end else begin
        _EVAL_64 <= _EVAL_242;
      end
    end
    if (_EVAL_14) begin
      _EVAL_69 <= 1'h0;
    end else if (_EVAL_221) begin
      if (_EVAL_162) begin
        _EVAL_69 <= 1'h0;
      end else begin
        _EVAL_69 <= _EVAL_27;
      end
    end
    if (_EVAL_14) begin
      _EVAL_78 <= 576'h0;
    end else begin
      _EVAL_78 <= _EVAL_35;
    end
    if (_EVAL_14) begin
      _EVAL_87 <= 32'h0;
    end else if (_EVAL_268) begin
      _EVAL_87 <= 32'h0;
    end else begin
      _EVAL_87 <= _EVAL_232;
    end
    if (_EVAL_161) begin
      _EVAL_96 <= _EVAL_4;
    end
    if (_EVAL_259) begin
      _EVAL_107 <= _EVAL_7;
    end
    if (_EVAL_161) begin
      _EVAL_122 <= _EVAL_12;
    end
    if (_EVAL_259) begin
      _EVAL_128 <= _EVAL_8;
    end
    if (_EVAL_161) begin
      _EVAL_137 <= _EVAL_0;
    end
    if (_EVAL_259) begin
      _EVAL_145 <= _EVAL;
    end
    if (_EVAL_161) begin
      _EVAL_175 <= _EVAL_6;
    end
    if (_EVAL_259) begin
      _EVAL_190 <= _EVAL_3;
    end
    if (_EVAL_259) begin
      _EVAL_193 <= _EVAL_5;
    end
    if (_EVAL_14) begin
      _EVAL_208 <= 1'h0;
    end else if (_EVAL_221) begin
      if (_EVAL_156) begin
        _EVAL_208 <= 1'h0;
      end else begin
        _EVAL_208 <= _EVAL_248;
      end
    end
    if (_EVAL_259) begin
      _EVAL_211 <= _EVAL_11;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c01cae7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd37cea9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(feff41ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d2f3466)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_250) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1088a42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d114cc0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(117d87c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(260fd863)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_253) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77f61228)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59bf152b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76f71e1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(540f64aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(665b4840)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce85b946)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4290de67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b95532ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa421194)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1de76200)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52b2e2a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(819a2667)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82c0c7c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37aea240)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_220) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_220) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94e120a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(404320b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5288db8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4faa77aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ae0290e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa3a434)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48ab0bbc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_275) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b961c1c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d64764d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfd461e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d9387b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ad6b0b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_255) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95953ca3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_30) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e48de12e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7fa6ce29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d8738a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9fd7f7ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca52da7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1325c2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ab42f07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aebff07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_253) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9921abef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7645bedf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81204d87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_275) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84b10db1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_30) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a2ff4b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_81) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e14afdc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3f03f68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3c82d7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_53) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3846071)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_247) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3570f9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61d2bd1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(523f6eb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45efb0a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35dad8c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_53) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec00e024)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_81) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7136261)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1d676e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(565068fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b8df004)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(875fb59b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(565f446d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4edf73a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_253) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8caa653f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a05bed93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_255) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(359740a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45a2f2fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_255) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f44d19b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c335f8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdb9af3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ec3cb3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d2057d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89b3f946)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32e46135)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fab4aa5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_253) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f948134)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_125) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(104d3db0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fab4aa5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce022162)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d810586d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0e2b021)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a4c1697)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17e259db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28f58f60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28f24e70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_110) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_255) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c817084d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ce0f04b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_271 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_277 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_247) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ead8b2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9990aef4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_250) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17b669c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f52b81f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_110) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ddb184e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96c58310)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1ac0a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_56 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_62 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_64 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_69 = _RAND_3[0:0];
  _RAND_4 = {18{`RANDOM}};
  _EVAL_78 = _RAND_4[575:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_87 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_96 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_107 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_122 = _RAND_8[29:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_128 = _RAND_9[9:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_137 = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_145 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_175 = _RAND_12[9:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_190 = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_193 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_208 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_211 = _RAND_16[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
