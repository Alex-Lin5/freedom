//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_151_assert(
  input  [1:0]  _EVAL,
  input  [3:0]  _EVAL_0,
  input  [2:0]  _EVAL_1,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [9:0]  _EVAL_7,
  input  [25:0] _EVAL_11,
  input         _EVAL_13,
  input  [2:0]  _EVAL_14,
  input         _EVAL_18,
  input         _EVAL_19,
  input         _EVAL_31,
  input         _EVAL_36,
  input         _EVAL_40,
  input         _EVAL_42,
  input         _EVAL_50,
  input         _EVAL_55,
  input         _EVAL_57,
  input  [7:0]  _EVAL_70,
  input         _EVAL_75,
  input         _EVAL_80,
  input         _EVAL_83,
  input  [7:0]  _EVAL_99,
  input         _EVAL_102,
  input         _EVAL_107,
  input  [31:0] _EVAL_115,
  input         _EVAL_117,
  input  [7:0]  _EVAL_123,
  input         _EVAL_131,
  input  [7:0]  _EVAL_138,
  input         _EVAL_139,
  input         _EVAL_145,
  input         _EVAL_147,
  input         _EVAL_150,
  input         _EVAL_160,
  input         _EVAL_163,
  input         _EVAL_164,
  input         _EVAL_169,
  input         _EVAL_178,
  input         _EVAL_181,
  input         _EVAL_191,
  input         _EVAL_196,
  input         _EVAL_198
);
  wire  _EVAL_22;
  wire  _EVAL_24;
  wire  _EVAL_29;
  wire  _EVAL_32;
  wire  _EVAL_43;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_61;
  wire  _EVAL_65;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_73;
  wire  _EVAL_82;
  wire  _EVAL_84;
  wire  _EVAL_87;
  wire  _EVAL_90;
  wire  _EVAL_95;
  wire  _EVAL_100;
  wire  _EVAL_112;
  wire  monitor__EVAL;
  wire [1:0] monitor__EVAL_0;
  wire [9:0] monitor__EVAL_1;
  wire [2:0] monitor__EVAL_2;
  wire  monitor__EVAL_3;
  wire [25:0] monitor__EVAL_4;
  wire [2:0] monitor__EVAL_5;
  wire  monitor__EVAL_6;
  wire  monitor__EVAL_7;
  wire  monitor__EVAL_8;
  wire [9:0] monitor__EVAL_9;
  wire  monitor__EVAL_10;
  wire [3:0] monitor__EVAL_11;
  wire [2:0] monitor__EVAL_12;
  wire [1:0] monitor__EVAL_13;
  wire  monitor__EVAL_14;
  wire  _EVAL_116;
  wire  _EVAL_120;
  wire  _EVAL_126;
  wire  _EVAL_133;
  wire  _EVAL_140;
  wire  _EVAL_148;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_159;
  wire [30:0] _EVAL_165;
  wire  _EVAL_170;
  wire  _EVAL_173;
  wire  _EVAL_176;
  wire  _EVAL_182;
  wire  _EVAL_184;
  wire  _EVAL_188;
  wire  _EVAL_194;
  wire  _EVAL_201;
  _EVAL_150_assert monitor (
    ._EVAL(monitor__EVAL),
    ._EVAL_0(monitor__EVAL_0),
    ._EVAL_1(monitor__EVAL_1),
    ._EVAL_2(monitor__EVAL_2),
    ._EVAL_3(monitor__EVAL_3),
    ._EVAL_4(monitor__EVAL_4),
    ._EVAL_5(monitor__EVAL_5),
    ._EVAL_6(monitor__EVAL_6),
    ._EVAL_7(monitor__EVAL_7),
    ._EVAL_8(monitor__EVAL_8),
    ._EVAL_9(monitor__EVAL_9),
    ._EVAL_10(monitor__EVAL_10),
    ._EVAL_11(monitor__EVAL_11),
    ._EVAL_12(monitor__EVAL_12),
    ._EVAL_13(monitor__EVAL_13),
    ._EVAL_14(monitor__EVAL_14)
  );
  assign _EVAL_90 = _EVAL_140 & _EVAL_126;
  assign _EVAL_112 = _EVAL_140 & _EVAL_95;
  assign monitor__EVAL_5 = _EVAL_1;
  assign _EVAL_61 = _EVAL_148 & _EVAL_95;
  assign _EVAL_73 = _EVAL_53 & _EVAL_50;
  assign _EVAL_194 = _EVAL_155 & _EVAL_69;
  assign _EVAL_133 = _EVAL_155 & _EVAL_188;
  assign _EVAL_173 = _EVAL_53 & _EVAL_55;
  assign _EVAL_116 = _EVAL_54 & _EVAL_126;
  assign _EVAL_43 = _EVAL_54 & _EVAL_95;
  assign _EVAL_95 = |_EVAL_70;
  assign _EVAL_148 = _EVAL_120 & _EVAL_191;
  assign _EVAL_120 = _EVAL_53 & _EVAL_196;
  assign _EVAL_65 = _EVAL_53 & _EVAL_169;
  assign _EVAL_53 = _EVAL_42 & _EVAL_83;
  assign _EVAL_84 = _EVAL_154 & _EVAL_126;
  assign _EVAL_126 = |_EVAL_123;
  assign _EVAL_32 = _EVAL_148 & _EVAL_126;
  assign _EVAL_154 = _EVAL_68 & _EVAL_191;
  assign monitor__EVAL_11 = _EVAL_0;
  assign _EVAL_24 = _EVAL_154 & _EVAL_100;
  assign monitor__EVAL_6 = _EVAL_6;
  assign _EVAL_82 = _EVAL_140 & _EVAL_201;
  assign _EVAL_176 = _EVAL_140 & _EVAL_100;
  assign monitor__EVAL_9 = _EVAL_7;
  assign monitor__EVAL_2 = {{2'd0}, _EVAL_83};
  assign _EVAL_54 = _EVAL_65 & _EVAL_147;
  assign _EVAL_155 = _EVAL_73 & _EVAL_147;
  assign _EVAL_87 = _EVAL_148 & _EVAL_201;
  assign _EVAL_69 = |_EVAL_145;
  assign monitor__EVAL_8 = _EVAL_19;
  assign monitor__EVAL_13 = _EVAL;
  assign monitor__EVAL_10 = _EVAL_19;
  assign monitor__EVAL_14 = _EVAL_18;
  assign _EVAL_170 = _EVAL_154 & _EVAL_201;
  assign _EVAL_159 = _EVAL_54 & _EVAL_201;
  assign monitor__EVAL_0 = _EVAL;
  assign monitor__EVAL_4 = _EVAL_11;
  assign _EVAL_100 = |_EVAL_138;
  assign _EVAL_184 = _EVAL_154 & _EVAL_95;
  assign _EVAL_140 = _EVAL_173 & _EVAL_147;
  assign _EVAL_182 = _EVAL_148 & _EVAL_100;
  assign monitor__EVAL_1 = _EVAL_7;
  assign monitor__EVAL_3 = _EVAL_13;
  assign _EVAL_165 = _EVAL_115[31:1];
  assign _EVAL_22 = ~_EVAL_18;
  assign monitor__EVAL = _EVAL_5;
  assign _EVAL_188 = |_EVAL_165;
  assign _EVAL_68 = _EVAL_53 & _EVAL_163;
  assign monitor__EVAL_12 = _EVAL_14;
  assign _EVAL_201 = |_EVAL_99;
  assign _EVAL_29 = _EVAL_54 & _EVAL_100;
  assign monitor__EVAL_7 = _EVAL_6;
  always @(posedge _EVAL_13) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d728da28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a93fa1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0ccaf87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4bb50746)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1e2b9de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a066dad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_87 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(892a9b02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84e08e5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_160 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c76ebb8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1b1984c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b68130b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c642a68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efffd529)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba8a47cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e8de179)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac31dbf3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84f58be9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44ae3a00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(920a5bc3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6aae87f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9c8527c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8659adfd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f92651f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7681f14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ddb81638)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b112b89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95eca6d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c7743c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a0330cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d84d4652)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e505de33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(345372dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8766607)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24e71c4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c578052)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7381506f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(416aa22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_84 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(909a4a55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(654354f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_150 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9826ea9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22693138)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9e4ad4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a42f00b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8e1b6fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d63a1b53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_131 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(295d3f37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd99d295)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67dfa2bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(265f29f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18d118e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9412e4e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72950ec8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea06257a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(359a9d36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_24 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8f3414e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6b501c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a16c6f8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20398d6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f951af43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfdeba96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4fee2156)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_57 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90930b85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52c12412)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa9065f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee1668a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(725b18e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_164 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bd80af0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce39add9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be8f674c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_116 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e09d4cec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
