//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_114(
  output [31:0] _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  output        _EVAL_2,
  output [31:0] _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [1:0]  _EVAL_7,
  input  [1:0]  _EVAL_8,
  input  [31:0] _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input  [31:0] _EVAL_13,
  input         _EVAL_14,
  input  [31:0] _EVAL_15,
  output [7:0]  _EVAL_16,
  input         _EVAL_17,
  output [4:0]  _EVAL_18,
  output        _EVAL_19,
  input         _EVAL_20,
  input  [31:0] _EVAL_21,
  output        _EVAL_22,
  output        _EVAL_23,
  input  [4:0]  _EVAL_24,
  input  [7:0]  _EVAL_25,
  input         _EVAL_26,
  input  [31:0] _EVAL_27,
  output        _EVAL_28
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_120;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
`endif // RANDOMIZE_REG_INIT
  reg [12:0] _EVAL_29;
  wire  _EVAL_30;
  reg  _EVAL_31;
  reg [12:0] _EVAL_32;
  wire [13:0] _EVAL_33;
  wire [3:0] _EVAL_34;
  reg [12:0] _EVAL_35;
  wire  _EVAL_36;
  reg [12:0] _EVAL_37;
  reg  _EVAL_38;
  wire  _EVAL_39;
  wire [2:0] _EVAL_40;
  wire [17:0] _EVAL_41;
  wire [2:0] _EVAL_42;
  reg [2:0] _EVAL_43;
  wire  _EVAL_44;
  reg [1:0] _EVAL_45;
  reg [2:0] _EVAL_46;
  wire [12:0] _EVAL_48;
  reg [31:0] _EVAL_50;
  wire  _EVAL_52;
  wire [6:0] _EVAL_54;
  wire [2:0] _EVAL_55;
  wire [26:0] _EVAL_56;
  wire  _EVAL_57;
  wire [8:0] _EVAL_58;
  wire  _EVAL_59;
  wire [7:0] _EVAL_61;
  wire  _EVAL_62;
  reg  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  reg  _EVAL_72;
  reg [1:0] _EVAL_73;
  reg [2:0] _EVAL_76;
  wire  _EVAL_77;
  wire [9:0] _EVAL_79;
  wire [2:0] _EVAL_80;
  reg [1:0] _EVAL_82;
  wire [2:0] _EVAL_83;
  wire  _EVAL_84;
  reg  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire [17:0] _EVAL_89;
  wire [27:0] _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire [7:0] _EVAL_95;
  reg [2:0] _EVAL_97;
  wire  _EVAL_98;
  reg [12:0] _EVAL_99;
  wire  _EVAL_100;
  wire [2:0] _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  reg  _EVAL_104;
  wire  _EVAL_106;
  reg [12:0] _EVAL_107;
  wire  _EVAL_108;
  wire [2:0] _EVAL_109;
  wire [7:0] _EVAL_110;
  wire [6:0] _EVAL_112;
  wire [2:0] _EVAL_114;
  wire [1:0] _EVAL_115;
  wire [2:0] _EVAL_116;
  wire  _EVAL_118;
  wire [12:0] _EVAL_119;
  wire [2:0] _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  reg [12:0] _EVAL_123;
  wire  _EVAL_125;
  reg [2:0] _EVAL_127;
  wire [2:0] _EVAL_128;
  reg  _EVAL_129;
  wire [2:0] _EVAL_130;
  reg [9:0] _EVAL_131;
  wire  _EVAL_132;
  reg [1:0] _EVAL_133;
  wire [2:0] _EVAL_134;
  reg [1:0] _EVAL_135;
  wire [1:0] _EVAL_136;
  wire  _EVAL_137;
  wire [3:0] _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire [2:0] _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire [7:0] _EVAL_149;
  wire [2:0] _EVAL_150;
  reg [12:0] _EVAL_151;
  wire  _EVAL_152;
  wire [2:0] _EVAL_153;
  reg [12:0] _EVAL_155;
  wire [12:0] _EVAL_156;
  wire [12:0] _EVAL_157;
  wire [2:0] _EVAL_158;
  reg [12:0] _EVAL_159;
  wire [1:0] _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire [2:0] _EVAL_166;
  wire  _EVAL_167;
  wire [7:0] _EVAL_168;
  wire [1:0] _EVAL_170;
  reg [2:0] _EVAL_171;
  reg [2:0] _EVAL_172;
  reg [2:0] _EVAL_173;
  reg [1:0] _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire [12:0] _EVAL_177;
  wire [2:0] _EVAL_178;
  wire [31:0] _EVAL_179;
  wire [3:0] _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire [2:0] _EVAL_186;
  wire  _EVAL_187;
  wire [2:0] _EVAL_189;
  wire  _EVAL_190;
  wire [2:0] _EVAL_193;
  reg [17:0] _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  reg [12:0] _EVAL_199;
  wire [12:0] _EVAL_201;
  wire [12:0] _EVAL_202;
  wire [2:0] _EVAL_203;
  reg [31:0] _EVAL_204;
  wire [7:0] _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  reg [12:0] _EVAL_209;
  wire  _EVAL_210;
  wire [12:0] _EVAL_211;
  wire [2:0] _EVAL_212;
  reg [12:0] _EVAL_213;
  wire [12:0] _EVAL_215;
  wire [31:0] _EVAL_216;
  wire  _EVAL_217;
  wire [12:0] _EVAL_218;
  wire  _EVAL_219;
  wire [17:0] _EVAL_222;
  reg [2:0] _EVAL_223;
  wire [17:0] _EVAL_224;
  wire  _EVAL_226;
  wire [2:0] _EVAL_228;
  wire [2:0] _EVAL_229;
  wire  _EVAL_230;
  reg [2:0] _EVAL_231;
  wire [6:0] _EVAL_232;
  reg [1:0] _EVAL_233;
  wire [8:0] _EVAL_234;
  wire  _EVAL_236;
  wire [12:0] _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire [1:0] _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire [1:0] _EVAL_248;
  wire [2:0] _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_253;
  wire [31:0] _EVAL_254;
  wire  _EVAL_256;
  wire [2:0] _EVAL_257;
  wire  _EVAL_258;
  wire [6:0] _EVAL_259;
  wire  _EVAL_260;
  wire [2:0] _EVAL_261;
  wire [2:0] _EVAL_262;
  wire [31:0] _EVAL_263;
  wire  _EVAL_264;
  wire [6:0] _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire [27:0] _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire [2:0] _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_278;
  reg [1:0] _EVAL_279;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire [1:0] _EVAL_283;
  wire  _EVAL_284;
  reg [12:0] _EVAL_285;
  reg [12:0] _EVAL_286;
  reg [31:0] _EVAL_287;
  wire [2:0] _EVAL_289;
  wire [10:0] _EVAL_291;
  wire [6:0] _EVAL_293;
  reg [12:0] _EVAL_294;
  reg [12:0] _EVAL_295;
  wire  _EVAL_296;
  wire [2:0] _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_300;
  reg  _EVAL_301;
  wire  _EVAL_304;
  reg [2:0] _EVAL_305;
  wire [17:0] _EVAL_306;
  wire [27:0] _EVAL_307;
  wire [2:0] _EVAL_310;
  wire [8:0] _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_314;
  wire [12:0] _EVAL_316;
  wire  _EVAL_317;
  wire [12:0] _EVAL_318;
  wire [2:0] _EVAL_319;
  reg [2:0] _EVAL_321;
  wire  _EVAL_322;
  reg [1:0] _EVAL_323;
  wire [3:0] _EVAL_324;
  wire [20:0] _EVAL_326;
  wire [12:0] _EVAL_327;
  reg [12:0] _EVAL_328;
  wire [27:0] _EVAL_329;
  wire  _EVAL_330;
  wire [7:0] _EVAL_331;
  wire [2:0] _EVAL_333;
  wire  _EVAL_334;
  wire  _EVAL_336;
  wire  _EVAL_337;
  wire [2:0] _EVAL_338;
  reg [31:0] _EVAL_339;
  reg [2:0] _EVAL_341;
  wire  _EVAL_342;
  wire  _EVAL_344;
  reg [1:0] _EVAL_345;
  reg [5:0] _EVAL_347;
  reg [2:0] _EVAL_348;
  wire [14:0] _EVAL_349;
  wire  _EVAL_350;
  wire  _EVAL_351;
  wire  _EVAL_352;
  wire [2:0] _EVAL_355;
  reg [12:0] _EVAL_356;
  wire  _EVAL_357;
  wire [27:0] _EVAL_359;
  wire [2:0] _EVAL_360;
  wire  _EVAL_361;
  wire [12:0] _EVAL_362;
  wire [2:0] _EVAL_364;
  wire [3:0] _EVAL_365;
  wire [31:0] _EVAL_366;
  wire  _EVAL_367;
  wire  _EVAL_368;
  wire  _EVAL_369;
  wire [2:0] _EVAL_370;
  wire [12:0] _EVAL_371;
  wire  _EVAL_372;
  wire  _EVAL_373;
  wire  _EVAL_374;
  wire [17:0] _EVAL_375;
  wire [31:0] _EVAL_377;
  reg [12:0] _EVAL_378;
  wire [5:0] _EVAL_379;
  wire  _EVAL_380;
  wire  _EVAL_381;
  wire  _EVAL_382;
  wire  _EVAL_384;
  wire  _EVAL_385;
  wire [2:0] _EVAL_386;
  reg [12:0] _EVAL_387;
  wire [2:0] _EVAL_388;
  wire [6:0] _EVAL_389;
  wire [12:0] _EVAL_390;
  wire  _EVAL_391;
  wire [12:0] _EVAL_393;
  reg  _EVAL_394;
  wire [2:0] _EVAL_395;
  wire  _EVAL_396;
  wire  _EVAL_397;
  wire [6:0] _EVAL_398;
  wire [2:0] _EVAL_399;
  wire [4:0] _EVAL_400;
  reg [2:0] _EVAL_401;
  wire [17:0] _EVAL_402;
  wire [3:0] _EVAL_403;
  wire  _EVAL_405;
  reg [12:0] _EVAL_406;
  wire  _EVAL_407;
  wire [29:0] _EVAL_408;
  wire [1:0] _EVAL_409;
  wire  _EVAL_410;
  wire [7:0] _EVAL_411;
  wire [13:0] _EVAL_412;
  wire  _EVAL_413;
  reg [2:0] _EVAL_414;
  reg  _EVAL_415;
  wire [12:0] _EVAL_416;
  wire [1:0] _EVAL_417;
  wire  _EVAL_418;
  wire  _EVAL_419;
  wire [1:0] _EVAL_420;
  wire [2:0] _EVAL_422;
  wire [12:0] _EVAL_425;
  wire [15:0] _EVAL_426;
  wire  _EVAL_427;
  wire  _EVAL_432;
  wire [3:0] _EVAL_433;
  wire [2:0] _EVAL_436;
  wire  _EVAL_437;
  wire  _EVAL_439;
  wire [6:0] _EVAL_440;
  wire  _EVAL_442;
  wire [2:0] _EVAL_444;
  wire [2:0] _EVAL_445;
  wire [6:0] _EVAL_446;
  wire [27:0] _EVAL_448;
  wire  _EVAL_449;
  wire  _EVAL_451;
  reg [2:0] _EVAL_452;
  wire  _EVAL_453;
  wire [6:0] _EVAL_454;
  wire  _EVAL_455;
  reg [2:0] _EVAL_456;
  wire [6:0] _EVAL_458;
  wire [2:0] _EVAL_459;
  wire [2:0] _EVAL_460;
  wire  _EVAL_461;
  wire [1:0] _EVAL_464;
  reg [2:0] _EVAL_465;
  wire [7:0] _EVAL_466;
  reg [1:0] _EVAL_467;
  wire  _EVAL_468;
  wire [1:0] _EVAL_469;
  wire  _EVAL_470;
  wire  _EVAL_471;
  wire  _EVAL_472;
  wire  _EVAL_473;
  reg  _EVAL_474;
  wire [2:0] _EVAL_475;
  wire [12:0] _EVAL_476;
  wire  _EVAL_477;
  wire [31:0] _EVAL_478;
  reg [12:0] _EVAL_479;
  wire [2:0] _EVAL_480;
  reg [1:0] _EVAL_481;
  wire [12:0] _EVAL_482;
  wire [2:0] _EVAL_483;
  wire  _EVAL_484;
  wire  _EVAL_485;
  reg [1:0] _EVAL_486;
  reg  _EVAL_487;
  reg [1:0] _EVAL_488;
  wire  _EVAL_489;
  wire [2:0] _EVAL_490;
  wire  _EVAL_494;
  reg [12:0] _EVAL_495;
  wire [2:0] _EVAL_496;
  wire  _EVAL_497;
  wire  _EVAL_498;
  wire  _EVAL_499;
  wire [2:0] _EVAL_500;
  wire  _EVAL_501;
  wire  _EVAL_502;
  wire [12:0] _EVAL_503;
  wire [2:0] _EVAL_504;
  wire [27:0] _EVAL_505;
  wire  _EVAL_506;
  reg [12:0] _EVAL_507;
  wire [2:0] _EVAL_508;
  wire  _EVAL_509;
  reg [17:0] _EVAL_510;
  wire  _EVAL_511;
  wire  _EVAL_512;
  wire  _EVAL_513;
  reg [12:0] _EVAL_515;
  wire  _EVAL_516;
  reg [12:0] _EVAL_517;
  wire [12:0] _EVAL_519;
  wire  _EVAL_520;
  wire  _EVAL_522;
  wire [2:0] _EVAL_523;
  wire [2:0] _EVAL_524;
  wire  _EVAL_525;
  wire [2:0] _EVAL_526;
  wire [2:0] _EVAL_527;
  wire  _EVAL_528;
  wire [3:0] _EVAL_529;
  wire  _EVAL_530;
  wire  _EVAL_531;
  wire [2:0] _EVAL_532;
  wire  _EVAL_533;
  wire  _EVAL_534;
  wire [7:0] _EVAL_535;
  reg [31:0] _EVAL_536;
  reg [12:0] _EVAL_537;
  wire  _EVAL_538;
  wire  _EVAL_539;
  wire  _EVAL_540;
  wire  _EVAL_541;
  wire [3:0] _EVAL_542;
  wire  _EVAL_543;
  wire [1:0] _EVAL_544;
  wire [6:0] _EVAL_545;
  wire  _EVAL_546;
  wire [1:0] _EVAL_547;
  wire  _EVAL_548;
  reg  _EVAL_549;
  wire  _EVAL_550;
  reg [1:0] _EVAL_551;
  wire [12:0] _EVAL_552;
  reg [12:0] _EVAL_553;
  wire [5:0] _EVAL_554;
  wire  _EVAL_556;
  wire  _EVAL_557;
  wire [2:0] _EVAL_558;
  wire  _EVAL_559;
  reg [12:0] _EVAL_560;
  wire [2:0] _EVAL_561;
  wire  _EVAL_562;
  wire  _EVAL_563;
  wire  _EVAL_564;
  wire  _EVAL_565;
  wire [12:0] _EVAL_566;
  wire [8:0] _EVAL_567;
  wire  _EVAL_568;
  reg  _EVAL_569;
  wire [11:0] _EVAL_570;
  wire [3:0] _EVAL_571;
  wire [15:0] _EVAL_572;
  wire  _EVAL_573;
  wire [12:0] _EVAL_574;
  wire  _EVAL_575;
  reg [12:0] _EVAL_576;
  wire [12:0] _EVAL_577;
  wire  _EVAL_578;
  wire  _EVAL_579;
  wire [7:0] _EVAL_580;
  wire  _EVAL_581;
  wire  _EVAL_582;
  wire  _EVAL_583;
  wire [3:0] _EVAL_584;
  wire [2:0] _EVAL_585;
  reg [17:0] _EVAL_586;
  wire [1:0] _EVAL_587;
  wire [2:0] _EVAL_588;
  wire [2:0] _EVAL_589;
  wire  _EVAL_590;
  wire  _EVAL_592;
  reg [2:0] _EVAL_593;
  wire  _EVAL_594;
  reg  _EVAL_595;
  wire  _EVAL_598;
  wire [31:0] _EVAL_599;
  wire [1:0] _EVAL_600;
  wire  _EVAL_601;
  wire  _EVAL_602;
  wire [2:0] _EVAL_603;
  wire [2:0] _EVAL_604;
  wire  _EVAL_605;
  wire [8:0] _EVAL_606;
  wire  _EVAL_607;
  wire [7:0] _EVAL_609;
  wire [2:0] _EVAL_610;
  wire [2:0] _EVAL_612;
  wire  _EVAL_613;
  wire  _EVAL_614;
  wire [7:0] _EVAL_617;
  reg [2:0] _EVAL_619;
  wire [12:0] _EVAL_620;
  wire [17:0] _EVAL_621;
  reg  _EVAL_622;
  wire [10:0] _EVAL_624;
  wire [2:0] _EVAL_625;
  wire  _EVAL_626;
  reg [2:0] _EVAL_627;
  reg [12:0] _EVAL_628;
  wire  _EVAL_631;
  wire  _EVAL_632;
  reg  _EVAL_633;
  reg [31:0] _EVAL_634;
  wire [3:0] _EVAL_635;
  reg [2:0] _EVAL_636;
  wire  _EVAL_638;
  wire  _EVAL_639;
  wire [2:0] _EVAL_640;
  wire [1:0] _EVAL_641;
  reg [12:0] _EVAL_642;
  wire  _EVAL_643;
  wire  _EVAL_644;
  wire  _EVAL_645;
  wire [2:0] _EVAL_649;
  wire [2:0] _EVAL_651;
  wire  _EVAL_652;
  wire  _EVAL_653;
  wire  _EVAL_654;
  wire  _EVAL_657;
  wire  _EVAL_658;
  wire  _EVAL_660;
  wire [1:0] _EVAL_661;
  wire  _EVAL_662;
  wire  _EVAL_663;
  reg [2:0] _EVAL_664;
  reg [2:0] _EVAL_665;
  wire  _EVAL_667;
  wire [3:0] _EVAL_668;
  wire  _EVAL_670;
  wire  _EVAL_671;
  wire [27:0] _EVAL_672;
  reg [1:0] _EVAL_673;
  wire [17:0] _EVAL_674;
  wire  _EVAL_675;
  reg [12:0] _EVAL_676;
  wire  _EVAL_677;
  wire  _EVAL_678;
  reg [12:0] _EVAL_679;
  wire  _EVAL_680;
  wire  _EVAL_681;
  wire  _EVAL_682;
  wire  _EVAL_683;
  wire  _EVAL_684;
  wire [14:0] _EVAL_685;
  wire  _EVAL_686;
  wire [2:0] _EVAL_688;
  reg  _EVAL_689;
  wire [2:0] _EVAL_690;
  wire  _EVAL_691;
  wire [2:0] _EVAL_692;
  wire  _EVAL_694;
  wire  _EVAL_695;
  wire  _EVAL_696;
  wire [7:0] _EVAL_697;
  wire [2:0] _EVAL_698;
  wire [12:0] _EVAL_700;
  wire [2:0] _EVAL_701;
  reg [1:0] _EVAL_703;
  wire [3:0] _EVAL_704;
  wire [1:0] _EVAL_706;
  wire  _EVAL_707;
  wire [13:0] _EVAL_708;
  wire  _EVAL_709;
  wire [9:0] _EVAL_710;
  wire  _EVAL_711;
  wire [2:0] _EVAL_712;
  wire  _EVAL_714;
  reg [2:0] _EVAL_715;
  wire [2:0] _EVAL_717;
  wire  _EVAL_718;
  reg [2:0] _EVAL_719;
  wire  _EVAL_720;
  wire  _EVAL_721;
  wire  _EVAL_722;
  wire  _EVAL_723;
  wire  _EVAL_724;
  wire  _EVAL_725;
  reg [12:0] _EVAL_726;
  reg [2:0] _EVAL_729;
  reg [12:0] _EVAL_730;
  wire  _EVAL_731;
  wire [2:0] _EVAL_732;
  wire [3:0] _EVAL_733;
  wire [2:0] _EVAL_734;
  wire [1:0] _EVAL_735;
  wire  _EVAL_736;
  wire  _EVAL_737;
  wire  _EVAL_738;
  wire  _EVAL_740;
  reg [12:0] _EVAL_741;
  wire  _EVAL_743;
  wire [1:0] _EVAL_744;
  wire [4:0] _EVAL_745;
  wire [12:0] _EVAL_746;
  wire [5:0] _EVAL_747;
  wire [6:0] _EVAL_748;
  wire [15:0] _EVAL_750;
  wire  _EVAL_751;
  wire  _EVAL_752;
  reg [12:0] _EVAL_753;
  wire [12:0] _EVAL_754;
  wire  _EVAL_756;
  wire [2:0] _EVAL_757;
  wire  _EVAL_758;
  reg  _EVAL_759;
  wire  _EVAL_760;
  wire  _EVAL_762;
  wire [7:0] _EVAL_763;
  wire  _EVAL_764;
  wire [15:0] _EVAL_765;
  wire  _EVAL_766;
  wire  _EVAL_767;
  wire [2:0] _EVAL_768;
  reg [1:0] _EVAL_769;
  wire [1:0] _EVAL_770;
  wire [3:0] _EVAL_771;
  wire  _EVAL_772;
  wire [2:0] _EVAL_773;
  wire [12:0] _EVAL_774;
  wire [1:0] _EVAL_775;
  wire [2:0] _EVAL_776;
  wire [2:0] _EVAL_777;
  wire  _EVAL_778;
  reg [12:0] _EVAL_779;
  wire [2:0] _EVAL_780;
  wire  _EVAL_782;
  wire [2:0] _EVAL_783;
  reg  _EVAL_784;
  wire [6:0] _EVAL_785;
  wire  _EVAL_786;
  wire [3:0] _EVAL_787;
  wire [7:0] _EVAL_788;
  wire [12:0] _EVAL_789;
  wire  _EVAL_790;
  reg [2:0] _EVAL_791;
  wire  _EVAL_792;
  wire [12:0] _EVAL_793;
  reg [7:0] _EVAL_794;
  wire [6:0] _EVAL_795;
  wire  _EVAL_796;
  wire [3:0] _EVAL_797;
  wire [1:0] _EVAL_798;
  wire [8:0] _EVAL_799;
  wire  _EVAL_800;
  wire  _EVAL_801;
  wire [2:0] _EVAL_803;
  reg [12:0] _EVAL_804;
  wire  _EVAL_805;
  wire [2:0] _EVAL_806;
  wire [1:0] _EVAL_807;
  reg  _EVAL_808 [0:511];
  wire  _EVAL_808__EVAL_809_data;
  wire [8:0] _EVAL_808__EVAL_809_addr;
  wire  _EVAL_808__EVAL_810_data;
  wire [8:0] _EVAL_808__EVAL_810_addr;
  wire  _EVAL_808__EVAL_810_mask;
  wire  _EVAL_808__EVAL_810_en;
  reg  _EVAL_811;
  wire  _EVAL_812;
  wire [31:0] _EVAL_813;
  wire [3:0] _EVAL_814;
  wire  _EVAL_815;
  reg [2:0] _EVAL_816;
  wire [2:0] _EVAL_818;
  reg [12:0] _EVAL_819;
  wire  _EVAL_820;
  wire  _EVAL_821;
  reg [2:0] _EVAL_823;
  reg [1:0] _EVAL_824;
  reg [2:0] _EVAL_825;
  reg [2:0] _EVAL_826;
  wire  _EVAL_827;
  wire [1:0] _EVAL_829;
  wire [7:0] _EVAL_830;
  reg [2:0] _EVAL_831;
  wire [1:0] _EVAL_832;
  reg  _EVAL_833;
  reg [1:0] _EVAL_835;
  wire [2:0] _EVAL_836;
  wire  _EVAL_838;
  wire [12:0] _EVAL_840;
  reg [1:0] _EVAL_842;
  reg  _EVAL_843;
  wire  _EVAL_845;
  wire [2:0] _EVAL_847;
  reg [12:0] _EVAL_848;
  wire [3:0] _EVAL_849;
  wire [12:0] _EVAL_850;
  wire  _EVAL_851;
  wire [2:0] _EVAL_852;
  reg [26:0] _EVAL_853;
  wire [2:0] _EVAL_855;
  wire [12:0] _EVAL_856;
  reg [2:0] _EVAL_857;
  wire  _EVAL_858;
  wire  _EVAL_859;
  wire  _EVAL_860;
  wire  _EVAL_862;
  wire [2:0] _EVAL_864;
  wire  _EVAL_865;
  wire  _EVAL_866;
  wire  _EVAL_867;
  wire [14:0] _EVAL_868;
  wire [2:0] _EVAL_869;
  wire  _EVAL_870;
  wire [2:0] _EVAL_872;
  wire  _EVAL_873;
  wire  _EVAL_874;
  wire [2:0] _EVAL_875;
  wire [17:0] _EVAL_876;
  wire  _EVAL_877;
  wire [2:0] _EVAL_878;
  wire [1:0] _EVAL_879;
  wire [10:0] _EVAL_882;
  wire  _EVAL_884;
  wire  _EVAL_885;
  reg [2:0] _EVAL_886;
  wire  _EVAL_887;
  wire [2:0] _EVAL_888;
  wire [2:0] _EVAL_889;
  wire [2:0] _EVAL_890;
  reg [2:0] _EVAL_891;
  wire [2:0] _EVAL_893;
  wire [20:0] _EVAL_895;
  wire  _EVAL_896;
  wire  _EVAL_897;
  wire [2:0] _EVAL_899;
  wire [17:0] _EVAL_900;
  wire [3:0] _EVAL_901;
  wire  _EVAL_902;
  wire  _EVAL_903;
  wire [2:0] _EVAL_904;
  wire  _EVAL_905;
  wire  _EVAL_906;
  wire [10:0] _EVAL_907;
  wire [12:0] _EVAL_908;
  wire [2:0] _EVAL_909;
  wire [2:0] _EVAL_911;
  wire  _EVAL_912;
  wire [2:0] _EVAL_913;
  wire  _EVAL_914;
  wire  _EVAL_916;
  wire [17:0] _EVAL_917;
  reg [1:0] _EVAL_918;
  reg [2:0] _EVAL_919;
  wire  _EVAL_920;
  reg [27:0] _EVAL_921;
  wire  _EVAL_922;
  wire [12:0] _EVAL_923;
  wire [2:0] _EVAL_925;
  wire  _EVAL_926;
  wire  _EVAL_927;
  wire  _EVAL_928;
  wire  _EVAL_929;
  reg [2:0] _EVAL_930;
  wire  _EVAL_931;
  wire [12:0] _EVAL_932;
  wire [1:0] _EVAL_934;
  wire  _EVAL_935;
  wire  _EVAL_936;
  wire  _EVAL_937;
  wire  _EVAL_939;
  wire  _EVAL_940;
  wire  _EVAL_941;
  wire [31:0] _EVAL_943;
  wire [2:0] _EVAL_944;
  wire [6:0] _EVAL_945;
  reg [4:0] _EVAL_946;
  wire  _EVAL_947;
  wire  _EVAL_948;
  wire  _EVAL_949;
  wire [6:0] _EVAL_950;
  reg [12:0] _EVAL_951;
  reg [2:0] _EVAL_952;
  reg [12:0] _EVAL_954;
  reg [2:0] _EVAL_955;
  wire  _EVAL_956;
  wire  _EVAL_957;
  wire  _EVAL_958;
  wire  _EVAL_959;
  reg  _EVAL_960;
  wire [12:0] _EVAL_961;
  wire  _EVAL_962;
  wire  _EVAL_963;
  wire  _EVAL_966;
  wire [7:0] _EVAL_967;
  wire  _EVAL_968;
  wire [5:0] _EVAL_969;
  wire [2:0] _EVAL_970;
  reg [2:0] _EVAL_971;
  reg  _EVAL_972;
  reg [2:0] _EVAL_973;
  wire [12:0] _EVAL_974;
  reg [2:0] _EVAL_976;
  wire  _EVAL_977;
  reg [4:0] _EVAL_978;
  wire [9:0] _EVAL_979;
  wire  _EVAL_982;
  wire  _EVAL_983;
  wire [3:0] _EVAL_984;
  wire [2:0] _EVAL_985;
  wire [2:0] _EVAL_986;
  wire [30:0] _EVAL_987;
  wire  _EVAL_988;
  wire  _EVAL_989;
  reg  _EVAL_990;
  wire  _EVAL_991;
  wire  _EVAL_992;
  reg [12:0] _EVAL_993;
  wire [17:0] _EVAL_994;
  wire  _EVAL_995;
  wire  _EVAL_996;
  wire  _EVAL_997;
  wire [6:0] _EVAL_998;
  wire [7:0] _EVAL_1000;
  wire  _EVAL_1003;
  wire  _EVAL_1004;
  wire  _EVAL_1005;
  reg  _EVAL_1006;
  reg [12:0] _EVAL_1007;
  wire  _EVAL_1008;
  wire [1:0] _EVAL_1009;
  reg [1:0] _EVAL_1010;
  wire [12:0] _EVAL_1011;
  reg [2:0] _EVAL_1012;
  wire [7:0] _EVAL_1013;
  wire  _EVAL_1014;
  reg  _EVAL_1016;
  wire  _EVAL_1018;
  wire [2:0] _EVAL_1020;
  wire  _EVAL_1021;
  wire [7:0] _EVAL_1022;
  wire [2:0] _EVAL_1024;
  wire  _EVAL_1025;
  reg [31:0] _EVAL_1026;
  wire [6:0] _EVAL_1027;
  wire  _EVAL_1028;
  reg [12:0] _EVAL_1030;
  wire  _EVAL_1031;
  wire  _EVAL_1032;
  wire [1:0] _EVAL_1033;
  wire  _EVAL_1034;
  wire [2:0] _EVAL_1035;
  wire [31:0] _EVAL_1036;
  wire [2:0] _EVAL_1037;
  wire [2:0] _EVAL_1038;
  wire  _EVAL_1039;
  wire [12:0] _EVAL_1040;
  wire [2:0] _EVAL_1041;
  wire [13:0] _EVAL_1042;
  wire [2:0] _EVAL_1043;
  wire  _EVAL_1044;
  wire  _EVAL_1045;
  reg [12:0] _EVAL_1048;
  wire [2:0] _EVAL_1049;
  wire  _EVAL_1050;
  wire  _EVAL_1051;
  wire [5:0] _EVAL_1052;
  wire [12:0] _EVAL_1053;
  reg [2:0] _EVAL_1054;
  reg [1:0] _EVAL_1055;
  reg [12:0] _EVAL_1057;
  wire [7:0] _EVAL_1058;
  wire [12:0] _EVAL_1059;
  wire [2:0] _EVAL_1060;
  wire [2:0] _EVAL_1063;
  wire  _EVAL_1064;
  wire [2:0] _EVAL_1065;
  wire [2:0] _EVAL_1067;
  wire [1:0] _EVAL_1068;
  reg [31:0] _EVAL_1069;
  wire [12:0] _EVAL_1070;
  wire [1:0] _EVAL_1072;
  wire  _EVAL_1074;
  wire  _EVAL_1075;
  wire  _EVAL_1076;
  wire [2:0] _EVAL_1077;
  reg [12:0] _EVAL_1078;
  wire  _EVAL_1079;
  wire [31:0] _EVAL_1082;
  reg [2:0] _EVAL_1084;
  reg  _EVAL_1085;
  wire [2:0] _EVAL_1087;
  wire  _EVAL_1088;
  wire [31:0] _EVAL_1089;
  wire  _EVAL_1090;
  wire  _EVAL_1091;
  wire [2:0] _EVAL_1092;
  reg [2:0] _EVAL_1093;
  reg [2:0] _EVAL_1094;
  reg [2:0] _EVAL_1095;
  wire [2:0] _EVAL_1096;
  wire  _EVAL_1098;
  wire [2:0] _EVAL_1100;
  reg [12:0] _EVAL_1101;
  wire [3:0] _EVAL_1102;
  wire  _EVAL_1103;
  wire  _EVAL_1104;
  wire  _EVAL_1105;
  wire [12:0] _EVAL_1106;
  wire  _EVAL_1107;
  reg [12:0] _EVAL_1108;
  reg [17:0] _EVAL_1109;
  wire  _EVAL_1110;
  wire  _EVAL_1111;
  wire  _EVAL_1112;
  wire  _EVAL_1113;
  wire [8:0] _EVAL_1114;
  wire  _EVAL_1115;
  wire [31:0] _EVAL_1116;
  wire [13:0] _EVAL_1117;
  wire  _EVAL_1118;
  reg [17:0] _EVAL_1119;
  reg [12:0] _EVAL_1121;
  wire  _EVAL_1123;
  wire [29:0] _EVAL_1124;
  wire [12:0] _EVAL_1125;
  wire  _EVAL_1126;
  wire [1:0] _EVAL_1127;
  wire  _EVAL_1128;
  wire [8:0] _EVAL_1129;
  wire [2:0] _EVAL_1131;
  wire  _EVAL_1132;
  reg [2:0] _EVAL_1134;
  wire [4:0] _EVAL_1136;
  wire  _EVAL_1137;
  reg [2:0] _EVAL_1138;
  wire  _EVAL_1139;
  wire [12:0] _EVAL_1140;
  wire [2:0] _EVAL_1141;
  wire [2:0] _EVAL_1142;
  reg [12:0] _EVAL_1143;
  wire [6:0] _EVAL_1144;
  wire  _EVAL_1145;
  wire  _EVAL_1147;
  reg [1:0] _EVAL_1148;
  wire  _EVAL_1149;
  wire [4:0] _EVAL_1150;
  wire  _EVAL_1151;
  wire  _EVAL_1152;
  wire  _EVAL_1153;
  wire [12:0] _EVAL_1154;
  wire [8:0] _EVAL_1155;
  wire [6:0] _EVAL_1156;
  wire  _EVAL_1157;
  wire [15:0] _EVAL_1158;
  reg [2:0] _EVAL_1160;
  wire  _EVAL_1163;
  wire [12:0] _EVAL_1165;
  wire [4:0] _EVAL_1167;
  wire  _EVAL_1168;
  wire  _EVAL_1169;
  wire [12:0] _EVAL_1170;
  wire  _EVAL_1171;
  reg [2:0] _EVAL_1172;
  wire [5:0] _EVAL_1173;
  wire [9:0] _EVAL_1174;
  wire [2:0] _EVAL_1175;
  wire [2:0] _EVAL_1176;
  wire  _EVAL_1178;
  wire  _EVAL_1179;
  wire  _EVAL_1180;
  reg [1:0] _EVAL_1181;
  wire  _EVAL_1182;
  wire [1:0] _EVAL_1183;
  wire  _EVAL_1185;
  wire  _EVAL_1186;
  wire [2:0] _EVAL_1187;
  wire [6:0] _EVAL_1188;
  wire  _EVAL_1189;
  wire [3:0] _EVAL_1190;
  wire [2:0] _EVAL_1192;
  reg [2:0] _EVAL_1193;
  wire [2:0] _EVAL_1195;
  wire [13:0] _EVAL_1196;
  wire [17:0] _EVAL_1197;
  reg [2:0] _EVAL_1198;
  wire [2:0] _EVAL_1199;
  reg [1:0] _EVAL_1200;
  wire [2:0] _EVAL_1202;
  reg [2:0] _EVAL_1203;
  wire [2:0] _EVAL_1204;
  wire  _EVAL_1205;
  wire [2:0] _EVAL_1207;
  reg [2:0] _EVAL_1208;
  wire  _EVAL_1209;
  reg  _EVAL_1210;
  reg [2:0] _EVAL_1211;
  reg [12:0] _EVAL_1212;
  wire [17:0] _EVAL_1213;
  reg [17:0] _EVAL_1214;
  wire  _EVAL_1215;
  wire [2:0] _EVAL_1217;
  wire  _EVAL_1218;
  wire [2:0] _EVAL_1219;
  reg [1:0] _EVAL_1220;
  wire [31:0] _EVAL_1222;
  wire  _EVAL_1223;
  wire [1:0] _EVAL_1224;
  reg [1:0] _EVAL_1225;
  wire  _EVAL_1226;
  wire  _EVAL_1227;
  wire [7:0] _EVAL_1228;
  wire [2:0] _EVAL_1229;
  wire  _EVAL_1230;
  wire [2:0] _EVAL_1231;
  wire  _EVAL_1232;
  wire  _EVAL_1233;
  wire  _EVAL_1234;
  wire  _EVAL_1235;
  wire [2:0] _EVAL_1236;
  wire [12:0] _EVAL_1238;
  wire  _EVAL_1239;
  reg  _EVAL_1240;
  reg  _EVAL_1241;
  wire  _EVAL_1242;
  wire  _EVAL_1244;
  wire  _EVAL_1246;
  wire  _EVAL_1247;
  wire [2:0] _EVAL_1248;
  wire [12:0] _EVAL_1249;
  wire [2:0] _EVAL_1250;
  wire [12:0] _EVAL_1251;
  wire [2:0] _EVAL_1253;
  assign _EVAL_808__EVAL_809_addr = _EVAL_58 ^ _EVAL_1114;
  assign _EVAL_808__EVAL_809_data = _EVAL_808[_EVAL_808__EVAL_809_addr];
  assign _EVAL_808__EVAL_810_data = _EVAL_1 & _EVAL_838;
  assign _EVAL_808__EVAL_810_addr = _EVAL_79[8:0];
  assign _EVAL_808__EVAL_810_mask = 1'h1;
  assign _EVAL_808__EVAL_810_en = _EVAL_1 ? _EVAL_530 : _EVAL_756;
  assign _EVAL_179 = ~_EVAL_1089;
  assign _EVAL_1250 = _EVAL_962 ? _EVAL_893 : _EVAL_826;
  assign _EVAL_326 = _EVAL_408[29:9];
  assign _EVAL_805 = _EVAL_673 == 2'h0;
  assign _EVAL_196 = _EVAL_1034 | _EVAL_137;
  assign _EVAL_795 = {_EVAL_1173, 1'h0};
  assign _EVAL_987 = _EVAL_204[31:1];
  assign _EVAL_734 = _EVAL_635[2:0];
  assign _EVAL_359 = ~_EVAL_269;
  assign _EVAL_959 = _EVAL_1101 == _EVAL_1070;
  assign _EVAL_501 = _EVAL_1055 == 2'h3;
  assign _EVAL_398 = {_EVAL_330,_EVAL_342,_EVAL_805,_EVAL_1111,_EVAL_484,_EVAL_70,_EVAL_607};
  assign _EVAL_932 = _EVAL_1151 ? _EVAL_1078 : 13'h0;
  assign _EVAL_641 = _EVAL_34[1:0];
  assign _EVAL_1038 = _EVAL_718 ? _EVAL_911 : _EVAL_120;
  assign _EVAL = 3'h5 == _EVAL_456 ? _EVAL_634 : _EVAL_216;
  assign _EVAL_366 = 3'h5 == _EVAL_456 ? _EVAL_634 : _EVAL_216;
  assign _EVAL_69 = _EVAL_903 ? _EVAL_419 : _EVAL_122;
  assign _EVAL_869 = _EVAL_899 | _EVAL_1142;
  assign _EVAL_52 = _EVAL_1181 == 2'h3;
  assign _EVAL_1000 = _EVAL_763 | _EVAL_1058;
  assign _EVAL_814 = {_EVAL_472,_EVAL_333};
  assign _EVAL_974 = _EVAL_1040 | _EVAL_620;
  assign _EVAL_535 = _EVAL_697 | _EVAL_1013;
  assign _EVAL_920 = _EVAL_1148 == 2'h3;
  assign _EVAL_402 = _EVAL_410 ? _EVAL_41 : _EVAL_222;
  assign _EVAL_625 = _EVAL_948 ? _EVAL_1084 : 3'h0;
  assign _EVAL_572 = 8'hdd * _EVAL_25;
  assign _EVAL_516 = _EVAL_756 ? 1'h0 : _EVAL_808__EVAL_809_data;
  assign _EVAL_39 = _EVAL_515 == _EVAL_1070;
  assign _EVAL_1082 = _EVAL_549 ? _EVAL_377 : {{4'd0}, _EVAL_921};
  assign _EVAL_136 = {_EVAL_1226,_EVAL_282};
  assign _EVAL_526 = _EVAL_1248 | _EVAL_475;
  assign _EVAL_22 = _EVAL_1113 ? 1'h0 : 1'h1;
  assign _EVAL_573 = _EVAL_532[0];
  assign _EVAL_1152 = _EVAL_1068[0];
  assign _EVAL_95 = {_EVAL_14,_EVAL_265};
  assign _EVAL_1137 = _EVAL_1233 | _EVAL_939;
  assign _EVAL_543 = _EVAL_88 | _EVAL_272;
  assign _EVAL_1091 = _EVAL_997 & _EVAL_394;
  assign _EVAL_928 = ~_EVAL_756;
  assign _EVAL_1230 = _EVAL_102 | _EVAL_427;
  assign _EVAL_851 = _EVAL_947 | _EVAL_271;
  assign _EVAL_454 = {_EVAL_528,_EVAL_94,_EVAL_767,_EVAL_244,_EVAL_1246,_EVAL_276,_EVAL_533};
  assign _EVAL_1189 = ~_EVAL_1021;
  assign _EVAL_1218 = |_EVAL_735;
  assign _EVAL_1044 = _EVAL_558[2];
  assign _EVAL_743 = _EVAL_1150[4];
  assign _EVAL_375 = _EVAL_1018 ? _EVAL_900 : _EVAL_674;
  assign _EVAL_588 = _EVAL_1035 | _EVAL_1067;
  assign _EVAL_418 = _EVAL_269[1];
  assign _EVAL_289 = {_EVAL_903,_EVAL_563,_EVAL_256};
  assign _EVAL_319 = _EVAL_525 ? _EVAL_636 : 3'h0;
  assign _EVAL_460 = _EVAL_418 ? _EVAL_1138 : 3'h0;
  assign _EVAL_480 = _EVAL_459 | _EVAL_768;
  assign _EVAL_84 = _EVAL_583 & _EVAL_963;
  assign _EVAL_582 = _EVAL_547[1];
  assign _EVAL_1154 = _EVAL_840 | _EVAL_932;
  assign _EVAL_603 = _EVAL_249 | _EVAL_780;
  assign _EVAL_1087 = _EVAL_440[2:0];
  assign _EVAL_61 = 8'h1 << _EVAL_665;
  assign _EVAL_1040 = _EVAL_482 | _EVAL_1011;
  assign _EVAL_1173 = _EVAL_347 & _EVAL_1052;
  assign _EVAL_77 = _EVAL_347[3];
  assign _EVAL_988 = _EVAL_1108 == _EVAL_1070;
  assign _EVAL_494 = _EVAL_413 ? _EVAL_1189 : _EVAL_579;
  assign _EVAL_137 = _EVAL_374 & _EVAL_906;
  assign _EVAL_336 = _EVAL_35 == _EVAL_1070;
  assign _EVAL_1128 = _EVAL_987[0];
  assign _EVAL_528 = _EVAL_1048 == _EVAL_1070;
  assign _EVAL_390 = _EVAL_974 | _EVAL_1053;
  assign _EVAL_888 = _EVAL_867 ? _EVAL_823 : 3'h0;
  assign _EVAL_706 = _EVAL_787[3:2];
  assign _EVAL_55 = _EVAL_1065 | _EVAL_460;
  assign _EVAL_1224 = _EVAL_571[3:2];
  assign _EVAL_684 = _EVAL_133 == 2'h3;
  assign _EVAL_966 = _EVAL_270 ? _EVAL_1234 : _EVAL_605;
  assign _EVAL_1186 = _EVAL_819 == _EVAL_1070;
  assign _EVAL_1202 = _EVAL_1050 ? _EVAL_930 : 3'h0;
  assign _EVAL_245 = _EVAL_269[19];
  assign _EVAL_228 = _EVAL_525 ? _EVAL_414 : 3'h0;
  assign _EVAL_940 = _EVAL_951 == _EVAL_1070;
  assign _EVAL_140 = _EVAL_233 == 2'h3;
  assign _EVAL_724 = _EVAL_506 & _EVAL_1104;
  assign _EVAL_407 = |_EVAL_1173;
  assign _EVAL_232 = _EVAL_795 >> _EVAL_40;
  assign _EVAL_598 = _EVAL_509 | _EVAL_1178;
  assign _EVAL_485 = _EVAL_860 | _EVAL_373;
  assign _EVAL_256 = _EVAL_903 ? _EVAL_122 : _EVAL_278;
  assign _EVAL_1236 = _EVAL_144 ? _EVAL_664 : 3'h0;
  assign _EVAL_1100 = _EVAL_164 ? _EVAL_952 : 3'h0;
  assign _EVAL_900 = _EVAL_77 ? _EVAL_510 : 18'h0;
  assign _EVAL_497 = _EVAL_469[0];
  assign _EVAL_337 = _EVAL_1185 & _EVAL_784;
  assign _EVAL_427 = _EVAL_1233 & _EVAL_939;
  assign _EVAL_803 = _EVAL_1223 ? _EVAL_1208 : 3'h0;
  assign _EVAL_866 = _EVAL_725 | _EVAL_455;
  assign _EVAL_1196 = {_EVAL_437,_EVAL_461,_EVAL_684,_EVAL_643,_EVAL_241,_EVAL_877,_EVAL_827,_EVAL_950};
  assign _EVAL_640 = _EVAL_565 ? _EVAL_223 : 3'h0;
  assign _EVAL_461 = _EVAL_323 == 2'h3;
  assign _EVAL_62 = _EVAL_594 & _EVAL_752;
  assign _EVAL_917 = _EVAL_142 ? _EVAL_994 : _EVAL_621;
  assign _EVAL_1036 = 3'h1 == _EVAL_456 ? _EVAL_50 : _EVAL_287;
  assign _EVAL_962 = ~_EVAL_1032;
  assign _EVAL_1075 = _EVAL_1057 == _EVAL_1070;
  assign _EVAL_873 = _EVAL_724 | _EVAL_1132;
  assign _EVAL_895 = _EVAL_1124[29:9];
  assign _EVAL_297 = _EVAL_890 | _EVAL_524;
  assign _EVAL_614 = |_EVAL_329;
  assign _EVAL_1011 = _EVAL_1014 ? _EVAL_954 : 13'h0;
  assign _EVAL_649 = _EVAL_399 | _EVAL_925;
  assign _EVAL_472 = _EVAL_882[10];
  assign _EVAL_318 = _EVAL_626 ? _EVAL_151 : 13'h0;
  assign _EVAL_102 = _EVAL_1232 | _EVAL_1004;
  assign _EVAL_420 = _EVAL_34[3:2];
  assign _EVAL_801 = _EVAL_928 & _EVAL_17;
  assign _EVAL_484 = _EVAL_1055 == 2'h0;
  assign _EVAL_678 = _EVAL_115[1];
  assign _EVAL_793 = _EVAL_700 | _EVAL_425;
  assign _EVAL_840 = _EVAL_552 | _EVAL_211;
  assign _EVAL_207 = _EVAL_345 == 2'h3;
  assign _EVAL_65 = _EVAL_174 == 2'h3;
  assign _EVAL_1043 = _EVAL_158 | _EVAL_1236;
  assign _EVAL_567 = _EVAL_1124[8:0];
  assign _EVAL_382 = _EVAL_134[2];
  assign _EVAL_167 = _EVAL_344 & _EVAL_740;
  assign _EVAL_879 = _EVAL_403[1:0];
  assign _EVAL_979 = _EVAL_624[9:0];
  assign _EVAL_400 = _EVAL_1173[4:0];
  assign _EVAL_906 = _EVAL_453 | _EVAL_958;
  assign _EVAL_890 = _EVAL_496 | _EVAL_229;
  assign _EVAL_490 = _EVAL_44 ? _EVAL_1203 : 3'h0;
  assign _EVAL_405 = _EVAL_948 & _EVAL_833;
  assign _EVAL_1027 = _EVAL_33[6:0];
  assign _EVAL_253 = _EVAL_903 ? _EVAL_122 : _EVAL_184;
  assign _EVAL_937 = _EVAL_486 == 2'h3;
  assign _EVAL_547 = _EVAL_735 | _EVAL_1033;
  assign _EVAL_1033 = _EVAL_433[1:0];
  assign _EVAL_1005 = _EVAL_804 == _EVAL_1070;
  assign _EVAL_215 = _EVAL_442 ? _EVAL_517 : 13'h0;
  assign _EVAL_764 = _EVAL_832[0];
  assign _EVAL_912 = _EVAL_504[1];
  assign _EVAL_1205 = _EVAL_357 ? _EVAL_419 : _EVAL_266;
  assign _EVAL_388 = _EVAL_245 ? _EVAL_321 : 3'h0;
  assign _EVAL_786 = _EVAL_115[0];
  assign _EVAL_1110 = _EVAL_144 & _EVAL_990;
  assign _EVAL_662 = _EVAL_195 == _EVAL_1213;
  assign _EVAL_601 = _EVAL_269[6];
  assign _EVAL_949 = _EVAL_1014 & _EVAL_72;
  assign _EVAL_1025 = _EVAL_1168 | _EVAL_1110;
  assign _EVAL_998 = {_EVAL_718,_EVAL_114,_EVAL_193};
  assign _EVAL_607 = _EVAL_551 == 2'h0;
  assign _EVAL_714 = _EVAL_1025 | _EVAL_1169;
  assign _EVAL_1018 = _EVAL_166 == 3'h3;
  assign _EVAL_1176 = {_EVAL_903,_EVAL_198,_EVAL_246};
  assign _EVAL_1156 = {_EVAL_718,_EVAL_1038,_EVAL_1229};
  assign _EVAL_1065 = _EVAL_380 ? _EVAL_341 : 3'h0;
  assign _EVAL_170 = _EVAL_1199[2:1];
  assign _EVAL_284 = _EVAL_269[3];
  assign _EVAL_317 = _EVAL_534 & _EVAL_175;
  assign _EVAL_540 = _EVAL_190 | _EVAL_541;
  assign _EVAL_903 = ~_EVAL_670;
  assign _EVAL_1170 = _EVAL_156 | _EVAL_48;
  assign _EVAL_737 = _EVAL_1200 == 2'h3;
  assign _EVAL_262 = {_EVAL_792,_EVAL_751,_EVAL_711};
  assign _EVAL_259 = _EVAL_33[13:7];
  assign _EVAL_91 = {_EVAL_989,_EVAL_65,_EVAL_920,_EVAL_859,_EVAL_52,_EVAL_983,_EVAL_937,_EVAL_389,_EVAL_1196};
  assign _EVAL_164 = _EVAL_269[12];
  assign _EVAL_86 = _EVAL_551 == 2'h3;
  assign _EVAL_360 = _EVAL_766 ? _EVAL_401 : 3'h0;
  assign _EVAL_722 = _EVAL_347[0];
  assign _EVAL_30 = _EVAL_1112 & _EVAL_865;
  assign _EVAL_211 = _EVAL_396 ? _EVAL_285 : 13'h0;
  assign _EVAL_40 = _EVAL_1217 | _EVAL_444;
  assign _EVAL_28 = _EVAL_314 | _EVAL_185;
  assign _EVAL_436 = _EVAL_483 | _EVAL_109;
  assign _EVAL_733 = _EVAL_293[6:3];
  assign _EVAL_311 = _EVAL_408[8:0];
  assign _EVAL_409 = _EVAL_733[3:2];
  assign _EVAL_357 = _EVAL_1175[2];
  assign _EVAL_1163 = _EVAL_723 | _EVAL_1145;
  assign _EVAL_416 = _EVAL_1251 | _EVAL_1125;
  assign _EVAL_957 = _EVAL_885 & _EVAL_569;
  assign _EVAL_868 = _EVAL_539 ? _EVAL_349 : _EVAL_685;
  assign _EVAL_748 = _EVAL_882[6:0];
  assign _EVAL_373 = _EVAL_1118 & _EVAL_71;
  assign _EVAL_663 = _EVAL_123 == _EVAL_1070;
  assign _EVAL_139 = _EVAL_902 | _EVAL_1091;
  assign _EVAL_153 = _EVAL_855 | _EVAL_228;
  assign _EVAL_281 = _EVAL_1182 & _EVAL_260;
  assign _EVAL_1207 = {{1'd0}, _EVAL_744};
  assign _EVAL_1238 = _EVAL_789 | _EVAL_850;
  assign _EVAL_1123 = _EVAL_166 == 3'h4;
  assign _EVAL_1174 = _EVAL_928 ? {{1'd0}, _EVAL_1155} : _EVAL_131;
  assign _EVAL_1209 = _EVAL_471 | _EVAL_1230;
  assign _EVAL_489 = _EVAL_1183[0];
  assign _EVAL_1092 = _EVAL_718 ? _EVAL_818 : _EVAL_504;
  assign _EVAL_201 = _EVAL_284 ? _EVAL_99 : 13'h0;
  assign _EVAL_923 = _EVAL_565 ? _EVAL_378 : 13'h0;
  assign _EVAL_1232 = _EVAL_183 | _EVAL_167;
  assign _EVAL_1141 = _EVAL_626 ? _EVAL_919 : 3'h0;
  assign _EVAL_1076 = _EVAL_1031 | _EVAL_549;
  assign _EVAL_772 = _EVAL_956 | _EVAL_949;
  assign _EVAL_271 = _EVAL_694 & _EVAL_811;
  assign _EVAL_246 = _EVAL_903 ? _EVAL_122 : _EVAL_605;
  assign _EVAL_746 = _EVAL_867 ? _EVAL_1143 : 13'h0;
  assign _EVAL_849 = _EVAL_440[6:3];
  assign _EVAL_234 = {_EVAL_889, 6'h0};
  assign _EVAL_762 = _EVAL_1223 & _EVAL_1085;
  assign _EVAL_1142 = _EVAL_144 ? _EVAL_973 : 3'h0;
  assign _EVAL_274 = _EVAL_657 ? _EVAL_734 : 3'h5;
  assign _EVAL_342 = _EVAL_73 == 2'h0;
  assign _EVAL_613 = _EVAL_769 == 2'h3;
  assign _EVAL_694 = _EVAL_269[25];
  assign _EVAL_426 = 8'hdd * _EVAL_794;
  assign _EVAL_1105 = _EVAL_317 | _EVAL_916;
  assign _EVAL_2 = _EVAL_232[0];
  assign _EVAL_1158 = _EVAL_269[15:0];
  assign _EVAL_787 = _EVAL_1027[6:3];
  assign _EVAL_247 = _EVAL_286 == _EVAL_1070;
  assign _EVAL_875 = _EVAL_601 ? _EVAL_715 : 3'h0;
  assign _EVAL_147 = _EVAL_903 ? _EVAL_122 : _EVAL_1090;
  assign _EVAL_683 = _EVAL_911[2];
  assign _EVAL_542 = _EVAL_580[3:0];
  assign _EVAL_244 = _EVAL_726 == _EVAL_1070;
  assign _EVAL_18 = {_EVAL_941,_EVAL_180};
  assign _EVAL_612 = _EVAL_601 ? _EVAL_619 : 3'h0;
  assign _EVAL_550 = _EVAL_131[9];
  assign _EVAL_367 = _EVAL_667 | _EVAL_564;
  assign _EVAL_773 = _EVAL_869 | _EVAL_1202;
  assign _EVAL_1118 = _EVAL_786 | _EVAL_678;
  assign _EVAL_206 = _EVAL_323 == 2'h0;
  assign _EVAL_157 = _EVAL_44 ? _EVAL_848 : 13'h0;
  assign _EVAL_1022 = _EVAL_765[7:0];
  assign _EVAL_672 = _EVAL_269 & _EVAL_91;
  assign _EVAL_1003 = _EVAL_178[0];
  assign _EVAL_1089 = 32'h1 << _EVAL_1136;
  assign _EVAL_229 = _EVAL_626 ? _EVAL_857 : 3'h0;
  assign _EVAL_121 = ~_EVAL_407;
  assign _EVAL_556 = _EVAL_679 == _EVAL_1070;
  assign _EVAL_1028 = |_EVAL_984;
  assign _EVAL_697 = {{2'd0}, _EVAL_554};
  assign _EVAL_554 = {_EVAL_400,_EVAL_66};
  assign _EVAL_1072 = _EVAL_812 ? _EVAL_1009 : _EVAL_798;
  assign _EVAL_329 = _EVAL_269 & _EVAL_505;
  assign _EVAL_985 = {_EVAL_93,_EVAL_661};
  assign _EVAL_766 = _EVAL_269[24];
  assign _EVAL_411 = _EVAL_407 ? 8'h0 : _EVAL_617;
  assign _EVAL_218 = _EVAL_694 ? _EVAL_209 : 13'h0;
  assign _EVAL_482 = _EVAL_1154 | _EVAL_318;
  assign _EVAL_1233 = _EVAL_344 | _EVAL_740;
  assign _EVAL_56 = {_EVAL_539,_EVAL_907,_EVAL_868};
  assign _EVAL_1197 = _EVAL_1239 ? _EVAL_224 : _EVAL_917;
  assign _EVAL_268 = _EVAL_269[7];
  assign _EVAL_1144 = {_EVAL_59,_EVAL_298,_EVAL_695,_EVAL_929,_EVAL_821,_EVAL_210,_EVAL_350};
  assign _EVAL_1145 = _EVAL_409[1];
  assign _EVAL_500 = _EVAL_882[9:7];
  assign _EVAL_1077 = _EVAL_284 ? _EVAL_825 : 3'h0;
  assign _EVAL_1106 = _EVAL_144 ? _EVAL_1007 : 13'h0;
  assign _EVAL_190 = _EVAL_874 | _EVAL_230;
  assign _EVAL_240 = {_EVAL_1045,_EVAL_513};
  assign _EVAL_1021 = _EVAL_879[0];
  assign _EVAL_982 = _EVAL_1214 == _EVAL_306;
  assign _EVAL_296 = _EVAL_1064 | _EVAL_782;
  assign _EVAL_584 = _EVAL_631 ? _EVAL_814 : _EVAL_668;
  assign _EVAL_639 = _EVAL_30 | _EVAL_267;
  assign _EVAL_847 = _EVAL_1171 ? _EVAL_891 : 3'h0;
  assign _EVAL_941 = |_EVAL_570;
  assign _EVAL_263 = _EVAL_478 | _EVAL_1089;
  assign _EVAL_266 = _EVAL_1175[0];
  assign _EVAL_870 = _EVAL_369 | _EVAL_1247;
  assign _EVAL_561 = _EVAL_55 | _EVAL_261;
  assign _EVAL_1153 = _EVAL_135 == 2'h3;
  assign _EVAL_750 = {{4'd0}, _EVAL_570};
  assign _EVAL_1249 = _EVAL_268 ? _EVAL_107 : 13'h0;
  assign _EVAL_533 = _EVAL_779 == _EVAL_1070;
  assign _EVAL_983 = _EVAL_481 == 2'h3;
  assign _EVAL_893 = _EVAL_704[2:0];
  assign _EVAL_909 = _EVAL_130 | _EVAL_625;
  assign _EVAL_1034 = _EVAL_163 | _EVAL_632;
  assign _EVAL_544 = _EVAL_696 ? _EVAL_240 : _EVAL_136;
  assign _EVAL_413 = ~_EVAL_87;
  assign _EVAL_522 = _EVAL_356 == _EVAL_1070;
  assign _EVAL_448 = {_EVAL_988,_EVAL_522,_EVAL_1074,_EVAL_592,_EVAL_959,_EVAL_247,_EVAL_336,_EVAL_454,_EVAL_708};
  assign _EVAL_149 = _EVAL_549 ? _EVAL_830 : {{2'd0}, _EVAL_347};
  assign _EVAL_645 = _EVAL_106 | _EVAL_1137;
  assign _EVAL_1169 = _EVAL_1050 & _EVAL_487;
  assign _EVAL_830 = _EVAL_1000 | _EVAL_609;
  assign _EVAL_122 = ~_EVAL_764;
  assign _EVAL_451 = ~_EVAL_103;
  assign _EVAL_505 = {_EVAL_352,_EVAL_815,_EVAL_368,_EVAL_720,_EVAL_473,_EVAL_548,_EVAL_675,_EVAL_1144,_EVAL_1042};
  assign _EVAL_471 = _EVAL_300 | _EVAL_432;
  assign _EVAL_464 = {_EVAL_92,_EVAL_652};
  assign _EVAL_991 = _EVAL_683 ? _EVAL_1107 : _EVAL_118;
  assign _EVAL_532 = _EVAL_771[2:0];
  assign _EVAL_1183 = _EVAL_849[3:2];
  assign _EVAL_70 = _EVAL_279 == 2'h0;
  assign _EVAL_680 = _EVAL_549 & _EVAL_1227;
  assign _EVAL_989 = _EVAL_467 == 2'h3;
  assign _EVAL_1182 = ~_EVAL_152;
  assign _EVAL_712 = _EVAL_396 ? _EVAL_1160 : 3'h0;
  assign _EVAL_477 = _EVAL_1213 == _EVAL_306;
  assign _EVAL_249 = _EVAL_143 | _EVAL_847;
  assign _EVAL_386 = {_EVAL_903,_EVAL_322,_EVAL_253};
  assign _EVAL_1185 = _EVAL_269[17];
  assign _EVAL_557 = _EVAL_133 == 2'h0;
  assign _EVAL_1042 = {_EVAL_681,_EVAL_206,_EVAL_557,_EVAL_1179,_EVAL_887,_EVAL_671,_EVAL_602,_EVAL_398};
  assign _EVAL_469 = _EVAL_1087[2:1];
  assign _EVAL_939 = _EVAL_583 | _EVAL_963;
  assign _EVAL_770 = _EVAL_895[1:0];
  assign _EVAL_468 = _EVAL_558[1];
  assign _EVAL_996 = _EVAL_1214 == _EVAL_1213;
  assign _EVAL_466 = _EVAL_765[15:8];
  assign _EVAL_396 = _EVAL_269[8];
  assign _EVAL_738 = _EVAL_786 & _EVAL_678;
  assign _EVAL_264 = _EVAL_531 | _EVAL_1149;
  assign _EVAL_1190 = _EVAL_259[6:3];
  assign _EVAL_372 = _EVAL_347[1];
  assign _EVAL_34 = _EVAL_138 | _EVAL_529;
  assign _EVAL_265 = _EVAL_794[7:1];
  assign _EVAL_272 = _EVAL_525 & _EVAL_104;
  assign _EVAL_410 = _EVAL_166 == 3'h1;
  assign _EVAL_89 = _EVAL_1123 ? _EVAL_994 : _EVAL_375;
  assign _EVAL_1217 = _EVAL_526 | _EVAL_888;
  assign _EVAL_98 = _EVAL_586 == _EVAL_1213;
  assign _EVAL_59 = _EVAL_842 == 2'h0;
  assign _EVAL_119 = _EVAL_1059 | _EVAL_574;
  assign _EVAL_681 = _EVAL_835 == 2'h0;
  assign _EVAL_236 = _EVAL_667 & _EVAL_564;
  assign _EVAL_310 = _EVAL_324[2:0];
  assign _EVAL_546 = _EVAL_1225 == 2'h3;
  assign _EVAL_66 = _EVAL_1173[5];
  assign _EVAL_1014 = _EVAL_269[11];
  assign _EVAL_224 = _EVAL_914 ? _EVAL_1214 : 18'h0;
  assign _EVAL_160 = _EVAL_326[1:0];
  assign _EVAL_432 = _EVAL_800 & _EVAL_499;
  assign _EVAL_168 = {{2'd0}, _EVAL_1173};
  assign _EVAL_478 = {{4'd0}, _EVAL_921};
  assign _EVAL_1126 = _EVAL_1105 | _EVAL_575;
  assign _EVAL_575 = _EVAL_905 & _EVAL_1163;
  assign _EVAL_600 = _EVAL_913[2:1];
  assign _EVAL_581 = ~_EVAL_477;
  assign _EVAL_54 = _EVAL_162 ? _EVAL_785 : _EVAL_945;
  assign _EVAL_970 = _EVAL_1014 ? _EVAL_831 : 3'h0;
  assign _EVAL_1009 = {_EVAL_683,_EVAL_991};
  assign _EVAL_1149 = _EVAL_1127[1];
  assign _EVAL_369 = _EVAL_721 | _EVAL_927;
  assign _EVAL_178 = _EVAL_259[2:0];
  assign _EVAL_80 = _EVAL_948 ? _EVAL_43 : 3'h0;
  assign _EVAL_558 = _EVAL_748[2:0];
  assign _EVAL_538 = _EVAL_73 == 2'h3;
  assign _EVAL_254 = 3'h2 == _EVAL_456 ? _EVAL_1069 : _EVAL_1036;
  assign _EVAL_110 = _EVAL_20 ? _EVAL_95 : _EVAL_794;
  assign _EVAL_587 = {_EVAL_270,_EVAL_966};
  assign _EVAL_344 = _EVAL_1087[0];
  assign _EVAL_605 = _EVAL_717[0];
  assign _EVAL_148 = _EVAL_685[14];
  assign _EVAL_799 = _EVAL_311 ^ _EVAL_1129;
  assign _EVAL_626 = _EVAL_269[10];
  assign _EVAL_1102 = _EVAL_826 + 3'h1;
  assign _EVAL_42 = {_EVAL_1028,_EVAL_1218,_EVAL_582};
  assign _EVAL_203 = _EVAL_164 ? _EVAL_76 : 3'h0;
  assign _EVAL_440 = _EVAL_412[13:7];
  assign _EVAL_1187 = _EVAL_565 ? _EVAL_465 : 3'h0;
  assign _EVAL_1088 = _EVAL_540 | _EVAL_935;
  assign _EVAL_483 = _EVAL_944 | _EVAL_388;
  assign _EVAL_1251 = _EVAL_1165 | _EVAL_362;
  assign _EVAL_956 = _EVAL_1088 | _EVAL_258;
  assign _EVAL_453 = _EVAL_1003 | _EVAL_264;
  assign _EVAL_282 = _EVAL_1226 ? _EVAL_912 : _EVAL_1090;
  assign _EVAL_355 = _EVAL_1037 | _EVAL_116;
  assign _EVAL_1104 = _EVAL_170[1];
  assign _EVAL_796 = _EVAL_226 | _EVAL_957;
  assign _EVAL_437 = _EVAL_835 == 2'h3;
  assign _EVAL_907 = _EVAL_539 ? _EVAL_882 : _EVAL_291;
  assign _EVAL_792 = |_EVAL_138;
  assign _EVAL_1111 = _EVAL_345 == 2'h0;
  assign _EVAL_667 = _EVAL_807[0];
  assign _EVAL_36 = _EVAL_926 & _EVAL_239;
  assign _EVAL_180 = {_EVAL_862,_EVAL_313,_EVAL_1079,_EVAL_686};
  assign _EVAL_661 = _EVAL_93 ? _EVAL_587 : _EVAL_829;
  assign _EVAL_1008 = _EVAL_531 & _EVAL_1149;
  assign _EVAL_818 = {_EVAL_903,_EVAL_181,_EVAL_147};
  assign _EVAL_927 = _EVAL_418 & _EVAL_38;
  assign _EVAL_1219 = _EVAL_1185 ? _EVAL_1198 : 3'h0;
  assign _EVAL_181 = _EVAL_903 ? _EVAL_912 : _EVAL_122;
  assign _EVAL_144 = _EVAL_269[4];
  assign _EVAL_57 = ~_EVAL_516;
  assign _EVAL_100 = _EVAL_706[0];
  assign _EVAL_710 = _EVAL_26 ? _EVAL_1174 : _EVAL_131;
  assign _EVAL_585 = _EVAL_885 ? _EVAL_172 : 3'h0;
  assign _EVAL_118 = _EVAL_911[0];
  assign _EVAL_293 = _EVAL_412[6:0];
  assign _EVAL_1107 = _EVAL_911[1];
  assign _EVAL_902 = _EVAL_866 | _EVAL_1157;
  assign _EVAL_653 = _EVAL_453 & _EVAL_958;
  assign _EVAL_632 = _EVAL_896 | _EVAL_653;
  assign _EVAL_458 = _EVAL_25[7:1];
  assign _EVAL_304 = _EVAL_1199[0];
  assign _EVAL_590 = _EVAL_543 | _EVAL_337;
  assign _EVAL_609 = _EVAL_1182 ? _EVAL_535 : 8'h0;
  assign _EVAL_751 = |_EVAL_420;
  assign _EVAL_539 = ~_EVAL_743;
  assign _EVAL_412 = _EVAL_269[13:0];
  assign _EVAL_33 = _EVAL_269[27:14];
  assign _EVAL_141 = _EVAL_946 < 5'h1c;
  assign _EVAL_644 = _EVAL_106 & _EVAL_1137;
  assign _EVAL_116 = _EVAL_1151 ? _EVAL_791 : 3'h0;
  assign _EVAL_856 = _EVAL_948 ? _EVAL_406 : 13'h0;
  assign _EVAL_397 = _EVAL_269[2];
  assign _EVAL_449 = _EVAL_347[4];
  assign _EVAL_815 = _EVAL_174 == 2'h0;
  assign _EVAL_146 = _EVAL_506 | _EVAL_1104;
  assign _EVAL_134 = _EVAL_403[2:0];
  assign _EVAL_1113 = _EVAL_57 & _EVAL_614;
  assign _EVAL_93 = _EVAL_446[6];
  assign _EVAL_92 = _EVAL_500[2];
  assign _EVAL_721 = _EVAL_380 & _EVAL_972;
  assign _EVAL_1041 = _EVAL_694 ? _EVAL_593 : 3'h0;
  assign _EVAL_904 = _EVAL_380 ? _EVAL_1172 : 3'h0;
  assign _EVAL_867 = _EVAL_269[26];
  assign _EVAL_1178 = _EVAL_384 & _EVAL_367;
  assign _EVAL_226 = _EVAL_139 | _EVAL_568;
  assign _EVAL_994 = _EVAL_449 ? _EVAL_195 : 18'h0;
  assign _EVAL_660 = _EVAL_532 >= 3'h6;
  assign _EVAL_115 = _EVAL_787[1:0];
  assign _EVAL_422 = _EVAL_867 ? _EVAL_1095 : 3'h0;
  assign _EVAL_967 = _EVAL_168 | _EVAL_411;
  assign _EVAL_1247 = _EVAL_397 & _EVAL_64;
  assign _EVAL_241 = _EVAL_918 == 2'h3;
  assign _EVAL_882 = _EVAL_853[25:15];
  assign _EVAL_1013 = _EVAL_407 ? 8'h0 : _EVAL_61;
  assign _EVAL_275 = _EVAL_164 & _EVAL_595;
  assign _EVAL_691 = _EVAL_903 ? _EVAL_122 : _EVAL_118;
  assign _EVAL_624 = _EVAL_131 + 10'h1;
  assign _EVAL_571 = _EVAL_797 | _EVAL_542;
  assign _EVAL_475 = _EVAL_694 ? _EVAL_231 : 3'h0;
  assign _EVAL_442 = _EVAL_269[27];
  assign _EVAL_926 = _EVAL_913[0];
  assign _EVAL_788 = _EVAL_451 ? _EVAL_609 : _EVAL_1058;
  assign _EVAL_380 = _EVAL_269[0];
  assign _EVAL_513 = _EVAL_1045 ? _EVAL_578 : _EVAL_278;
  assign _EVAL_158 = _EVAL_776 | _EVAL_604;
  assign _EVAL_524 = _EVAL_1014 ? _EVAL_1134 : 3'h0;
  assign _EVAL_897 = _EVAL_1109 == _EVAL_1213;
  assign _EVAL_251 = _EVAL_510 == _EVAL_1213;
  assign _EVAL_947 = _EVAL_796 | _EVAL_1244;
  assign _EVAL_995 = _EVAL_1228[3];
  assign _EVAL_1063 = _EVAL_418 ? _EVAL_46 : 3'h0;
  assign _EVAL_88 = _EVAL_219 | _EVAL_405;
  assign _EVAL_79 = _EVAL_1 ? _EVAL_710 : _EVAL_131;
  assign _EVAL_800 = _EVAL_926 | _EVAL_239;
  assign _EVAL_1053 = _EVAL_1223 ? _EVAL_730 : 13'h0;
  assign _EVAL_674 = _EVAL_936 ? _EVAL_876 : _EVAL_402;
  assign _EVAL_338 = {_EVAL_413,_EVAL_1242,_EVAL_494};
  assign _EVAL_239 = _EVAL_594 | _EVAL_752;
  assign _EVAL_845 = _EVAL_1118 | _EVAL_71;
  assign _EVAL_1253 = _EVAL_718 ? _EVAL_189 : _EVAL_289;
  assign _EVAL_610 = _EVAL_962 ? _EVAL_274 : _EVAL_456;
  assign _EVAL_1124 = _EVAL_21[31:2];
  assign _EVAL_128 = _EVAL_83 | _EVAL_395;
  assign _EVAL_187 = _EVAL_867 & _EVAL_415;
  assign _EVAL_152 = |_EVAL_379;
  assign _EVAL_499 = _EVAL_905 | _EVAL_1163;
  assign _EVAL_459 = _EVAL_651 | _EVAL_612;
  assign _EVAL_1070 = _EVAL_21[13:1];
  assign _EVAL_142 = _EVAL_166 == 3'h6;
  assign _EVAL_374 = _EVAL_778 | _EVAL_845;
  assign _EVAL_754 = _EVAL_119 | _EVAL_218;
  assign _EVAL_865 = _EVAL_417[1];
  assign _EVAL_352 = _EVAL_467 == 2'h0;
  assign _EVAL_760 = _EVAL_1119 == _EVAL_1213;
  assign _EVAL_156 = _EVAL_503 | _EVAL_202;
  assign _EVAL_707 = _EVAL_7 == 2'h3;
  assign _EVAL_212 = _EVAL_1024 | _EVAL_1041;
  assign _EVAL_283 = _EVAL_1224 | _EVAL_248;
  assign _EVAL_617 = _EVAL_477 ? _EVAL_331 : {{2'd0}, _EVAL_969};
  assign _EVAL_455 = _EVAL_245 & _EVAL_1006;
  assign _EVAL_161 = _EVAL_826 < 3'h6;
  assign _EVAL_250 = _EVAL_456 < 3'h5;
  assign _EVAL_473 = _EVAL_1181 == 2'h0;
  assign _EVAL_765 = _EVAL_750 | _EVAL_1158;
  assign _EVAL_701 = _EVAL_186 | _EVAL_490;
  assign _EVAL_732 = _EVAL_212 | _EVAL_422;
  assign _EVAL_48 = _EVAL_1185 ? _EVAL_553 : 13'h0;
  assign _EVAL_1244 = _EVAL_766 & _EVAL_843;
  assign _EVAL_333 = _EVAL_472 ? {{1'd0}, _EVAL_464} : _EVAL_1231;
  assign _EVAL_1179 = _EVAL_824 == 2'h0;
  assign _EVAL_349 = {_EVAL_162,_EVAL_54,_EVAL_1188};
  assign _EVAL_943 = _EVAL_478 & _EVAL_179;
  assign _EVAL_785 = _EVAL_685[13:7];
  assign _EVAL_862 = |_EVAL_466;
  assign _EVAL_901 = _EVAL_967[3:0];
  assign _EVAL_606 = {{7'd0}, _EVAL_770};
  assign _EVAL_334 = _EVAL_1228[5];
  assign _EVAL_740 = _EVAL_497 | _EVAL_658;
  assign _EVAL_408 = _EVAL_27[31:2];
  assign _EVAL_1242 = _EVAL_413 ? _EVAL_858 : _EVAL_1189;
  assign _EVAL_685 = _EVAL_853[14:0];
  assign _EVAL_1204 = _EVAL_806 | _EVAL_1219;
  assign _EVAL_1037 = _EVAL_588 | _EVAL_1049;
  assign _EVAL_578 = _EVAL_189[1];
  assign _EVAL_1226 = _EVAL_504[2];
  assign _EVAL_548 = _EVAL_481 == 2'h0;
  assign _EVAL_670 = _EVAL_832[1];
  assign _EVAL_1229 = _EVAL_718 ? _EVAL_386 : _EVAL_558;
  assign _EVAL_529 = _EVAL_331[3:0];
  assign _EVAL_1125 = _EVAL_601 ? _EVAL_576 : 13'h0;
  assign _EVAL_682 = _EVAL_788[2];
  assign _EVAL_316 = _EVAL_885 ? _EVAL_213 : 13'h0;
  assign _EVAL_905 = _EVAL_534 | _EVAL_175;
  assign _EVAL_267 = _EVAL_489 & _EVAL_758;
  assign _EVAL_216 = 3'h4 == _EVAL_456 ? _EVAL_536 : _EVAL_813;
  assign _EVAL_389 = {_EVAL_520,_EVAL_559,_EVAL_1153,_EVAL_613,_EVAL_140,_EVAL_385,_EVAL_546};
  assign _EVAL_364 = _EVAL_250 ? _EVAL_1195 : 3'h0;
  assign _EVAL_1136 = _EVAL_141 ? _EVAL_946 : _EVAL_745;
  assign _EVAL_527 = {_EVAL_696,_EVAL_544};
  assign _EVAL_330 = _EVAL_1200 == 2'h0;
  assign _EVAL_621 = _EVAL_125 ? _EVAL_224 : _EVAL_89;
  assign _EVAL_1090 = _EVAL_504[0];
  assign _EVAL_512 = _EVAL_217 & _EVAL_960;
  assign _EVAL_574 = _EVAL_766 ? _EVAL_328 : 13'h0;
  assign _EVAL_445 = {_EVAL_903,_EVAL_69,_EVAL_1139};
  assign _EVAL_504 = _EVAL_785[2:0];
  assign _EVAL_1064 = _EVAL_709 | _EVAL_196;
  assign _EVAL_103 = _EVAL_262[0];
  assign _EVAL_361 = _EVAL_565 & _EVAL_1016;
  assign _EVAL_1132 = _EVAL_304 & _EVAL_146;
  assign _EVAL_731 = _EVAL_279 == 2'h3;
  assign _EVAL_986 = _EVAL_397 ? _EVAL_976 : 3'h0;
  assign _EVAL_1052 = {_EVAL_982,_EVAL_884,_EVAL_439,_EVAL_736,_EVAL_677,_EVAL_273};
  assign _EVAL_1035 = _EVAL_773 | _EVAL_875;
  assign _EVAL_1192 = _EVAL_44 ? _EVAL_1012 : 3'h0;
  assign _EVAL_403 = _EVAL_1150[3:0];
  assign _EVAL_744 = _EVAL_281 ? 2'h2 : 2'h1;
  assign _EVAL_248 = _EVAL_571[1:0];
  assign _EVAL_23 = _EVAL_756 ? 1'h0 : _EVAL_808__EVAL_809_data;
  assign _EVAL_150 = _EVAL_836 | _EVAL_523;
  assign _EVAL_735 = _EVAL_433[3:2];
  assign _EVAL_1139 = _EVAL_903 ? _EVAL_122 : _EVAL_266;
  assign _EVAL_509 = _EVAL_502 | _EVAL_236;
  assign _EVAL_718 = ~_EVAL_382;
  assign _EVAL_758 = _EVAL_1183[1];
  assign _EVAL_1050 = _EVAL_269[5];
  assign _EVAL_270 = _EVAL_717[2];
  assign _EVAL_87 = _EVAL_879[1];
  assign _EVAL_948 = _EVAL_269[15];
  assign _EVAL_371 = _EVAL_245 ? _EVAL_537 : 13'h0;
  assign _EVAL_997 = _EVAL_269[21];
  assign _EVAL_534 = _EVAL_775[0];
  assign _EVAL_327 = _EVAL_237 | _EVAL_215;
  assign _EVAL_884 = _EVAL_195 == _EVAL_306;
  assign _EVAL_370 = _EVAL_701 | _EVAL_585;
  assign _EVAL_916 = _EVAL_723 & _EVAL_1145;
  assign _EVAL_198 = _EVAL_903 ? _EVAL_1234 : _EVAL_122;
  assign _EVAL_273 = _EVAL_586 == _EVAL_306;
  assign _EVAL_1248 = _EVAL_370 | _EVAL_360;
  assign _EVAL_690 = _EVAL_1102[2:0];
  assign _EVAL_314 = _EVAL_851 | _EVAL_187;
  assign _EVAL_936 = _EVAL_166 == 3'h2;
  assign _EVAL_1175 = _EVAL_446[2:0];
  assign _EVAL_589 = _EVAL_442 ? _EVAL_171 : 3'h0;
  assign _EVAL_498 = _EVAL_294 == _EVAL_1070;
  assign _EVAL_210 = _EVAL_703 == 2'h0;
  assign _EVAL_620 = _EVAL_164 ? _EVAL_753 : 13'h0;
  assign _EVAL_1096 = _EVAL_904 | _EVAL_1063;
  assign _EVAL_1051 = _EVAL_788[4];
  assign _EVAL_1235 = _EVAL_903 ? _EVAL_1107 : _EVAL_122;
  assign _EVAL_520 = _EVAL_842 == 2'h3;
  assign _EVAL_564 = _EVAL_807[1];
  assign _EVAL_205 = {_EVAL_17,_EVAL_458};
  assign _EVAL_291 = {_EVAL_162,_EVAL_257,_EVAL_112};
  assign _EVAL_977 = _EVAL_387 == _EVAL_1070;
  assign _EVAL_182 = _EVAL_931 | _EVAL_762;
  assign _EVAL_565 = _EVAL_269[18];
  assign _EVAL_813 = 3'h3 == _EVAL_456 ? _EVAL_339 : _EVAL_254;
  assign _EVAL_176 = _EVAL_706[1];
  assign _EVAL_635 = _EVAL_456 - 3'h1;
  assign _EVAL_1171 = _EVAL_269[20];
  assign _EVAL_782 = _EVAL_645 & _EVAL_1215;
  assign _EVAL_312 = _EVAL_62 | _EVAL_36;
  assign _EVAL_1167 = _EVAL_331[4:0];
  assign _EVAL_836 = _EVAL_878 | _EVAL_803;
  assign _EVAL_992 = _EVAL_601 & _EVAL_622;
  assign _EVAL_877 = _EVAL_45 == 2'h3;
  assign _EVAL_968 = _EVAL_347[2];
  assign _EVAL_1098 = _EVAL_778 & _EVAL_845;
  assign _EVAL_922 = _EVAL_331[5];
  assign _EVAL_112 = _EVAL_162 ? _EVAL_1156 : _EVAL_748;
  assign _EVAL_444 = _EVAL_442 ? _EVAL_729 : 3'h0;
  assign _EVAL_963 = _EVAL_489 | _EVAL_758;
  assign _EVAL_878 = _EVAL_297 | _EVAL_203;
  assign _EVAL_530 = _EVAL_26 | _EVAL_756;
  assign _EVAL_1215 = _EVAL_374 | _EVAL_906;
  assign _EVAL_592 = _EVAL_1121 == _EVAL_1070;
  assign _EVAL_604 = _EVAL_284 ? _EVAL_627 : 3'h0;
  assign _EVAL_797 = _EVAL_580[7:4];
  assign _EVAL_58 = _EVAL_567 ^ _EVAL_606;
  assign _EVAL_961 = _EVAL_390 | _EVAL_177;
  assign _EVAL_777 = _EVAL_692 | _EVAL_640;
  assign _EVAL_1168 = _EVAL_870 | _EVAL_1039;
  assign _EVAL_1157 = _EVAL_1171 & _EVAL_759;
  assign _EVAL_1231 = {_EVAL_812,_EVAL_1072};
  assign _EVAL_790 = _EVAL_962 & _EVAL_238;
  assign _EVAL_313 = |_EVAL_797;
  assign _EVAL_260 = _EVAL_581 & _EVAL_121;
  assign _EVAL_717 = _EVAL_446[5:3];
  assign _EVAL_476 = _EVAL_1170 | _EVAL_923;
  assign _EVAL_577 = _EVAL_793 | _EVAL_566;
  assign _EVAL_747 = {_EVAL_996,_EVAL_662,_EVAL_251,_EVAL_760,_EVAL_897,_EVAL_98};
  assign _EVAL_720 = _EVAL_1220 == 2'h0;
  assign _EVAL_638 = _EVAL_32 == _EVAL_1070;
  assign _EVAL_929 = _EVAL_769 == 2'h0;
  assign _EVAL_783 = _EVAL_1151 ? _EVAL_816 : 3'h0;
  assign _EVAL_1227 = _EVAL_1182 | _EVAL_260;
  assign _EVAL_399 = _EVAL_603 | _EVAL_1192;
  assign _EVAL_945 = {_EVAL_718,_EVAL_1253,_EVAL_1092};
  assign _EVAL_820 = _EVAL_29 == _EVAL_1070;
  assign _EVAL_120 = {_EVAL_903,_EVAL_1235,_EVAL_691};
  assign _EVAL_775 = _EVAL_733[1:0];
  assign _EVAL_108 = _EVAL_37 == _EVAL_1070;
  assign _EVAL_552 = _EVAL_416 | _EVAL_1249;
  assign _EVAL_860 = _EVAL_738 | _EVAL_1147;
  assign _EVAL_1031 = _EVAL_1240 & _EVAL_1241;
  assign _EVAL_776 = _EVAL_1096 | _EVAL_986;
  assign _EVAL_219 = _EVAL_182 | _EVAL_512;
  assign _EVAL_602 = _EVAL_1010 == 2'h0;
  assign _EVAL_381 = _EVAL_1008 | _EVAL_1115;
  assign _EVAL_16 = _EVAL_794;
  assign _EVAL_1199 = _EVAL_1027[2:0];
  assign _EVAL_562 = _EVAL_7 == 2'h2;
  assign _EVAL_433 = _EVAL_984 | _EVAL_901;
  assign _EVAL_1165 = _EVAL_393 | _EVAL_1106;
  assign _EVAL_599 = {_EVAL_1197,_EVAL_1117};
  assign _EVAL_657 = _EVAL_456 > 3'h0;
  assign _EVAL_643 = _EVAL_824 == 2'h3;
  assign _EVAL_278 = _EVAL_189[0];
  assign _EVAL_1239 = _EVAL_166 == 3'h7;
  assign _EVAL_935 = _EVAL_1151 & _EVAL_474;
  assign _EVAL_106 = _EVAL_800 | _EVAL_499;
  assign _EVAL_887 = _EVAL_918 == 2'h0;
  assign _EVAL_298 = _EVAL_488 == 2'h0;
  assign _EVAL_696 = _EVAL_785[6];
  assign _EVAL_222 = _EVAL_722 ? _EVAL_586 : 18'h0;
  assign _EVAL_439 = _EVAL_510 == _EVAL_306;
  assign _EVAL_175 = _EVAL_775[1];
  assign _EVAL_568 = _EVAL_44 & _EVAL_31;
  assign _EVAL_767 = _EVAL_479 == _EVAL_1070;
  assign _EVAL_789 = _EVAL_908 | _EVAL_774;
  assign _EVAL_519 = _EVAL_577 | _EVAL_157;
  assign _EVAL_1116 = _EVAL_296 ? {{4'd0}, _EVAL_307} : _EVAL_1082;
  assign _EVAL_166 = _EVAL_732 | _EVAL_589;
  assign _EVAL_1131 = _EVAL_217 ? _EVAL_886 : 3'h0;
  assign _EVAL_257 = _EVAL_162 ? _EVAL_500 : _EVAL_338;
  assign _EVAL_583 = _EVAL_1112 | _EVAL_865;
  assign _EVAL_350 = _EVAL_1225 == 2'h0;
  assign _EVAL_1188 = _EVAL_162 ? _EVAL_998 : _EVAL_446;
  assign _EVAL_177 = _EVAL_217 ? _EVAL_741 : 13'h0;
  assign _EVAL_798 = {_EVAL_1044,_EVAL_511};
  assign _EVAL_708 = {_EVAL_638,_EVAL_498,_EVAL_940,_EVAL_39,_EVAL_663,_EVAL_470,_EVAL_1103,_EVAL_545};
  assign _EVAL_525 = _EVAL_269[16];
  assign _EVAL_331 = _EVAL_152 ? {{2'd0}, _EVAL_379} : _EVAL_535;
  assign _EVAL_768 = _EVAL_268 ? _EVAL_955 : 3'h0;
  assign _EVAL_269 = _EVAL_448 & _EVAL_921;
  assign _EVAL_71 = _EVAL_100 | _EVAL_176;
  assign _EVAL_1060 = _EVAL_1185 ? _EVAL_97 : 3'h0;
  assign _EVAL_757 = _EVAL_355 | _EVAL_1141;
  assign _EVAL_876 = _EVAL_968 ? _EVAL_1119 : 18'h0;
  assign _EVAL_362 = _EVAL_1050 ? _EVAL_155 : 13'h0;
  assign _EVAL_1195 = _EVAL_365[2:0];
  assign _EVAL_1045 = _EVAL_189[2];
  assign _EVAL_832 = _EVAL_134[1:0];
  assign _EVAL_852 = _EVAL_426[7:5];
  assign _EVAL_1140 = _EVAL_1026[13:1];
  assign _EVAL_384 = _EVAL_1152 | _EVAL_132;
  assign _EVAL_189 = _EVAL_785[5:3];
  assign _EVAL_806 = _EVAL_909 | _EVAL_319;
  assign _EVAL_723 = _EVAL_409[0];
  assign _EVAL_3 = _EVAL_790 ? _EVAL_366 : _EVAL_599;
  assign _EVAL_237 = _EVAL_754 | _EVAL_746;
  assign _EVAL_807 = _EVAL_1190[3:2];
  assign _EVAL_984 = _EVAL_967[7:4];
  assign _EVAL_1112 = _EVAL_417[0];
  assign _EVAL_594 = _EVAL_600[0];
  assign _EVAL_1150 = _EVAL_549 ? _EVAL_1136 : _EVAL_978;
  assign _EVAL_821 = _EVAL_233 == 2'h0;
  assign _EVAL_1222 = _EVAL_10 ? 32'h0 : _EVAL_1116;
  assign _EVAL_125 = _EVAL_166 == 3'h5;
  assign _EVAL_889 = _EVAL_572[7:5];
  assign _EVAL_677 = _EVAL_1109 == _EVAL_306;
  assign _EVAL_864 = _EVAL_766 ? _EVAL_173 : 3'h0;
  assign _EVAL_752 = _EVAL_600[1];
  assign _EVAL_1058 = _EVAL_260 ? _EVAL_617 : 8'h0;
  assign _EVAL_872 = _EVAL_148 ? _EVAL_527 : _EVAL_985;
  assign _EVAL_1180 = _EVAL_873 | _EVAL_485;
  assign _EVAL_700 = _EVAL_476 | _EVAL_371;
  assign _EVAL_184 = _EVAL_558[0];
  assign _EVAL_911 = _EVAL_748[5:3];
  assign _EVAL_780 = _EVAL_997 ? _EVAL_1211 : 3'h0;
  assign _EVAL_566 = _EVAL_997 ? _EVAL_199 : 13'h0;
  assign _EVAL_496 = _EVAL_688 | _EVAL_783;
  assign _EVAL_531 = _EVAL_1127[0];
  assign _EVAL_523 = _EVAL_217 ? _EVAL_1093 : 3'h0;
  assign _EVAL_101 = _EVAL_997 ? _EVAL_127 : 3'h0;
  assign _EVAL_391 = _EVAL_403[3];
  assign _EVAL_1059 = _EVAL_519 | _EVAL_316;
  assign _EVAL_1103 = _EVAL_560 == _EVAL_1070;
  assign _EVAL_1117 = {_EVAL_327, 1'h0};
  assign _EVAL_559 = _EVAL_488 == 2'h3;
  assign _EVAL_114 = _EVAL_718 ? _EVAL_717 : _EVAL_1176;
  assign _EVAL_1151 = _EVAL_269[9];
  assign _EVAL_563 = _EVAL_903 ? _EVAL_578 : _EVAL_122;
  assign _EVAL_570 = _EVAL_269[27:16];
  assign _EVAL_368 = _EVAL_1148 == 2'h0;
  assign _EVAL_829 = {_EVAL_357,_EVAL_1205};
  assign _EVAL_1147 = _EVAL_100 & _EVAL_176;
  assign _EVAL_709 = _EVAL_1209 | _EVAL_644;
  assign _EVAL_307 = _EVAL_921 & _EVAL_359;
  assign _EVAL_688 = _EVAL_480 | _EVAL_712;
  assign _EVAL_19 = ~_EVAL_1032;
  assign _EVAL_94 = _EVAL_1212 == _EVAL_1070;
  assign _EVAL_351 = _EVAL_1228[1];
  assign _EVAL_186 = _EVAL_436 | _EVAL_101;
  assign _EVAL_419 = _EVAL_1175[1];
  assign _EVAL_83 = _EVAL_698 | _EVAL_1100;
  assign _EVAL_185 = _EVAL_442 & _EVAL_301;
  assign _EVAL_1213 = _EVAL_1026[31:14];
  assign _EVAL_1020 = _EVAL_1050 ? _EVAL_1094 : 3'h0;
  assign _EVAL_163 = _EVAL_1180 | _EVAL_1098;
  assign _EVAL_41 = _EVAL_372 ? _EVAL_1109 : 18'h0;
  assign _EVAL_1115 = _EVAL_1003 & _EVAL_264;
  assign _EVAL_1074 = _EVAL_507 == _EVAL_1070;
  assign _EVAL_276 = _EVAL_993 == _EVAL_1070;
  assign _EVAL_958 = _EVAL_384 | _EVAL_367;
  assign _EVAL_899 = _EVAL_561 | _EVAL_1077;
  assign _EVAL_671 = _EVAL_45 == 2'h0;
  assign _EVAL_44 = _EVAL_269[22];
  assign _EVAL_508 = _EVAL_245 ? _EVAL_305 : 3'h0;
  assign _EVAL_1114 = {_EVAL_852, 6'h0};
  assign _EVAL_306 = _EVAL_21[31:14];
  assign _EVAL_756 = ~_EVAL_550;
  assign _EVAL_1127 = _EVAL_178[2:1];
  assign _EVAL_1039 = _EVAL_284 & _EVAL_689;
  assign _EVAL_925 = _EVAL_885 ? _EVAL_348 : 3'h0;
  assign _EVAL_395 = _EVAL_1223 ? _EVAL_1054 : 3'h0;
  assign _EVAL_692 = _EVAL_153 | _EVAL_1060;
  assign _EVAL_579 = _EVAL_500[0];
  assign _EVAL_217 = _EVAL_269[14];
  assign _EVAL_827 = _EVAL_1010 == 2'h3;
  assign _EVAL_931 = _EVAL_772 | _EVAL_275;
  assign _EVAL_944 = _EVAL_1204 | _EVAL_1187;
  assign _EVAL_470 = _EVAL_676 == _EVAL_1070;
  assign _EVAL_745 = {_EVAL_631,_EVAL_584};
  assign _EVAL_908 = _EVAL_380 ? _EVAL_159 : 13'h0;
  assign _EVAL_261 = _EVAL_397 ? _EVAL_719 : 3'h0;
  assign _EVAL_109 = _EVAL_1171 ? _EVAL_452 : 3'h0;
  assign _EVAL_950 = {_EVAL_737,_EVAL_538,_EVAL_654,_EVAL_207,_EVAL_501,_EVAL_731,_EVAL_86};
  assign _EVAL_658 = _EVAL_469[1];
  assign _EVAL_503 = _EVAL_961 | _EVAL_856;
  assign _EVAL_580 = _EVAL_466 | _EVAL_1022;
  assign _EVAL_1228 = _EVAL_451 ? _EVAL_1058 : _EVAL_609;
  assign _EVAL_686 = _EVAL_283[1];
  assign _EVAL_874 = _EVAL_714 | _EVAL_992;
  assign _EVAL_1234 = _EVAL_717[1];
  assign _EVAL_850 = _EVAL_397 ? _EVAL_642 : 13'h0;
  assign _EVAL_763 = {{2'd0}, _EVAL_347};
  assign _EVAL_1032 = _EVAL_826 == 3'h0;
  assign _EVAL_258 = _EVAL_626 & _EVAL_1210;
  assign _EVAL_377 = _EVAL_129 ? _EVAL_263 : _EVAL_943;
  assign _EVAL_1024 = _EVAL_649 | _EVAL_864;
  assign _EVAL_725 = _EVAL_590 | _EVAL_361;
  assign _EVAL_1067 = _EVAL_268 ? _EVAL_971 : 3'h0;
  assign _EVAL_969 = {_EVAL_1167,_EVAL_922};
  assign _EVAL_736 = _EVAL_1119 == _EVAL_306;
  assign _EVAL_913 = _EVAL_293[2:0];
  assign _EVAL_193 = _EVAL_718 ? _EVAL_445 : _EVAL_1175;
  assign _EVAL_1068 = _EVAL_1190[1:0];
  assign _EVAL_425 = _EVAL_1171 ? _EVAL_1030 : 13'h0;
  assign _EVAL_896 = _EVAL_381 | _EVAL_598;
  assign _EVAL_934 = _EVAL_420 | _EVAL_641;
  assign _EVAL_506 = _EVAL_170[0];
  assign _EVAL_202 = _EVAL_525 ? _EVAL_495 : 13'h0;
  assign _EVAL_511 = _EVAL_1044 ? _EVAL_468 : _EVAL_184;
  assign _EVAL_230 = _EVAL_268 & _EVAL_85;
  assign _EVAL_838 = _EVAL_26 & _EVAL_801;
  assign _EVAL_162 = ~_EVAL_391;
  assign _EVAL_541 = _EVAL_396 & _EVAL_633;
  assign _EVAL_545 = {_EVAL_820,_EVAL_977,_EVAL_1186,_EVAL_108,_EVAL_556,_EVAL_1005,_EVAL_1075};
  assign _EVAL_652 = _EVAL_92 ? _EVAL_858 : _EVAL_579;
  assign _EVAL_130 = _EVAL_128 | _EVAL_1131;
  assign _EVAL_379 = _EVAL_347 & _EVAL_747;
  assign _EVAL_855 = _EVAL_150 | _EVAL_80;
  assign _EVAL_914 = _EVAL_347[5];
  assign _EVAL_322 = _EVAL_903 ? _EVAL_468 : _EVAL_122;
  assign _EVAL_393 = _EVAL_1238 | _EVAL_201;
  assign _EVAL_698 = _EVAL_757 | _EVAL_970;
  assign _EVAL_812 = _EVAL_748[6];
  assign _EVAL_1223 = _EVAL_269[13];
  assign _EVAL_695 = _EVAL_135 == 2'h0;
  assign _EVAL_324 = _EVAL_262 + 3'h1;
  assign _EVAL_365 = _EVAL_456 + 3'h1;
  assign _EVAL_1155 = _EVAL_799 ^ _EVAL_234;
  assign _EVAL_859 = _EVAL_1220 == 2'h3;
  assign _EVAL_654 = _EVAL_673 == 2'h3;
  assign _EVAL_885 = _EVAL_269[23];
  assign _EVAL_238 = |_EVAL_672;
  assign _EVAL_1129 = {{7'd0}, _EVAL_160};
  assign _EVAL_183 = _EVAL_497 & _EVAL_658;
  assign _EVAL_132 = _EVAL_1068[1];
  assign _EVAL_502 = _EVAL_1152 & _EVAL_132;
  assign _EVAL_143 = _EVAL_777 | _EVAL_508;
  assign _EVAL_778 = _EVAL_304 | _EVAL_146;
  assign _EVAL_446 = _EVAL_685[6:0];
  assign _EVAL_858 = _EVAL_500[1];
  assign _EVAL_651 = _EVAL_1043 | _EVAL_1020;
  assign _EVAL_138 = _EVAL_331[7:4];
  assign _EVAL_300 = _EVAL_312 | _EVAL_1126;
  assign _EVAL_675 = _EVAL_486 == 2'h0;
  assign _EVAL_774 = _EVAL_418 ? _EVAL_295 : 13'h0;
  assign _EVAL_1246 = _EVAL_628 == _EVAL_1070;
  assign _EVAL_771 = _EVAL_665 + _EVAL_1207;
  assign _EVAL_417 = _EVAL_849[1:0];
  assign _EVAL_711 = _EVAL_934[1];
  assign _EVAL_631 = _EVAL_853[26];
  assign _EVAL_197 = _EVAL_788[0];
  assign _EVAL_1079 = |_EVAL_1224;
  assign _EVAL_704 = _EVAL_826 - 3'h1;
  assign _EVAL_1004 = _EVAL_639 | _EVAL_84;
  assign _EVAL_668 = {_EVAL_148,_EVAL_872};
  assign _EVAL_1049 = _EVAL_396 ? _EVAL_1193 : 3'h0;
  assign _EVAL_385 = _EVAL_703 == 2'h3;
  always @(posedge _EVAL_5) begin
    if (_EVAL_549) begin
      if (5'h6 == _EVAL_1136) begin
        _EVAL_29 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (5'h16 == _EVAL_1136) begin
        _EVAL_31 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'hd == _EVAL_1136) begin
        _EVAL_32 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (5'h15 == _EVAL_1136) begin
        _EVAL_35 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (5'h3 == _EVAL_1136) begin
        _EVAL_37 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (5'h1 == _EVAL_1136) begin
        _EVAL_38 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'hf == _EVAL_1136) begin
        _EVAL_43 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'h8 == _EVAL_1136) begin
        _EVAL_45 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'h1 == _EVAL_1136) begin
        _EVAL_46 <= _EVAL_42;
      end
    end
    if (_EVAL_6) begin
      if (_EVAL_562) begin
        if (3'h1 == _EVAL_364) begin
          _EVAL_50 <= _EVAL_13;
        end
      end
    end
    if (_EVAL_549) begin
      if (5'h2 == _EVAL_1136) begin
        _EVAL_64 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'hb == _EVAL_1136) begin
        _EVAL_72 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'h5 == _EVAL_1136) begin
        _EVAL_73 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'hc == _EVAL_1136) begin
        _EVAL_76 <= _EVAL_42;
      end
    end
    if (_EVAL_4) begin
      _EVAL_82 <= _EVAL_8;
    end
    if (_EVAL_549) begin
      if (5'h7 == _EVAL_1136) begin
        _EVAL_85 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'h11 == _EVAL_1136) begin
        _EVAL_97 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'h3 == _EVAL_1136) begin
        _EVAL_99 <= _EVAL_1070;
      end
    end
    if (_EVAL_549) begin
      if (5'h10 == _EVAL_1136) begin
        _EVAL_104 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'h7 == _EVAL_1136) begin
        _EVAL_107 <= _EVAL_1070;
      end
    end
    if (_EVAL_549) begin
      if (5'h9 == _EVAL_1136) begin
        _EVAL_123 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (5'h15 == _EVAL_1136) begin
        _EVAL_127 <= _EVAL_310;
      end
    end
    if (_EVAL_4) begin
      _EVAL_129 <= _EVAL_12;
    end
    if (_EVAL_11) begin
      _EVAL_131 <= 10'h0;
    end else if (_EVAL_756) begin
      _EVAL_131 <= _EVAL_979;
    end
    if (_EVAL_549) begin
      if (5'hb == _EVAL_1136) begin
        _EVAL_133 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'h12 == _EVAL_1136) begin
        _EVAL_135 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'ha == _EVAL_1136) begin
        _EVAL_151 <= _EVAL_1070;
      end
    end
    if (_EVAL_549) begin
      if (5'h5 == _EVAL_1136) begin
        _EVAL_155 <= _EVAL_1070;
      end
    end
    if (_EVAL_549) begin
      if (5'h0 == _EVAL_1136) begin
        _EVAL_159 <= _EVAL_1070;
      end
    end
    if (_EVAL_549) begin
      if (5'h1b == _EVAL_1136) begin
        _EVAL_171 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'h17 == _EVAL_1136) begin
        _EVAL_172 <= _EVAL_310;
      end
    end
    if (_EVAL_549) begin
      if (5'h18 == _EVAL_1136) begin
        _EVAL_173 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'h1a == _EVAL_1136) begin
        _EVAL_174 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (_EVAL_1051) begin
        if (_EVAL_451) begin
          _EVAL_195 <= _EVAL_1213;
        end else begin
          _EVAL_195 <= _EVAL_306;
        end
      end
    end
    if (_EVAL_549) begin
      if (5'h15 == _EVAL_1136) begin
        _EVAL_199 <= _EVAL_1070;
      end
    end
    if (_EVAL_4) begin
      _EVAL_204 <= _EVAL_9;
    end
    if (_EVAL_549) begin
      if (5'h19 == _EVAL_1136) begin
        _EVAL_209 <= _EVAL_1070;
      end
    end
    if (_EVAL_549) begin
      if (5'h17 == _EVAL_1136) begin
        _EVAL_213 <= _EVAL_1070;
      end
    end
    if (_EVAL_549) begin
      if (5'h12 == _EVAL_1136) begin
        _EVAL_223 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'h19 == _EVAL_1136) begin
        _EVAL_231 <= _EVAL_310;
      end
    end
    if (_EVAL_549) begin
      if (5'h10 == _EVAL_1136) begin
        _EVAL_233 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'h1 == _EVAL_1136) begin
        _EVAL_279 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'h8 == _EVAL_1136) begin
        _EVAL_285 <= _EVAL_1070;
      end
    end
    if (_EVAL_549) begin
      if (5'h16 == _EVAL_1136) begin
        _EVAL_286 <= _EVAL_1140;
      end
    end
    if (_EVAL_6) begin
      if (_EVAL_562) begin
        if (3'h0 == _EVAL_364) begin
          _EVAL_287 <= _EVAL_13;
        end
      end
    end
    if (_EVAL_549) begin
      if (5'hc == _EVAL_1136) begin
        _EVAL_294 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (5'h1 == _EVAL_1136) begin
        _EVAL_295 <= _EVAL_1070;
      end
    end
    if (_EVAL_549) begin
      if (5'h1b == _EVAL_1136) begin
        _EVAL_301 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'h13 == _EVAL_1136) begin
        _EVAL_305 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'h13 == _EVAL_1136) begin
        _EVAL_321 <= _EVAL_310;
      end
    end
    if (_EVAL_549) begin
      if (5'hc == _EVAL_1136) begin
        _EVAL_323 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'h18 == _EVAL_1136) begin
        _EVAL_328 <= _EVAL_1070;
      end
    end
    if (_EVAL_6) begin
      if (_EVAL_562) begin
        if (3'h3 == _EVAL_364) begin
          _EVAL_339 <= _EVAL_13;
        end
      end
    end
    if (_EVAL_549) begin
      if (5'h0 == _EVAL_1136) begin
        _EVAL_341 <= _EVAL_310;
      end
    end
    if (_EVAL_549) begin
      if (5'h3 == _EVAL_1136) begin
        _EVAL_345 <= _EVAL_82;
      end
    end
    if (_EVAL_11) begin
      _EVAL_347 <= 6'h0;
    end else begin
      _EVAL_347 <= _EVAL_149[5:0];
    end
    if (_EVAL_549) begin
      if (5'h17 == _EVAL_1136) begin
        _EVAL_348 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'h1a == _EVAL_1136) begin
        _EVAL_356 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (5'h12 == _EVAL_1136) begin
        _EVAL_378 <= _EVAL_1070;
      end
    end
    if (_EVAL_549) begin
      if (5'h5 == _EVAL_1136) begin
        _EVAL_387 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (5'h15 == _EVAL_1136) begin
        _EVAL_394 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'h18 == _EVAL_1136) begin
        _EVAL_401 <= _EVAL_310;
      end
    end
    if (_EVAL_549) begin
      if (5'hf == _EVAL_1136) begin
        _EVAL_406 <= _EVAL_1070;
      end
    end
    if (_EVAL_549) begin
      if (5'h10 == _EVAL_1136) begin
        _EVAL_414 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'h1a == _EVAL_1136) begin
        _EVAL_415 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'h14 == _EVAL_1136) begin
        _EVAL_452 <= _EVAL_310;
      end
    end
    if (_EVAL_11) begin
      _EVAL_456 <= 3'h0;
    end else if (_EVAL_6) begin
      if (_EVAL_562) begin
        if (_EVAL_250) begin
          _EVAL_456 <= _EVAL_1195;
        end else begin
          _EVAL_456 <= 3'h0;
        end
      end else if (_EVAL_707) begin
        _EVAL_456 <= _EVAL_610;
      end
    end
    if (_EVAL_549) begin
      if (5'h12 == _EVAL_1136) begin
        _EVAL_465 <= _EVAL_310;
      end
    end
    if (_EVAL_549) begin
      if (5'h1b == _EVAL_1136) begin
        _EVAL_467 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'h9 == _EVAL_1136) begin
        _EVAL_474 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'h12 == _EVAL_1136) begin
        _EVAL_479 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (5'h16 == _EVAL_1136) begin
        _EVAL_481 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'h15 == _EVAL_1136) begin
        _EVAL_486 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'h5 == _EVAL_1136) begin
        _EVAL_487 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'h13 == _EVAL_1136) begin
        _EVAL_488 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'h10 == _EVAL_1136) begin
        _EVAL_495 <= _EVAL_1070;
      end
    end
    if (_EVAL_549) begin
      if (5'h19 == _EVAL_1136) begin
        _EVAL_507 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (_EVAL_995) begin
        if (_EVAL_451) begin
          _EVAL_510 <= _EVAL_306;
        end else begin
          _EVAL_510 <= _EVAL_1213;
        end
      end
    end
    if (_EVAL_549) begin
      if (5'ha == _EVAL_1136) begin
        _EVAL_515 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (5'h1b == _EVAL_1136) begin
        _EVAL_517 <= _EVAL_1070;
      end
    end
    if (_EVAL_6) begin
      if (_EVAL_562) begin
        if (3'h4 == _EVAL_364) begin
          _EVAL_536 <= _EVAL_13;
        end
      end
    end
    if (_EVAL_549) begin
      if (5'h13 == _EVAL_1136) begin
        _EVAL_537 <= _EVAL_1070;
      end
    end
    if (_EVAL_11) begin
      _EVAL_549 <= 1'h0;
    end else begin
      _EVAL_549 <= _EVAL_4;
    end
    if (_EVAL_549) begin
      if (5'h0 == _EVAL_1136) begin
        _EVAL_551 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'h11 == _EVAL_1136) begin
        _EVAL_553 <= _EVAL_1070;
      end
    end
    if (_EVAL_549) begin
      if (5'h7 == _EVAL_1136) begin
        _EVAL_560 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (5'h17 == _EVAL_1136) begin
        _EVAL_569 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'h6 == _EVAL_1136) begin
        _EVAL_576 <= _EVAL_1070;
      end
    end
    if (_EVAL_549) begin
      if (_EVAL_197) begin
        if (_EVAL_451) begin
          _EVAL_586 <= _EVAL_1213;
        end else begin
          _EVAL_586 <= _EVAL_306;
        end
      end
    end
    if (_EVAL_549) begin
      if (5'h19 == _EVAL_1136) begin
        _EVAL_593 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'hc == _EVAL_1136) begin
        _EVAL_595 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'h6 == _EVAL_1136) begin
        _EVAL_619 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'h6 == _EVAL_1136) begin
        _EVAL_622 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'h3 == _EVAL_1136) begin
        _EVAL_627 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'h10 == _EVAL_1136) begin
        _EVAL_628 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (5'h8 == _EVAL_1136) begin
        _EVAL_633 <= _EVAL_1128;
      end
    end
    if (_EVAL_6) begin
      if (_EVAL_562) begin
        if (3'h5 == _EVAL_364) begin
          _EVAL_634 <= _EVAL_13;
        end
      end
    end
    if (_EVAL_549) begin
      if (5'h10 == _EVAL_1136) begin
        _EVAL_636 <= _EVAL_310;
      end
    end
    if (_EVAL_549) begin
      if (5'h2 == _EVAL_1136) begin
        _EVAL_642 <= _EVAL_1070;
      end
    end
    if (_EVAL_549) begin
      if (5'h4 == _EVAL_1136) begin
        _EVAL_664 <= _EVAL_42;
      end
    end
    if (_EVAL_11) begin
      _EVAL_665 <= 3'h0;
    end else if (_EVAL_680) begin
      if (_EVAL_660) begin
        _EVAL_665 <= {{2'd0}, _EVAL_573};
      end else begin
        _EVAL_665 <= _EVAL_532;
      end
    end
    if (_EVAL_549) begin
      if (5'h4 == _EVAL_1136) begin
        _EVAL_673 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'h8 == _EVAL_1136) begin
        _EVAL_676 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (5'h2 == _EVAL_1136) begin
        _EVAL_679 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (5'h3 == _EVAL_1136) begin
        _EVAL_689 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'hf == _EVAL_1136) begin
        _EVAL_703 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'h6 == _EVAL_1136) begin
        _EVAL_715 <= _EVAL_310;
      end
    end
    if (_EVAL_549) begin
      if (5'h2 == _EVAL_1136) begin
        _EVAL_719 <= _EVAL_310;
      end
    end
    if (_EVAL_549) begin
      if (5'h11 == _EVAL_1136) begin
        _EVAL_726 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (5'h1b == _EVAL_1136) begin
        _EVAL_729 <= _EVAL_310;
      end
    end
    if (_EVAL_549) begin
      if (5'hd == _EVAL_1136) begin
        _EVAL_730 <= _EVAL_1070;
      end
    end
    if (_EVAL_549) begin
      if (5'he == _EVAL_1136) begin
        _EVAL_741 <= _EVAL_1070;
      end
    end
    if (_EVAL_549) begin
      if (5'hc == _EVAL_1136) begin
        _EVAL_753 <= _EVAL_1070;
      end
    end
    if (_EVAL_549) begin
      if (5'h14 == _EVAL_1136) begin
        _EVAL_759 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'h11 == _EVAL_1136) begin
        _EVAL_769 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'he == _EVAL_1136) begin
        _EVAL_779 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (5'h11 == _EVAL_1136) begin
        _EVAL_784 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'h9 == _EVAL_1136) begin
        _EVAL_791 <= _EVAL_310;
      end
    end
    if (_EVAL_11) begin
      _EVAL_794 <= 8'h0;
    end else if (_EVAL_1) begin
      if (_EVAL_26) begin
        if (_EVAL_0) begin
          _EVAL_794 <= _EVAL_205;
        end else begin
          _EVAL_794 <= _EVAL_110;
        end
      end else if (_EVAL_0) begin
        _EVAL_794 <= _EVAL_25;
      end else begin
        _EVAL_794 <= _EVAL_110;
      end
    end else begin
      _EVAL_794 <= _EVAL_110;
    end
    if (_EVAL_549) begin
      if (5'h1 == _EVAL_1136) begin
        _EVAL_804 <= _EVAL_1140;
      end
    end
    if(_EVAL_808__EVAL_810_en & _EVAL_808__EVAL_810_mask) begin
      _EVAL_808[_EVAL_808__EVAL_810_addr] <= _EVAL_808__EVAL_810_data;
    end
    if (_EVAL_549) begin
      if (5'h19 == _EVAL_1136) begin
        _EVAL_811 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'h9 == _EVAL_1136) begin
        _EVAL_816 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'h4 == _EVAL_1136) begin
        _EVAL_819 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (5'h1a == _EVAL_1136) begin
        _EVAL_823 <= _EVAL_310;
      end
    end
    if (_EVAL_549) begin
      if (5'ha == _EVAL_1136) begin
        _EVAL_824 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'h3 == _EVAL_1136) begin
        _EVAL_825 <= _EVAL_310;
      end
    end
    if (_EVAL_11) begin
      _EVAL_826 <= 3'h0;
    end else if (_EVAL_6) begin
      if (_EVAL_562) begin
        if (_EVAL_161) begin
          _EVAL_826 <= _EVAL_690;
        end
      end else if (_EVAL_707) begin
        _EVAL_826 <= _EVAL_1250;
      end
    end
    if (_EVAL_549) begin
      if (5'hb == _EVAL_1136) begin
        _EVAL_831 <= _EVAL_310;
      end
    end
    if (_EVAL_549) begin
      if (5'hf == _EVAL_1136) begin
        _EVAL_833 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'hd == _EVAL_1136) begin
        _EVAL_835 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'h14 == _EVAL_1136) begin
        _EVAL_842 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'h18 == _EVAL_1136) begin
        _EVAL_843 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'h16 == _EVAL_1136) begin
        _EVAL_848 <= _EVAL_1070;
      end
    end
    if (_EVAL_11) begin
      _EVAL_853 <= 27'h0;
    end else if (_EVAL_1076) begin
      _EVAL_853 <= _EVAL_56;
    end
    if (_EVAL_549) begin
      if (5'ha == _EVAL_1136) begin
        _EVAL_857 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'he == _EVAL_1136) begin
        _EVAL_886 <= _EVAL_310;
      end
    end
    if (_EVAL_549) begin
      if (5'h14 == _EVAL_1136) begin
        _EVAL_891 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'h9 == _EVAL_1136) begin
        _EVAL_918 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'ha == _EVAL_1136) begin
        _EVAL_919 <= _EVAL_310;
      end
    end
    if (_EVAL_11) begin
      _EVAL_921 <= 28'h0;
    end else begin
      _EVAL_921 <= _EVAL_1222[27:0];
    end
    if (_EVAL_549) begin
      if (5'h5 == _EVAL_1136) begin
        _EVAL_930 <= _EVAL_310;
      end
    end
    if (_EVAL_4) begin
      _EVAL_946 <= _EVAL_24;
    end
    if (_EVAL_549) begin
      if (5'hb == _EVAL_1136) begin
        _EVAL_951 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (5'hc == _EVAL_1136) begin
        _EVAL_952 <= _EVAL_310;
      end
    end
    if (_EVAL_549) begin
      if (5'hb == _EVAL_1136) begin
        _EVAL_954 <= _EVAL_1070;
      end
    end
    if (_EVAL_549) begin
      if (5'h7 == _EVAL_1136) begin
        _EVAL_955 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'he == _EVAL_1136) begin
        _EVAL_960 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'h7 == _EVAL_1136) begin
        _EVAL_971 <= _EVAL_310;
      end
    end
    if (_EVAL_549) begin
      if (5'h0 == _EVAL_1136) begin
        _EVAL_972 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'h4 == _EVAL_1136) begin
        _EVAL_973 <= _EVAL_310;
      end
    end
    if (_EVAL_549) begin
      if (5'h2 == _EVAL_1136) begin
        _EVAL_976 <= _EVAL_42;
      end
    end
    if (_EVAL_2) begin
      _EVAL_978 <= _EVAL_18;
    end
    if (_EVAL_549) begin
      if (5'h4 == _EVAL_1136) begin
        _EVAL_990 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'hf == _EVAL_1136) begin
        _EVAL_993 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (5'h13 == _EVAL_1136) begin
        _EVAL_1006 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'h4 == _EVAL_1136) begin
        _EVAL_1007 <= _EVAL_1070;
      end
    end
    if (_EVAL_549) begin
      if (5'h7 == _EVAL_1136) begin
        _EVAL_1010 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'h16 == _EVAL_1136) begin
        _EVAL_1012 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'h12 == _EVAL_1136) begin
        _EVAL_1016 <= _EVAL_1128;
      end
    end
    if (_EVAL_4) begin
      _EVAL_1026 <= _EVAL_15;
    end
    if (_EVAL_549) begin
      if (5'h14 == _EVAL_1136) begin
        _EVAL_1030 <= _EVAL_1070;
      end
    end
    if (_EVAL_549) begin
      if (5'h14 == _EVAL_1136) begin
        _EVAL_1048 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (5'hd == _EVAL_1136) begin
        _EVAL_1054 <= _EVAL_310;
      end
    end
    if (_EVAL_549) begin
      if (5'h2 == _EVAL_1136) begin
        _EVAL_1055 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'h0 == _EVAL_1136) begin
        _EVAL_1057 <= _EVAL_1140;
      end
    end
    if (_EVAL_6) begin
      if (_EVAL_562) begin
        if (3'h2 == _EVAL_364) begin
          _EVAL_1069 <= _EVAL_13;
        end
      end
    end
    if (_EVAL_549) begin
      if (5'h9 == _EVAL_1136) begin
        _EVAL_1078 <= _EVAL_1070;
      end
    end
    if (_EVAL_549) begin
      if (5'hf == _EVAL_1136) begin
        _EVAL_1084 <= _EVAL_310;
      end
    end
    if (_EVAL_549) begin
      if (5'hd == _EVAL_1136) begin
        _EVAL_1085 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'he == _EVAL_1136) begin
        _EVAL_1093 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'h5 == _EVAL_1136) begin
        _EVAL_1094 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'h1a == _EVAL_1136) begin
        _EVAL_1095 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'h17 == _EVAL_1136) begin
        _EVAL_1101 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (5'h1b == _EVAL_1136) begin
        _EVAL_1108 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (_EVAL_351) begin
        if (_EVAL_451) begin
          _EVAL_1109 <= _EVAL_306;
        end else begin
          _EVAL_1109 <= _EVAL_1213;
        end
      end
    end
    if (_EVAL_549) begin
      if (_EVAL_682) begin
        if (_EVAL_451) begin
          _EVAL_1119 <= _EVAL_1213;
        end else begin
          _EVAL_1119 <= _EVAL_306;
        end
      end
    end
    if (_EVAL_549) begin
      if (5'h18 == _EVAL_1136) begin
        _EVAL_1121 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (5'hb == _EVAL_1136) begin
        _EVAL_1134 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'h1 == _EVAL_1136) begin
        _EVAL_1138 <= _EVAL_310;
      end
    end
    if (_EVAL_549) begin
      if (5'h1a == _EVAL_1136) begin
        _EVAL_1143 <= _EVAL_1070;
      end
    end
    if (_EVAL_549) begin
      if (5'h19 == _EVAL_1136) begin
        _EVAL_1148 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'h8 == _EVAL_1136) begin
        _EVAL_1160 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'h0 == _EVAL_1136) begin
        _EVAL_1172 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'h17 == _EVAL_1136) begin
        _EVAL_1181 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'h8 == _EVAL_1136) begin
        _EVAL_1193 <= _EVAL_310;
      end
    end
    if (_EVAL_549) begin
      if (5'h11 == _EVAL_1136) begin
        _EVAL_1198 <= _EVAL_310;
      end
    end
    if (_EVAL_549) begin
      if (5'h6 == _EVAL_1136) begin
        _EVAL_1200 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'h16 == _EVAL_1136) begin
        _EVAL_1203 <= _EVAL_310;
      end
    end
    if (_EVAL_549) begin
      if (5'hd == _EVAL_1136) begin
        _EVAL_1208 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'ha == _EVAL_1136) begin
        _EVAL_1210 <= _EVAL_1128;
      end
    end
    if (_EVAL_549) begin
      if (5'h15 == _EVAL_1136) begin
        _EVAL_1211 <= _EVAL_42;
      end
    end
    if (_EVAL_549) begin
      if (5'h13 == _EVAL_1136) begin
        _EVAL_1212 <= _EVAL_1140;
      end
    end
    if (_EVAL_549) begin
      if (_EVAL_334) begin
        if (_EVAL_451) begin
          _EVAL_1214 <= _EVAL_306;
        end else begin
          _EVAL_1214 <= _EVAL_1213;
        end
      end
    end
    if (_EVAL_549) begin
      if (5'h18 == _EVAL_1136) begin
        _EVAL_1220 <= _EVAL_82;
      end
    end
    if (_EVAL_549) begin
      if (5'he == _EVAL_1136) begin
        _EVAL_1225 <= _EVAL_82;
      end
    end
    if (_EVAL_11) begin
      _EVAL_1240 <= 1'h0;
    end else begin
      _EVAL_1240 <= _EVAL_2;
    end
    if (_EVAL_2) begin
      _EVAL_1241 <= _EVAL_22;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_120 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    _EVAL_808[initvar] = _RAND_120[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_29 = _RAND_0[12:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_31 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_32 = _RAND_2[12:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_35 = _RAND_3[12:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_37 = _RAND_4[12:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_38 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_43 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_45 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_46 = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_50 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_64 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_72 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_73 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_76 = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_82 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_85 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_97 = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  _EVAL_99 = _RAND_17[12:0];
  _RAND_18 = {1{`RANDOM}};
  _EVAL_104 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  _EVAL_107 = _RAND_19[12:0];
  _RAND_20 = {1{`RANDOM}};
  _EVAL_123 = _RAND_20[12:0];
  _RAND_21 = {1{`RANDOM}};
  _EVAL_127 = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  _EVAL_129 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  _EVAL_131 = _RAND_23[9:0];
  _RAND_24 = {1{`RANDOM}};
  _EVAL_133 = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  _EVAL_135 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  _EVAL_151 = _RAND_26[12:0];
  _RAND_27 = {1{`RANDOM}};
  _EVAL_155 = _RAND_27[12:0];
  _RAND_28 = {1{`RANDOM}};
  _EVAL_159 = _RAND_28[12:0];
  _RAND_29 = {1{`RANDOM}};
  _EVAL_171 = _RAND_29[2:0];
  _RAND_30 = {1{`RANDOM}};
  _EVAL_172 = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  _EVAL_173 = _RAND_31[2:0];
  _RAND_32 = {1{`RANDOM}};
  _EVAL_174 = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  _EVAL_195 = _RAND_33[17:0];
  _RAND_34 = {1{`RANDOM}};
  _EVAL_199 = _RAND_34[12:0];
  _RAND_35 = {1{`RANDOM}};
  _EVAL_204 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  _EVAL_209 = _RAND_36[12:0];
  _RAND_37 = {1{`RANDOM}};
  _EVAL_213 = _RAND_37[12:0];
  _RAND_38 = {1{`RANDOM}};
  _EVAL_223 = _RAND_38[2:0];
  _RAND_39 = {1{`RANDOM}};
  _EVAL_231 = _RAND_39[2:0];
  _RAND_40 = {1{`RANDOM}};
  _EVAL_233 = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  _EVAL_279 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  _EVAL_285 = _RAND_42[12:0];
  _RAND_43 = {1{`RANDOM}};
  _EVAL_286 = _RAND_43[12:0];
  _RAND_44 = {1{`RANDOM}};
  _EVAL_287 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  _EVAL_294 = _RAND_45[12:0];
  _RAND_46 = {1{`RANDOM}};
  _EVAL_295 = _RAND_46[12:0];
  _RAND_47 = {1{`RANDOM}};
  _EVAL_301 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  _EVAL_305 = _RAND_48[2:0];
  _RAND_49 = {1{`RANDOM}};
  _EVAL_321 = _RAND_49[2:0];
  _RAND_50 = {1{`RANDOM}};
  _EVAL_323 = _RAND_50[1:0];
  _RAND_51 = {1{`RANDOM}};
  _EVAL_328 = _RAND_51[12:0];
  _RAND_52 = {1{`RANDOM}};
  _EVAL_339 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  _EVAL_341 = _RAND_53[2:0];
  _RAND_54 = {1{`RANDOM}};
  _EVAL_345 = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  _EVAL_347 = _RAND_55[5:0];
  _RAND_56 = {1{`RANDOM}};
  _EVAL_348 = _RAND_56[2:0];
  _RAND_57 = {1{`RANDOM}};
  _EVAL_356 = _RAND_57[12:0];
  _RAND_58 = {1{`RANDOM}};
  _EVAL_378 = _RAND_58[12:0];
  _RAND_59 = {1{`RANDOM}};
  _EVAL_387 = _RAND_59[12:0];
  _RAND_60 = {1{`RANDOM}};
  _EVAL_394 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  _EVAL_401 = _RAND_61[2:0];
  _RAND_62 = {1{`RANDOM}};
  _EVAL_406 = _RAND_62[12:0];
  _RAND_63 = {1{`RANDOM}};
  _EVAL_414 = _RAND_63[2:0];
  _RAND_64 = {1{`RANDOM}};
  _EVAL_415 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  _EVAL_452 = _RAND_65[2:0];
  _RAND_66 = {1{`RANDOM}};
  _EVAL_456 = _RAND_66[2:0];
  _RAND_67 = {1{`RANDOM}};
  _EVAL_465 = _RAND_67[2:0];
  _RAND_68 = {1{`RANDOM}};
  _EVAL_467 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  _EVAL_474 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  _EVAL_479 = _RAND_70[12:0];
  _RAND_71 = {1{`RANDOM}};
  _EVAL_481 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  _EVAL_486 = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  _EVAL_487 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  _EVAL_488 = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  _EVAL_495 = _RAND_75[12:0];
  _RAND_76 = {1{`RANDOM}};
  _EVAL_507 = _RAND_76[12:0];
  _RAND_77 = {1{`RANDOM}};
  _EVAL_510 = _RAND_77[17:0];
  _RAND_78 = {1{`RANDOM}};
  _EVAL_515 = _RAND_78[12:0];
  _RAND_79 = {1{`RANDOM}};
  _EVAL_517 = _RAND_79[12:0];
  _RAND_80 = {1{`RANDOM}};
  _EVAL_536 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  _EVAL_537 = _RAND_81[12:0];
  _RAND_82 = {1{`RANDOM}};
  _EVAL_549 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  _EVAL_551 = _RAND_83[1:0];
  _RAND_84 = {1{`RANDOM}};
  _EVAL_553 = _RAND_84[12:0];
  _RAND_85 = {1{`RANDOM}};
  _EVAL_560 = _RAND_85[12:0];
  _RAND_86 = {1{`RANDOM}};
  _EVAL_569 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  _EVAL_576 = _RAND_87[12:0];
  _RAND_88 = {1{`RANDOM}};
  _EVAL_586 = _RAND_88[17:0];
  _RAND_89 = {1{`RANDOM}};
  _EVAL_593 = _RAND_89[2:0];
  _RAND_90 = {1{`RANDOM}};
  _EVAL_595 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  _EVAL_619 = _RAND_91[2:0];
  _RAND_92 = {1{`RANDOM}};
  _EVAL_622 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  _EVAL_627 = _RAND_93[2:0];
  _RAND_94 = {1{`RANDOM}};
  _EVAL_628 = _RAND_94[12:0];
  _RAND_95 = {1{`RANDOM}};
  _EVAL_633 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  _EVAL_634 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  _EVAL_636 = _RAND_97[2:0];
  _RAND_98 = {1{`RANDOM}};
  _EVAL_642 = _RAND_98[12:0];
  _RAND_99 = {1{`RANDOM}};
  _EVAL_664 = _RAND_99[2:0];
  _RAND_100 = {1{`RANDOM}};
  _EVAL_665 = _RAND_100[2:0];
  _RAND_101 = {1{`RANDOM}};
  _EVAL_673 = _RAND_101[1:0];
  _RAND_102 = {1{`RANDOM}};
  _EVAL_676 = _RAND_102[12:0];
  _RAND_103 = {1{`RANDOM}};
  _EVAL_679 = _RAND_103[12:0];
  _RAND_104 = {1{`RANDOM}};
  _EVAL_689 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  _EVAL_703 = _RAND_105[1:0];
  _RAND_106 = {1{`RANDOM}};
  _EVAL_715 = _RAND_106[2:0];
  _RAND_107 = {1{`RANDOM}};
  _EVAL_719 = _RAND_107[2:0];
  _RAND_108 = {1{`RANDOM}};
  _EVAL_726 = _RAND_108[12:0];
  _RAND_109 = {1{`RANDOM}};
  _EVAL_729 = _RAND_109[2:0];
  _RAND_110 = {1{`RANDOM}};
  _EVAL_730 = _RAND_110[12:0];
  _RAND_111 = {1{`RANDOM}};
  _EVAL_741 = _RAND_111[12:0];
  _RAND_112 = {1{`RANDOM}};
  _EVAL_753 = _RAND_112[12:0];
  _RAND_113 = {1{`RANDOM}};
  _EVAL_759 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  _EVAL_769 = _RAND_114[1:0];
  _RAND_115 = {1{`RANDOM}};
  _EVAL_779 = _RAND_115[12:0];
  _RAND_116 = {1{`RANDOM}};
  _EVAL_784 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  _EVAL_791 = _RAND_117[2:0];
  _RAND_118 = {1{`RANDOM}};
  _EVAL_794 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  _EVAL_804 = _RAND_119[12:0];
  _RAND_121 = {1{`RANDOM}};
  _EVAL_811 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  _EVAL_816 = _RAND_122[2:0];
  _RAND_123 = {1{`RANDOM}};
  _EVAL_819 = _RAND_123[12:0];
  _RAND_124 = {1{`RANDOM}};
  _EVAL_823 = _RAND_124[2:0];
  _RAND_125 = {1{`RANDOM}};
  _EVAL_824 = _RAND_125[1:0];
  _RAND_126 = {1{`RANDOM}};
  _EVAL_825 = _RAND_126[2:0];
  _RAND_127 = {1{`RANDOM}};
  _EVAL_826 = _RAND_127[2:0];
  _RAND_128 = {1{`RANDOM}};
  _EVAL_831 = _RAND_128[2:0];
  _RAND_129 = {1{`RANDOM}};
  _EVAL_833 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  _EVAL_835 = _RAND_130[1:0];
  _RAND_131 = {1{`RANDOM}};
  _EVAL_842 = _RAND_131[1:0];
  _RAND_132 = {1{`RANDOM}};
  _EVAL_843 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  _EVAL_848 = _RAND_133[12:0];
  _RAND_134 = {1{`RANDOM}};
  _EVAL_853 = _RAND_134[26:0];
  _RAND_135 = {1{`RANDOM}};
  _EVAL_857 = _RAND_135[2:0];
  _RAND_136 = {1{`RANDOM}};
  _EVAL_886 = _RAND_136[2:0];
  _RAND_137 = {1{`RANDOM}};
  _EVAL_891 = _RAND_137[2:0];
  _RAND_138 = {1{`RANDOM}};
  _EVAL_918 = _RAND_138[1:0];
  _RAND_139 = {1{`RANDOM}};
  _EVAL_919 = _RAND_139[2:0];
  _RAND_140 = {1{`RANDOM}};
  _EVAL_921 = _RAND_140[27:0];
  _RAND_141 = {1{`RANDOM}};
  _EVAL_930 = _RAND_141[2:0];
  _RAND_142 = {1{`RANDOM}};
  _EVAL_946 = _RAND_142[4:0];
  _RAND_143 = {1{`RANDOM}};
  _EVAL_951 = _RAND_143[12:0];
  _RAND_144 = {1{`RANDOM}};
  _EVAL_952 = _RAND_144[2:0];
  _RAND_145 = {1{`RANDOM}};
  _EVAL_954 = _RAND_145[12:0];
  _RAND_146 = {1{`RANDOM}};
  _EVAL_955 = _RAND_146[2:0];
  _RAND_147 = {1{`RANDOM}};
  _EVAL_960 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  _EVAL_971 = _RAND_148[2:0];
  _RAND_149 = {1{`RANDOM}};
  _EVAL_972 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  _EVAL_973 = _RAND_150[2:0];
  _RAND_151 = {1{`RANDOM}};
  _EVAL_976 = _RAND_151[2:0];
  _RAND_152 = {1{`RANDOM}};
  _EVAL_978 = _RAND_152[4:0];
  _RAND_153 = {1{`RANDOM}};
  _EVAL_990 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  _EVAL_993 = _RAND_154[12:0];
  _RAND_155 = {1{`RANDOM}};
  _EVAL_1006 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  _EVAL_1007 = _RAND_156[12:0];
  _RAND_157 = {1{`RANDOM}};
  _EVAL_1010 = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  _EVAL_1012 = _RAND_158[2:0];
  _RAND_159 = {1{`RANDOM}};
  _EVAL_1016 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  _EVAL_1026 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  _EVAL_1030 = _RAND_161[12:0];
  _RAND_162 = {1{`RANDOM}};
  _EVAL_1048 = _RAND_162[12:0];
  _RAND_163 = {1{`RANDOM}};
  _EVAL_1054 = _RAND_163[2:0];
  _RAND_164 = {1{`RANDOM}};
  _EVAL_1055 = _RAND_164[1:0];
  _RAND_165 = {1{`RANDOM}};
  _EVAL_1057 = _RAND_165[12:0];
  _RAND_166 = {1{`RANDOM}};
  _EVAL_1069 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  _EVAL_1078 = _RAND_167[12:0];
  _RAND_168 = {1{`RANDOM}};
  _EVAL_1084 = _RAND_168[2:0];
  _RAND_169 = {1{`RANDOM}};
  _EVAL_1085 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  _EVAL_1093 = _RAND_170[2:0];
  _RAND_171 = {1{`RANDOM}};
  _EVAL_1094 = _RAND_171[2:0];
  _RAND_172 = {1{`RANDOM}};
  _EVAL_1095 = _RAND_172[2:0];
  _RAND_173 = {1{`RANDOM}};
  _EVAL_1101 = _RAND_173[12:0];
  _RAND_174 = {1{`RANDOM}};
  _EVAL_1108 = _RAND_174[12:0];
  _RAND_175 = {1{`RANDOM}};
  _EVAL_1109 = _RAND_175[17:0];
  _RAND_176 = {1{`RANDOM}};
  _EVAL_1119 = _RAND_176[17:0];
  _RAND_177 = {1{`RANDOM}};
  _EVAL_1121 = _RAND_177[12:0];
  _RAND_178 = {1{`RANDOM}};
  _EVAL_1134 = _RAND_178[2:0];
  _RAND_179 = {1{`RANDOM}};
  _EVAL_1138 = _RAND_179[2:0];
  _RAND_180 = {1{`RANDOM}};
  _EVAL_1143 = _RAND_180[12:0];
  _RAND_181 = {1{`RANDOM}};
  _EVAL_1148 = _RAND_181[1:0];
  _RAND_182 = {1{`RANDOM}};
  _EVAL_1160 = _RAND_182[2:0];
  _RAND_183 = {1{`RANDOM}};
  _EVAL_1172 = _RAND_183[2:0];
  _RAND_184 = {1{`RANDOM}};
  _EVAL_1181 = _RAND_184[1:0];
  _RAND_185 = {1{`RANDOM}};
  _EVAL_1193 = _RAND_185[2:0];
  _RAND_186 = {1{`RANDOM}};
  _EVAL_1198 = _RAND_186[2:0];
  _RAND_187 = {1{`RANDOM}};
  _EVAL_1200 = _RAND_187[1:0];
  _RAND_188 = {1{`RANDOM}};
  _EVAL_1203 = _RAND_188[2:0];
  _RAND_189 = {1{`RANDOM}};
  _EVAL_1208 = _RAND_189[2:0];
  _RAND_190 = {1{`RANDOM}};
  _EVAL_1210 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  _EVAL_1211 = _RAND_191[2:0];
  _RAND_192 = {1{`RANDOM}};
  _EVAL_1212 = _RAND_192[12:0];
  _RAND_193 = {1{`RANDOM}};
  _EVAL_1214 = _RAND_193[17:0];
  _RAND_194 = {1{`RANDOM}};
  _EVAL_1220 = _RAND_194[1:0];
  _RAND_195 = {1{`RANDOM}};
  _EVAL_1225 = _RAND_195[1:0];
  _RAND_196 = {1{`RANDOM}};
  _EVAL_1240 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  _EVAL_1241 = _RAND_197[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
