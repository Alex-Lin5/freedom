//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_152_assert(
  input  [2:0] _EVAL,
  input  [1:0] _EVAL_0,
  input        _EVAL_1,
  input        _EVAL_2,
  input  [1:0] _EVAL_3,
  input  [8:0] _EVAL_4,
  input        _EVAL_5,
  input  [2:0] _EVAL_6,
  input        _EVAL_7,
  input        _EVAL_8,
  input        _EVAL_9,
  input        _EVAL_10,
  input        _EVAL_11,
  input        _EVAL_12
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_13;
  wire  _EVAL_14;
  wire  _EVAL_15;
  wire [32:0] _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire [1:0] _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire [1:0] _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire [9:0] _EVAL_51;
  wire  _EVAL_52;
  reg  _EVAL_53;
  wire [1:0] _EVAL_54;
  wire  _EVAL_55;
  reg  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_65;
  wire  _EVAL_66;
  reg [1:0] _EVAL_67;
  wire [1:0] _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  reg [1:0] _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire [1:0] _EVAL_84;
  reg  _EVAL_85;
  wire [1:0] _EVAL_86;
  reg [2:0] _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire [9:0] _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  reg  _EVAL_108;
  wire  _EVAL_109;
  reg  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  reg [8:0] _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  reg  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire [31:0] _EVAL_139;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire [8:0] _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_148;
  reg [2:0] _EVAL_149;
  wire  _EVAL_150;
  wire [9:0] _EVAL_151;
  wire  _EVAL_152;
  reg  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  reg [31:0] _EVAL_161;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_101 = _EVAL_69 | _EVAL_58;
  assign _EVAL_26 = ~_EVAL_17;
  assign _EVAL_59 = _EVAL == 3'h5;
  assign _EVAL_106 = ~_EVAL_157;
  assign _EVAL_41 = ~_EVAL_58;
  assign _EVAL_69 = _EVAL_152 | _EVAL_5;
  assign _EVAL_66 = _EVAL_6 == 3'h4;
  assign _EVAL_30 = _EVAL_56 - 1'h1;
  assign _EVAL_102 = _EVAL_6 == 3'h2;
  assign _EVAL_148 = ~_EVAL_101;
  assign _EVAL_89 = _EVAL_0 != 2'h2;
  assign _EVAL_73 = _EVAL_21 | _EVAL_156;
  assign _EVAL_141 = _EVAL_4 == _EVAL_118;
  assign _EVAL_81 = _EVAL_21 & _EVAL_96;
  assign _EVAL_94 = _EVAL_79 | _EVAL_58;
  assign _EVAL_160 = _EVAL_156 & _EVAL_143;
  assign _EVAL_155 = _EVAL_1 & _EVAL_28;
  assign _EVAL_45 = ~_EVAL_75;
  assign _EVAL_15 = ~_EVAL_133;
  assign _EVAL_159 = _EVAL_55 | _EVAL_58;
  assign _EVAL_82 = _EVAL_12 & _EVAL_70;
  assign _EVAL_98 = _EVAL_21 & _EVAL_97;
  assign _EVAL_52 = ~_EVAL_136;
  assign _EVAL_79 = _EVAL == _EVAL_87;
  assign _EVAL_65 = _EVAL_6 <= 3'h6;
  assign _EVAL_135 = ~_EVAL_74;
  assign _EVAL_44 = _EVAL_126 - 1'h1;
  assign _EVAL_119 = _EVAL_54[0];
  assign _EVAL_39 = _EVAL_3 == _EVAL_80;
  assign _EVAL_46 = ~_EVAL_103;
  assign _EVAL_23 = _EVAL_130 | _EVAL_58;
  assign _EVAL_22 = _EVAL_6 == 3'h0;
  assign _EVAL_33 = _EVAL_12 & _EVAL_22;
  assign _EVAL_38 = _EVAL == 3'h2;
  assign _EVAL_13 = $signed(_EVAL_151) == 10'sh0;
  assign _EVAL_115 = ~_EVAL_146;
  assign _EVAL_132 = _EVAL_1 & _EVAL_129;
  assign _EVAL_105 = ~_EVAL_114;
  assign _EVAL_122 = _EVAL_1 & _EVAL_25;
  assign _EVAL_71 = ~_EVAL_5;
  assign _EVAL_152 = ~_EVAL_11;
  assign _EVAL_84 = _EVAL_98 ? 2'h1 : 2'h0;
  assign _EVAL_25 = _EVAL == 3'h6;
  assign _EVAL_62 = _EVAL_84[0];
  assign _EVAL_75 = _EVAL_92 | _EVAL_58;
  assign _EVAL_70 = _EVAL_6 == 3'h5;
  assign _EVAL_18 = ~_EVAL_145;
  assign _EVAL_86 = _EVAL_123 ? 2'h1 : 2'h0;
  assign _EVAL_131 = _EVAL_60 | _EVAL_58;
  assign _EVAL_130 = _EVAL_124 | _EVAL_109;
  assign _EVAL_37 = _EVAL_152 | _EVAL_58;
  assign _EVAL_128 = _EVAL == 3'h3;
  assign _EVAL_125 = _EVAL_1 & _EVAL_43;
  assign _EVAL_61 = _EVAL_7 == _EVAL_110;
  assign _EVAL_107 = _EVAL_144 == 9'h0;
  assign _EVAL_49 = _EVAL_141 | _EVAL_58;
  assign _EVAL_63 = _EVAL_1 & _EVAL_38;
  assign _EVAL_140 = _EVAL_156 & _EVAL_19;
  assign _EVAL_114 = _EVAL_93 | _EVAL_58;
  assign _EVAL_103 = _EVAL_116 | _EVAL_58;
  assign _EVAL_133 = _EVAL_40 | _EVAL_58;
  assign _EVAL_57 = _EVAL_30[0];
  assign _EVAL_27 = _EVAL == 3'h4;
  assign _EVAL_158 = plusarg_reader_out == 32'h0;
  assign _EVAL_14 = _EVAL_68[0];
  assign _EVAL_55 = _EVAL_3 >= 2'h2;
  assign _EVAL_50 = _EVAL == 3'h1;
  assign _EVAL_19 = ~_EVAL_153;
  assign _EVAL_54 = _EVAL_108 - 1'h1;
  assign _EVAL_116 = ~_EVAL_85;
  assign _EVAL_92 = _EVAL_11 == _EVAL_53;
  assign _EVAL_142 = _EVAL_1 & _EVAL_59;
  assign _EVAL_32 = _EVAL_6 == 3'h6;
  assign _EVAL_90 = _EVAL_12 & _EVAL_112;
  assign _EVAL_99 = {1'b0,$signed(_EVAL_4)};
  assign _EVAL_88 = ~_EVAL_134;
  assign _EVAL_154 = ~_EVAL_76;
  assign _EVAL_48 = _EVAL_1 & _EVAL_50;
  assign _EVAL_31 = _EVAL_12 & _EVAL_32;
  assign _EVAL_156 = _EVAL_9 & _EVAL_12;
  assign _EVAL_36 = ~_EVAL_111;
  assign _EVAL_113 = _EVAL_12 & _EVAL_66;
  assign _EVAL_123 = _EVAL_160 & _EVAL_83;
  assign _EVAL_136 = _EVAL_65 | _EVAL_58;
  assign _EVAL_21 = _EVAL_10 & _EVAL_1;
  assign _EVAL_139 = _EVAL_16[31:0];
  assign _EVAL_104 = ~_EVAL_137;
  assign _EVAL_137 = _EVAL_29 | _EVAL_58;
  assign _EVAL_129 = ~_EVAL_96;
  assign _EVAL_157 = _EVAL_71 | _EVAL_58;
  assign _EVAL_134 = _EVAL_13 | _EVAL_58;
  assign _EVAL_35 = ~_EVAL_94;
  assign _EVAL_112 = ~_EVAL_19;
  assign _EVAL_17 = _EVAL_100 | _EVAL_58;
  assign _EVAL_111 = _EVAL_86[0];
  assign _EVAL_96 = ~_EVAL_108;
  assign _EVAL_97 = ~_EVAL_126;
  assign _EVAL_24 = _EVAL_6 == 3'h1;
  assign _EVAL_29 = _EVAL_0 == _EVAL_67;
  assign _EVAL_91 = _EVAL_85 | _EVAL_62;
  assign _EVAL_77 = ~_EVAL_37;
  assign _EVAL_146 = _EVAL_107 | _EVAL_58;
  assign _EVAL_144 = _EVAL_4 & 9'h3;
  assign _EVAL_109 = _EVAL_161 < plusarg_reader_out;
  assign _EVAL_83 = ~_EVAL_32;
  assign _EVAL_51 = $signed(_EVAL_99) & 10'sh200;
  assign _EVAL_143 = ~_EVAL_56;
  assign _EVAL_93 = _EVAL_0 == 2'h0;
  assign _EVAL_60 = _EVAL_62 | _EVAL_85;
  assign _EVAL_58 = _EVAL_8;
  assign _EVAL_151 = _EVAL_51;
  assign _EVAL_124 = _EVAL_78 | _EVAL_158;
  assign _EVAL_28 = _EVAL == 3'h7;
  assign _EVAL_76 = _EVAL_61 | _EVAL_58;
  assign _EVAL_43 = _EVAL == 3'h0;
  assign _EVAL_74 = _EVAL_89 | _EVAL_58;
  assign _EVAL_72 = _EVAL_12 & _EVAL_24;
  assign _EVAL_68 = _EVAL_153 - 1'h1;
  assign _EVAL_100 = _EVAL_0 <= 2'h2;
  assign _EVAL_120 = ~_EVAL_49;
  assign _EVAL_34 = _EVAL_12 & _EVAL_102;
  assign _EVAL_150 = ~_EVAL_159;
  assign _EVAL_145 = _EVAL_39 | _EVAL_58;
  assign _EVAL_47 = ~_EVAL_131;
  assign _EVAL_78 = ~_EVAL_42;
  assign _EVAL_40 = _EVAL_6 == _EVAL_149;
  assign _EVAL_16 = _EVAL_161 + 32'h1;
  assign _EVAL_121 = _EVAL_1 & _EVAL_27;
  assign _EVAL_20 = _EVAL_1 & _EVAL_128;
  assign _EVAL_127 = _EVAL_44[0];
  assign _EVAL_42 = |_EVAL_85;
  assign _EVAL_138 = ~_EVAL_23;
  always @(posedge _EVAL_2) begin
    if (_EVAL_140) begin
      _EVAL_53 <= _EVAL_11;
    end
    if (_EVAL_140) begin
      _EVAL_67 <= _EVAL_0;
    end
    if (_EVAL_140) begin
      _EVAL_80 <= _EVAL_3;
    end
    if (_EVAL_81) begin
      _EVAL_87 <= _EVAL;
    end
    if (_EVAL_140) begin
      _EVAL_110 <= _EVAL_7;
    end
    if (_EVAL_81) begin
      _EVAL_118 <= _EVAL_4;
    end
    if (_EVAL_140) begin
      _EVAL_149 <= _EVAL_6;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3aee542b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(772f8319)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65775608)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(319ea5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b698dde)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ce31011)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84af9b1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_15) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61c94678)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8721726)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bcbc594)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49893af2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2b445fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1191d07f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5322a7e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26e88d53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_12 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56a24d86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc07e805)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5cbcb7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_46) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4720704)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_120) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9843739b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99edc8b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca3282f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5376508e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da3f8e6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26e80799)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf1a34cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca3282f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d381f3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bed26c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_15) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_45) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30dac7b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_120) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4cf17d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bcdba9bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d90ae2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a124a8ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34c673ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acc2be96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15d10b70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c76862a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c366bc0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_45) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c53019d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fc3371d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_46) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_12 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5ce58c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ab15b30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4207504)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_34 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d780153)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b005627)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da454d4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5598567)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a808db96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_48 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5620dca5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_155 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bee588f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_31 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1caefc3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge _EVAL_2 or posedge _EVAL_8) begin
    if (_EVAL_8) begin
      _EVAL_56 <= 1'h0;
    end else if (_EVAL_156) begin
      if (_EVAL_143) begin
        _EVAL_56 <= 1'h0;
      end else begin
        _EVAL_56 <= _EVAL_57;
      end
    end
  end
  always @(posedge _EVAL_2 or posedge _EVAL_8) begin
    if (_EVAL_8) begin
      _EVAL_85 <= 1'h0;
    end else begin
      _EVAL_85 <= _EVAL_91 & _EVAL_36;
    end
  end
  always @(posedge _EVAL_2 or posedge _EVAL_8) begin
    if (_EVAL_8) begin
      _EVAL_108 <= 1'h0;
    end else if (_EVAL_21) begin
      if (_EVAL_96) begin
        _EVAL_108 <= 1'h0;
      end else begin
        _EVAL_108 <= _EVAL_119;
      end
    end
  end
  always @(posedge _EVAL_2 or posedge _EVAL_8) begin
    if (_EVAL_8) begin
      _EVAL_126 <= 1'h0;
    end else if (_EVAL_21) begin
      if (_EVAL_97) begin
        _EVAL_126 <= 1'h0;
      end else begin
        _EVAL_126 <= _EVAL_127;
      end
    end
  end
  always @(posedge _EVAL_2 or posedge _EVAL_8) begin
    if (_EVAL_8) begin
      _EVAL_153 <= 1'h0;
    end else if (_EVAL_156) begin
      if (_EVAL_19) begin
        _EVAL_153 <= 1'h0;
      end else begin
        _EVAL_153 <= _EVAL_14;
      end
    end
  end
  always @(posedge _EVAL_2 or posedge _EVAL_8) begin
    if (_EVAL_8) begin
      _EVAL_161 <= 32'h0;
    end else if (_EVAL_73) begin
      _EVAL_161 <= 32'h0;
    end else begin
      _EVAL_161 <= _EVAL_139;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_53 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_56 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_67 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_80 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_85 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_87 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_108 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_110 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_118 = _RAND_8[8:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_126 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_149 = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_153 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_161 = _RAND_12[31:0];
`endif // RANDOMIZE_REG_INIT
  if (_EVAL_8) begin
    _EVAL_56 = 1'h0;
  end
  if (_EVAL_8) begin
    _EVAL_85 = 1'h0;
  end
  if (_EVAL_8) begin
    _EVAL_108 = 1'h0;
  end
  if (_EVAL_8) begin
    _EVAL_126 = 1'h0;
  end
  if (_EVAL_8) begin
    _EVAL_153 = 1'h0;
  end
  if (_EVAL_8) begin
    _EVAL_161 = 32'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
