//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_97(
  input  [2:0]   _EVAL,
  input  [2:0]   _EVAL_0,
  input  [2:0]   _EVAL_1,
  input  [2:0]   _EVAL_2,
  input  [2:0]   _EVAL_3,
  input  [2:0]   _EVAL_4,
  input  [2:0]   _EVAL_5,
  input  [2:0]   _EVAL_6,
  input  [2:0]   _EVAL_7,
  input  [2:0]   _EVAL_8,
  input  [2:0]   _EVAL_9,
  input  [2:0]   _EVAL_10,
  input  [2:0]   _EVAL_11,
  input  [2:0]   _EVAL_12,
  input  [2:0]   _EVAL_13,
  input  [2:0]   _EVAL_14,
  input  [2:0]   _EVAL_15,
  input  [2:0]   _EVAL_16,
  input  [2:0]   _EVAL_17,
  input  [2:0]   _EVAL_18,
  input  [2:0]   _EVAL_19,
  input  [2:0]   _EVAL_20,
  input  [2:0]   _EVAL_21,
  input  [2:0]   _EVAL_22,
  input  [2:0]   _EVAL_23,
  input  [2:0]   _EVAL_24,
  input  [2:0]   _EVAL_25,
  input  [2:0]   _EVAL_26,
  input  [2:0]   _EVAL_27,
  input  [2:0]   _EVAL_28,
  input  [2:0]   _EVAL_29,
  input  [2:0]   _EVAL_30,
  input  [2:0]   _EVAL_31,
  input  [2:0]   _EVAL_32,
  input  [2:0]   _EVAL_33,
  input  [2:0]   _EVAL_34,
  input  [2:0]   _EVAL_35,
  input  [2:0]   _EVAL_36,
  input  [2:0]   _EVAL_37,
  input  [2:0]   _EVAL_38,
  input  [2:0]   _EVAL_39,
  input  [2:0]   _EVAL_40,
  input  [2:0]   _EVAL_41,
  input  [2:0]   _EVAL_42,
  input  [2:0]   _EVAL_43,
  input  [2:0]   _EVAL_44,
  input  [2:0]   _EVAL_45,
  input  [2:0]   _EVAL_46,
  input  [2:0]   _EVAL_47,
  input  [126:0] _EVAL_48,
  input  [2:0]   _EVAL_49,
  input  [2:0]   _EVAL_50,
  input  [2:0]   _EVAL_51,
  input  [2:0]   _EVAL_52,
  input  [2:0]   _EVAL_53,
  input  [2:0]   _EVAL_54,
  input  [2:0]   _EVAL_55,
  input  [2:0]   _EVAL_56,
  input  [2:0]   _EVAL_57,
  input  [2:0]   _EVAL_58,
  input  [2:0]   _EVAL_59,
  input  [2:0]   _EVAL_60,
  input  [2:0]   _EVAL_61,
  input  [2:0]   _EVAL_62,
  input  [2:0]   _EVAL_63,
  input  [2:0]   _EVAL_64,
  output [2:0]   _EVAL_65,
  input  [2:0]   _EVAL_66,
  input  [2:0]   _EVAL_67,
  input  [2:0]   _EVAL_68,
  input  [2:0]   _EVAL_69,
  input  [2:0]   _EVAL_70,
  input  [2:0]   _EVAL_71,
  input  [2:0]   _EVAL_72,
  input  [2:0]   _EVAL_73,
  input  [2:0]   _EVAL_74,
  input  [2:0]   _EVAL_75,
  input  [2:0]   _EVAL_76,
  input  [2:0]   _EVAL_77,
  input  [2:0]   _EVAL_78,
  input  [2:0]   _EVAL_79,
  input  [2:0]   _EVAL_80,
  input  [2:0]   _EVAL_81,
  input  [2:0]   _EVAL_82,
  input  [2:0]   _EVAL_83,
  input  [2:0]   _EVAL_84,
  input  [2:0]   _EVAL_85,
  output [6:0]   _EVAL_86,
  input  [2:0]   _EVAL_87,
  input  [2:0]   _EVAL_88,
  input  [2:0]   _EVAL_89,
  input  [2:0]   _EVAL_90,
  input  [2:0]   _EVAL_91,
  input  [2:0]   _EVAL_92,
  input  [2:0]   _EVAL_93,
  input  [2:0]   _EVAL_94,
  input  [2:0]   _EVAL_95,
  input  [2:0]   _EVAL_96,
  input  [2:0]   _EVAL_97,
  input  [2:0]   _EVAL_98,
  input  [2:0]   _EVAL_99,
  input  [2:0]   _EVAL_100,
  input  [2:0]   _EVAL_101,
  input  [2:0]   _EVAL_102,
  input  [2:0]   _EVAL_103,
  input  [2:0]   _EVAL_104,
  input  [2:0]   _EVAL_105,
  input  [2:0]   _EVAL_106,
  input  [2:0]   _EVAL_107,
  input  [2:0]   _EVAL_108,
  input  [2:0]   _EVAL_109,
  input  [2:0]   _EVAL_110,
  input  [2:0]   _EVAL_111,
  input  [2:0]   _EVAL_112,
  input  [2:0]   _EVAL_113,
  input  [2:0]   _EVAL_114,
  input  [2:0]   _EVAL_115,
  input  [2:0]   _EVAL_116,
  input  [2:0]   _EVAL_117,
  input  [2:0]   _EVAL_118,
  input  [2:0]   _EVAL_119,
  input  [2:0]   _EVAL_120,
  input  [2:0]   _EVAL_121,
  input  [2:0]   _EVAL_122,
  input  [2:0]   _EVAL_123,
  input  [2:0]   _EVAL_124,
  input  [2:0]   _EVAL_125,
  input  [2:0]   _EVAL_126,
  input  [2:0]   _EVAL_127,
  input  [2:0]   _EVAL_128
);
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire [1:0] _EVAL_133;
  wire [2:0] _EVAL_134;
  wire [3:0] _EVAL_135;
  wire  _EVAL_136;
  wire [3:0] _EVAL_137;
  wire  _EVAL_138;
  wire [1:0] _EVAL_139;
  wire  _EVAL_140;
  wire [1:0] _EVAL_141;
  wire [2:0] _EVAL_142;
  wire  _EVAL_143;
  wire [3:0] _EVAL_144;
  wire [3:0] _EVAL_145;
  wire [4:0] _EVAL_146;
  wire [2:0] _EVAL_147;
  wire  _EVAL_148;
  wire [3:0] _EVAL_149;
  wire [2:0] _EVAL_150;
  wire [3:0] _EVAL_151;
  wire [3:0] _EVAL_152;
  wire  _EVAL_153;
  wire [3:0] _EVAL_154;
  wire [1:0] _EVAL_155;
  wire [3:0] _EVAL_156;
  wire  _EVAL_157;
  wire [3:0] _EVAL_158;
  wire [1:0] _EVAL_159;
  wire [1:0] _EVAL_160;
  wire  _EVAL_161;
  wire [3:0] _EVAL_162;
  wire [2:0] _EVAL_163;
  wire [3:0] _EVAL_164;
  wire  _EVAL_165;
  wire [3:0] _EVAL_166;
  wire [1:0] _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire [3:0] _EVAL_170;
  wire [1:0] _EVAL_171;
  wire [3:0] _EVAL_172;
  wire  _EVAL_173;
  wire [3:0] _EVAL_174;
  wire [1:0] _EVAL_175;
  wire [3:0] _EVAL_176;
  wire [3:0] _EVAL_177;
  wire [1:0] _EVAL_178;
  wire [1:0] _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire [2:0] _EVAL_182;
  wire  _EVAL_183;
  wire [2:0] _EVAL_184;
  wire [3:0] _EVAL_185;
  wire [3:0] _EVAL_186;
  wire [3:0] _EVAL_187;
  wire  _EVAL_188;
  wire [3:0] _EVAL_189;
  wire [3:0] _EVAL_190;
  wire [1:0] _EVAL_191;
  wire [3:0] _EVAL_192;
  wire [3:0] _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire [1:0] _EVAL_196;
  wire  _EVAL_197;
  wire [1:0] _EVAL_198;
  wire  _EVAL_199;
  wire [3:0] _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire [3:0] _EVAL_206;
  wire  _EVAL_207;
  wire [1:0] _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire [1:0] _EVAL_211;
  wire [3:0] _EVAL_212;
  wire [3:0] _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire [3:0] _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire [3:0] _EVAL_219;
  wire [3:0] _EVAL_220;
  wire  _EVAL_221;
  wire [2:0] _EVAL_222;
  wire  _EVAL_223;
  wire [1:0] _EVAL_224;
  wire  _EVAL_225;
  wire [3:0] _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire [1:0] _EVAL_229;
  wire [3:0] _EVAL_230;
  wire  _EVAL_231;
  wire [3:0] _EVAL_232;
  wire [4:0] _EVAL_233;
  wire [3:0] _EVAL_234;
  wire  _EVAL_235;
  wire [3:0] _EVAL_236;
  wire [3:0] _EVAL_237;
  wire  _EVAL_238;
  wire [3:0] _EVAL_239;
  wire  _EVAL_240;
  wire [2:0] _EVAL_241;
  wire [3:0] _EVAL_242;
  wire  _EVAL_243;
  wire [3:0] _EVAL_244;
  wire [2:0] _EVAL_245;
  wire  _EVAL_246;
  wire [3:0] _EVAL_247;
  wire [3:0] _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire [3:0] _EVAL_251;
  wire [3:0] _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire [3:0] _EVAL_257;
  wire  _EVAL_258;
  wire [3:0] _EVAL_259;
  wire [2:0] _EVAL_260;
  wire  _EVAL_261;
  wire [2:0] _EVAL_262;
  wire [3:0] _EVAL_263;
  wire  _EVAL_264;
  wire [3:0] _EVAL_265;
  wire [3:0] _EVAL_266;
  wire  _EVAL_267;
  wire [3:0] _EVAL_268;
  wire [3:0] _EVAL_269;
  wire  _EVAL_270;
  wire [3:0] _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire [3:0] _EVAL_274;
  wire [3:0] _EVAL_275;
  wire [3:0] _EVAL_276;
  wire [2:0] _EVAL_277;
  wire [3:0] _EVAL_278;
  wire  _EVAL_279;
  wire  _EVAL_280;
  wire [3:0] _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire [3:0] _EVAL_289;
  wire [1:0] _EVAL_290;
  wire [3:0] _EVAL_291;
  wire [3:0] _EVAL_292;
  wire [3:0] _EVAL_293;
  wire [3:0] _EVAL_294;
  wire [4:0] _EVAL_295;
  wire [3:0] _EVAL_296;
  wire  _EVAL_297;
  wire  _EVAL_298;
  wire [3:0] _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_302;
  wire [3:0] _EVAL_303;
  wire  _EVAL_304;
  wire [1:0] _EVAL_305;
  wire [3:0] _EVAL_306;
  wire  _EVAL_307;
  wire  _EVAL_308;
  wire  _EVAL_309;
  wire [5:0] _EVAL_310;
  wire  _EVAL_311;
  wire [1:0] _EVAL_312;
  wire [3:0] _EVAL_313;
  wire [3:0] _EVAL_314;
  wire [2:0] _EVAL_315;
  wire [3:0] _EVAL_316;
  wire [3:0] _EVAL_317;
  wire  _EVAL_318;
  wire [2:0] _EVAL_319;
  wire [3:0] _EVAL_320;
  wire [1:0] _EVAL_321;
  wire [1:0] _EVAL_322;
  wire [1:0] _EVAL_323;
  wire  _EVAL_324;
  wire [1:0] _EVAL_325;
  wire [3:0] _EVAL_326;
  wire  _EVAL_327;
  wire  _EVAL_328;
  wire [3:0] _EVAL_329;
  wire [3:0] _EVAL_330;
  wire [2:0] _EVAL_331;
  wire [3:0] _EVAL_332;
  wire [3:0] _EVAL_333;
  wire  _EVAL_334;
  wire  _EVAL_335;
  wire [3:0] _EVAL_336;
  wire [3:0] _EVAL_337;
  wire [2:0] _EVAL_338;
  wire  _EVAL_339;
  wire  _EVAL_340;
  wire [1:0] _EVAL_341;
  wire [3:0] _EVAL_342;
  wire  _EVAL_343;
  wire [3:0] _EVAL_344;
  wire [3:0] _EVAL_345;
  wire [3:0] _EVAL_346;
  wire [3:0] _EVAL_347;
  wire [3:0] _EVAL_348;
  wire [1:0] _EVAL_349;
  wire [3:0] _EVAL_350;
  wire  _EVAL_351;
  wire [2:0] _EVAL_352;
  wire [6:0] _EVAL_353;
  wire  _EVAL_354;
  wire [1:0] _EVAL_355;
  wire [3:0] _EVAL_356;
  wire  _EVAL_357;
  wire  _EVAL_358;
  wire  _EVAL_359;
  wire [1:0] _EVAL_360;
  wire  _EVAL_361;
  wire [1:0] _EVAL_362;
  wire [3:0] _EVAL_363;
  wire  _EVAL_364;
  wire  _EVAL_365;
  wire  _EVAL_366;
  wire  _EVAL_367;
  wire [1:0] _EVAL_368;
  wire  _EVAL_369;
  wire [3:0] _EVAL_370;
  wire [3:0] _EVAL_371;
  wire  _EVAL_372;
  wire [3:0] _EVAL_373;
  wire  _EVAL_374;
  wire  _EVAL_375;
  wire  _EVAL_376;
  wire  _EVAL_377;
  wire  _EVAL_378;
  wire [3:0] _EVAL_379;
  wire [3:0] _EVAL_380;
  wire  _EVAL_381;
  wire [3:0] _EVAL_382;
  wire [3:0] _EVAL_383;
  wire [3:0] _EVAL_384;
  wire  _EVAL_385;
  wire [3:0] _EVAL_386;
  wire [3:0] _EVAL_387;
  wire  _EVAL_388;
  wire  _EVAL_389;
  wire  _EVAL_390;
  wire [3:0] _EVAL_391;
  wire [3:0] _EVAL_392;
  wire  _EVAL_393;
  wire [3:0] _EVAL_394;
  wire  _EVAL_395;
  wire  _EVAL_396;
  wire [1:0] _EVAL_397;
  wire [1:0] _EVAL_398;
  wire [3:0] _EVAL_399;
  wire  _EVAL_400;
  wire [3:0] _EVAL_401;
  wire  _EVAL_402;
  wire [3:0] _EVAL_403;
  wire  _EVAL_404;
  wire  _EVAL_405;
  wire [3:0] _EVAL_406;
  wire [2:0] _EVAL_407;
  wire  _EVAL_408;
  wire [3:0] _EVAL_409;
  wire  _EVAL_410;
  wire [1:0] _EVAL_411;
  wire [3:0] _EVAL_412;
  wire [3:0] _EVAL_413;
  wire [2:0] _EVAL_414;
  wire [3:0] _EVAL_415;
  wire [3:0] _EVAL_416;
  wire [5:0] _EVAL_417;
  wire [3:0] _EVAL_418;
  wire  _EVAL_419;
  wire [3:0] _EVAL_420;
  wire [3:0] _EVAL_421;
  wire [3:0] _EVAL_422;
  wire  _EVAL_423;
  wire [1:0] _EVAL_424;
  wire [3:0] _EVAL_425;
  wire [1:0] _EVAL_426;
  wire  _EVAL_427;
  wire  _EVAL_428;
  wire  _EVAL_429;
  wire  _EVAL_430;
  wire [3:0] _EVAL_431;
  wire  _EVAL_432;
  wire [3:0] _EVAL_433;
  wire  _EVAL_434;
  wire [3:0] _EVAL_435;
  wire [3:0] _EVAL_436;
  wire [1:0] _EVAL_437;
  wire  _EVAL_438;
  wire  _EVAL_439;
  wire [3:0] _EVAL_440;
  wire [3:0] _EVAL_441;
  wire  _EVAL_442;
  wire [2:0] _EVAL_443;
  wire  _EVAL_444;
  wire  _EVAL_445;
  wire [2:0] _EVAL_446;
  wire  _EVAL_447;
  wire  _EVAL_448;
  wire  _EVAL_449;
  wire [3:0] _EVAL_450;
  wire [3:0] _EVAL_451;
  wire [3:0] _EVAL_452;
  wire  _EVAL_453;
  wire [1:0] _EVAL_454;
  wire  _EVAL_455;
  wire [2:0] _EVAL_456;
  wire [2:0] _EVAL_457;
  wire [3:0] _EVAL_458;
  wire  _EVAL_459;
  wire  _EVAL_460;
  wire [3:0] _EVAL_461;
  wire  _EVAL_462;
  wire  _EVAL_463;
  wire [3:0] _EVAL_464;
  wire  _EVAL_465;
  wire  _EVAL_466;
  wire  _EVAL_467;
  wire [1:0] _EVAL_468;
  wire  _EVAL_469;
  wire  _EVAL_470;
  wire  _EVAL_471;
  wire  _EVAL_472;
  wire [3:0] _EVAL_473;
  wire [1:0] _EVAL_474;
  wire [3:0] _EVAL_475;
  wire [3:0] _EVAL_476;
  wire [1:0] _EVAL_477;
  wire  _EVAL_478;
  wire [1:0] _EVAL_479;
  wire  _EVAL_480;
  wire  _EVAL_481;
  wire [3:0] _EVAL_482;
  wire [3:0] _EVAL_483;
  wire [1:0] _EVAL_484;
  wire [3:0] _EVAL_485;
  wire [1:0] _EVAL_486;
  wire [3:0] _EVAL_487;
  wire [1:0] _EVAL_488;
  wire  _EVAL_489;
  wire  _EVAL_490;
  wire  _EVAL_491;
  wire  _EVAL_492;
  wire  _EVAL_493;
  wire [3:0] _EVAL_494;
  wire [3:0] _EVAL_495;
  wire  _EVAL_496;
  wire [3:0] _EVAL_497;
  wire  _EVAL_498;
  wire [2:0] _EVAL_499;
  wire [3:0] _EVAL_500;
  wire [3:0] _EVAL_501;
  wire [4:0] _EVAL_502;
  wire  _EVAL_503;
  wire  _EVAL_504;
  wire [3:0] _EVAL_505;
  wire [3:0] _EVAL_506;
  wire  _EVAL_507;
  wire [3:0] _EVAL_508;
  wire [3:0] _EVAL_509;
  wire  _EVAL_510;
  wire  _EVAL_511;
  wire [3:0] _EVAL_512;
  wire  _EVAL_513;
  wire  _EVAL_514;
  wire  _EVAL_515;
  wire  _EVAL_516;
  wire  _EVAL_517;
  wire  _EVAL_518;
  wire  _EVAL_519;
  wire  _EVAL_520;
  wire [1:0] _EVAL_521;
  wire [3:0] _EVAL_522;
  wire  _EVAL_523;
  wire  _EVAL_524;
  wire [3:0] _EVAL_525;
  wire  _EVAL_526;
  wire [3:0] _EVAL_527;
  wire [3:0] _EVAL_528;
  wire [3:0] _EVAL_529;
  wire [3:0] _EVAL_530;
  wire  _EVAL_531;
  wire [3:0] _EVAL_532;
  wire  _EVAL_533;
  wire  _EVAL_534;
  wire  _EVAL_535;
  wire [3:0] _EVAL_536;
  wire [1:0] _EVAL_537;
  wire [3:0] _EVAL_538;
  wire  _EVAL_539;
  wire [3:0] _EVAL_540;
  wire  _EVAL_541;
  wire [3:0] _EVAL_542;
  wire [3:0] _EVAL_543;
  wire [3:0] _EVAL_544;
  wire  _EVAL_545;
  wire [3:0] _EVAL_546;
  wire  _EVAL_547;
  wire  _EVAL_548;
  wire [1:0] _EVAL_549;
  wire  _EVAL_550;
  wire [2:0] _EVAL_551;
  wire [3:0] _EVAL_552;
  wire [3:0] _EVAL_553;
  wire [1:0] _EVAL_554;
  wire [3:0] _EVAL_555;
  wire  _EVAL_556;
  wire [3:0] _EVAL_557;
  wire  _EVAL_558;
  wire  _EVAL_559;
  wire [3:0] _EVAL_560;
  wire [3:0] _EVAL_561;
  wire [3:0] _EVAL_562;
  wire [3:0] _EVAL_563;
  wire  _EVAL_564;
  wire  _EVAL_565;
  wire [3:0] _EVAL_566;
  wire [3:0] _EVAL_567;
  wire  _EVAL_568;
  wire [2:0] _EVAL_569;
  wire  _EVAL_570;
  wire [1:0] _EVAL_571;
  wire [3:0] _EVAL_572;
  wire [3:0] _EVAL_573;
  wire  _EVAL_574;
  wire  _EVAL_575;
  wire [3:0] _EVAL_576;
  wire [2:0] _EVAL_577;
  wire [3:0] _EVAL_578;
  wire  _EVAL_579;
  wire [1:0] _EVAL_580;
  wire [6:0] _EVAL_581;
  wire [3:0] _EVAL_582;
  wire [3:0] _EVAL_583;
  wire [3:0] _EVAL_584;
  wire  _EVAL_585;
  wire [4:0] _EVAL_586;
  wire [2:0] _EVAL_587;
  wire  _EVAL_588;
  wire [3:0] _EVAL_589;
  wire [3:0] _EVAL_590;
  wire [1:0] _EVAL_591;
  wire [3:0] _EVAL_592;
  wire [3:0] _EVAL_593;
  wire [1:0] _EVAL_594;
  wire [3:0] _EVAL_595;
  wire [3:0] _EVAL_596;
  wire [3:0] _EVAL_597;
  wire [3:0] _EVAL_598;
  wire [1:0] _EVAL_599;
  wire  _EVAL_600;
  wire [3:0] _EVAL_601;
  wire [4:0] _EVAL_602;
  wire  _EVAL_603;
  wire  _EVAL_604;
  wire [2:0] _EVAL_605;
  wire [3:0] _EVAL_606;
  wire  _EVAL_607;
  wire [4:0] _EVAL_608;
  wire  _EVAL_609;
  wire  _EVAL_610;
  wire [3:0] _EVAL_611;
  wire [3:0] _EVAL_612;
  wire [3:0] _EVAL_613;
  wire  _EVAL_614;
  wire [1:0] _EVAL_615;
  wire [3:0] _EVAL_616;
  wire [1:0] _EVAL_617;
  wire  _EVAL_618;
  wire [3:0] _EVAL_619;
  wire [3:0] _EVAL_620;
  wire  _EVAL_621;
  wire  _EVAL_622;
  wire  _EVAL_623;
  wire [1:0] _EVAL_624;
  wire  _EVAL_625;
  wire  _EVAL_626;
  wire  _EVAL_627;
  wire [1:0] _EVAL_628;
  wire [3:0] _EVAL_629;
  wire [3:0] _EVAL_630;
  wire [3:0] _EVAL_631;
  wire [3:0] _EVAL_632;
  wire [3:0] _EVAL_633;
  wire  _EVAL_634;
  wire [3:0] _EVAL_635;
  wire  _EVAL_636;
  wire  _EVAL_637;
  wire  _EVAL_638;
  wire [3:0] _EVAL_639;
  wire  _EVAL_640;
  wire [1:0] _EVAL_641;
  wire  _EVAL_642;
  wire  _EVAL_643;
  wire  _EVAL_644;
  wire [2:0] _EVAL_645;
  wire [3:0] _EVAL_646;
  wire [3:0] _EVAL_647;
  wire [3:0] _EVAL_648;
  wire [1:0] _EVAL_649;
  wire  _EVAL_650;
  wire  _EVAL_651;
  wire [3:0] _EVAL_652;
  wire  _EVAL_653;
  wire [3:0] _EVAL_654;
  wire [1:0] _EVAL_655;
  wire  _EVAL_656;
  wire [1:0] _EVAL_657;
  wire  _EVAL_658;
  wire [3:0] _EVAL_659;
  wire [3:0] _EVAL_660;
  wire [1:0] _EVAL_661;
  wire  _EVAL_662;
  wire [2:0] _EVAL_663;
  wire  _EVAL_664;
  wire  _EVAL_665;
  wire  _EVAL_666;
  wire [1:0] _EVAL_667;
  wire  _EVAL_668;
  wire [3:0] _EVAL_669;
  wire [4:0] _EVAL_670;
  wire [2:0] _EVAL_671;
  wire [3:0] _EVAL_672;
  wire [3:0] _EVAL_673;
  wire [3:0] _EVAL_674;
  wire [3:0] _EVAL_675;
  wire [1:0] _EVAL_676;
  wire [3:0] _EVAL_677;
  wire [3:0] _EVAL_678;
  wire [3:0] _EVAL_679;
  wire [3:0] _EVAL_680;
  wire  _EVAL_681;
  wire  _EVAL_682;
  wire  _EVAL_683;
  wire [3:0] _EVAL_684;
  wire [4:0] _EVAL_685;
  wire  _EVAL_686;
  wire  _EVAL_687;
  wire  _EVAL_688;
  wire  _EVAL_689;
  wire [4:0] _EVAL_690;
  wire  _EVAL_691;
  wire [3:0] _EVAL_692;
  wire  _EVAL_693;
  wire  _EVAL_694;
  wire [2:0] _EVAL_695;
  wire  _EVAL_696;
  wire [5:0] _EVAL_697;
  wire  _EVAL_698;
  wire [3:0] _EVAL_699;
  wire [3:0] _EVAL_700;
  wire  _EVAL_701;
  wire  _EVAL_702;
  wire [3:0] _EVAL_703;
  wire [3:0] _EVAL_704;
  wire  _EVAL_705;
  wire [2:0] _EVAL_706;
  wire [3:0] _EVAL_707;
  wire  _EVAL_708;
  wire [3:0] _EVAL_709;
  wire [1:0] _EVAL_710;
  wire [3:0] _EVAL_711;
  wire [3:0] _EVAL_712;
  wire [3:0] _EVAL_713;
  wire [2:0] _EVAL_714;
  wire  _EVAL_715;
  wire  _EVAL_716;
  wire [3:0] _EVAL_717;
  wire [1:0] _EVAL_718;
  wire  _EVAL_719;
  wire [3:0] _EVAL_720;
  wire [3:0] _EVAL_721;
  wire  _EVAL_722;
  wire  _EVAL_723;
  wire [3:0] _EVAL_724;
  wire  _EVAL_725;
  wire  _EVAL_726;
  wire [2:0] _EVAL_727;
  wire [3:0] _EVAL_728;
  wire [1:0] _EVAL_729;
  wire [4:0] _EVAL_730;
  wire [2:0] _EVAL_731;
  wire  _EVAL_732;
  wire [3:0] _EVAL_733;
  wire [1:0] _EVAL_734;
  wire [1:0] _EVAL_735;
  wire  _EVAL_736;
  wire  _EVAL_737;
  wire [3:0] _EVAL_738;
  wire [3:0] _EVAL_739;
  wire  _EVAL_740;
  wire  _EVAL_741;
  wire  _EVAL_742;
  wire [3:0] _EVAL_743;
  wire [2:0] _EVAL_744;
  wire [1:0] _EVAL_745;
  wire  _EVAL_746;
  wire  _EVAL_747;
  wire  _EVAL_748;
  wire [5:0] _EVAL_749;
  wire [3:0] _EVAL_750;
  wire  _EVAL_751;
  wire [1:0] _EVAL_752;
  wire  _EVAL_753;
  wire [3:0] _EVAL_754;
  wire  _EVAL_755;
  wire  _EVAL_756;
  wire [3:0] _EVAL_757;
  wire  _EVAL_758;
  wire  _EVAL_759;
  wire [3:0] _EVAL_760;
  wire [1:0] _EVAL_761;
  wire [3:0] _EVAL_762;
  wire  _EVAL_763;
  wire  _EVAL_764;
  wire [2:0] _EVAL_765;
  wire [3:0] _EVAL_766;
  wire [1:0] _EVAL_767;
  wire [3:0] _EVAL_768;
  wire [1:0] _EVAL_769;
  wire [3:0] _EVAL_770;
  wire [3:0] _EVAL_771;
  wire [3:0] _EVAL_772;
  wire  _EVAL_773;
  wire [2:0] _EVAL_774;
  wire [2:0] _EVAL_775;
  wire  _EVAL_776;
  wire [1:0] _EVAL_777;
  wire  _EVAL_778;
  wire [3:0] _EVAL_779;
  wire [3:0] _EVAL_780;
  wire  _EVAL_781;
  wire  _EVAL_782;
  wire  _EVAL_783;
  wire [3:0] _EVAL_784;
  wire [1:0] _EVAL_785;
  wire [3:0] _EVAL_786;
  wire  _EVAL_787;
  wire  _EVAL_788;
  wire [1:0] _EVAL_789;
  wire  _EVAL_790;
  wire  _EVAL_791;
  wire  _EVAL_792;
  wire [3:0] _EVAL_793;
  wire [3:0] _EVAL_794;
  wire  _EVAL_795;
  wire [3:0] _EVAL_796;
  wire [3:0] _EVAL_797;
  wire  _EVAL_798;
  wire  _EVAL_799;
  wire  _EVAL_800;
  wire [1:0] _EVAL_801;
  wire [3:0] _EVAL_802;
  wire  _EVAL_803;
  wire  _EVAL_804;
  wire [5:0] _EVAL_805;
  wire [3:0] _EVAL_806;
  wire [3:0] _EVAL_807;
  wire  _EVAL_808;
  wire [1:0] _EVAL_809;
  wire [3:0] _EVAL_810;
  wire [1:0] _EVAL_811;
  wire  _EVAL_812;
  wire [3:0] _EVAL_813;
  wire [2:0] _EVAL_814;
  wire [3:0] _EVAL_815;
  wire  _EVAL_816;
  wire  _EVAL_817;
  wire  _EVAL_818;
  wire [1:0] _EVAL_819;
  wire [1:0] _EVAL_820;
  wire [1:0] _EVAL_821;
  wire [3:0] _EVAL_822;
  wire [2:0] _EVAL_823;
  wire  _EVAL_824;
  wire [3:0] _EVAL_825;
  wire [4:0] _EVAL_826;
  wire [3:0] _EVAL_827;
  wire [1:0] _EVAL_828;
  wire [3:0] _EVAL_829;
  wire  _EVAL_830;
  wire  _EVAL_831;
  wire [1:0] _EVAL_832;
  wire  _EVAL_833;
  wire  _EVAL_834;
  wire [3:0] _EVAL_835;
  wire  _EVAL_836;
  wire [3:0] _EVAL_837;
  wire [3:0] _EVAL_838;
  wire  _EVAL_839;
  wire [5:0] _EVAL_840;
  wire  _EVAL_841;
  wire  _EVAL_842;
  wire [2:0] _EVAL_843;
  wire [2:0] _EVAL_844;
  wire  _EVAL_845;
  wire [3:0] _EVAL_846;
  wire  _EVAL_847;
  wire [3:0] _EVAL_848;
  wire  _EVAL_849;
  wire [3:0] _EVAL_850;
  wire  _EVAL_851;
  wire [1:0] _EVAL_852;
  wire [2:0] _EVAL_853;
  wire [1:0] _EVAL_854;
  wire [3:0] _EVAL_855;
  wire [1:0] _EVAL_856;
  wire  _EVAL_857;
  wire  _EVAL_858;
  wire  _EVAL_859;
  wire  _EVAL_860;
  wire [3:0] _EVAL_861;
  wire [1:0] _EVAL_862;
  wire  _EVAL_863;
  wire [3:0] _EVAL_864;
  wire  _EVAL_865;
  wire [1:0] _EVAL_866;
  wire  _EVAL_867;
  wire [3:0] _EVAL_868;
  wire [3:0] _EVAL_869;
  wire [3:0] _EVAL_870;
  wire  _EVAL_871;
  wire [3:0] _EVAL_872;
  wire [3:0] _EVAL_873;
  wire [2:0] _EVAL_874;
  wire  _EVAL_875;
  wire [1:0] _EVAL_876;
  wire  _EVAL_877;
  wire  _EVAL_878;
  wire  _EVAL_879;
  wire [1:0] _EVAL_880;
  wire [1:0] _EVAL_881;
  wire  _EVAL_882;
  wire  _EVAL_883;
  wire [3:0] _EVAL_884;
  wire [3:0] _EVAL_885;
  wire [1:0] _EVAL_886;
  wire  _EVAL_887;
  wire [1:0] _EVAL_888;
  assign _EVAL_610 = _EVAL_552 >= _EVAL_252;
  assign _EVAL_828 = 2'h2 | _EVAL_167;
  assign _EVAL_443 = 3'h4 | _EVAL_457;
  assign _EVAL_731 = _EVAL_453 ? {{1'd0}, _EVAL_323} : _EVAL_260;
  assign _EVAL_396 = _EVAL_48[96];
  assign _EVAL_608 = 5'h10 | _EVAL_730;
  assign _EVAL_215 = _EVAL_48[100];
  assign _EVAL_870 = _EVAL_834 ? _EVAL_348 : _EVAL_156;
  assign _EVAL_746 = _EVAL_565 ? 1'h0 : 1'h1;
  assign _EVAL_770 = {_EVAL_169,_EVAL_82};
  assign _EVAL_862 = {{1'd0}, _EVAL_419};
  assign _EVAL_478 = _EVAL_219 >= _EVAL_613;
  assign _EVAL_194 = _EVAL_48[55];
  assign _EVAL_884 = _EVAL_860 ? _EVAL_299 : _EVAL_717;
  assign _EVAL_511 = _EVAL_48[15];
  assign _EVAL_344 = _EVAL_808 ? _EVAL_170 : _EVAL_546;
  assign _EVAL_618 = _EVAL_48[74];
  assign _EVAL_570 = _EVAL_772 >= _EVAL_700;
  assign _EVAL_562 = {_EVAL_194,_EVAL_28};
  assign _EVAL_831 = _EVAL_48[11];
  assign _EVAL_773 = _EVAL_791 ? 1'h0 : 1'h1;
  assign _EVAL_188 = _EVAL_209 ? 1'h0 : 1'h1;
  assign _EVAL_813 = _EVAL_791 ? _EVAL_306 : _EVAL_869;
  assign _EVAL_277 = {{1'd0}, _EVAL_655};
  assign _EVAL_665 = _EVAL_183 ? 1'h0 : 1'h1;
  assign _EVAL_819 = _EVAL_287 ? {{1'd0}, _EVAL_254} : _EVAL_752;
  assign _EVAL_168 = _EVAL_458 >= _EVAL_596;
  assign _EVAL_630 = _EVAL_439 ? _EVAL_149 : _EVAL_601;
  assign _EVAL_399 = _EVAL_328 ? _EVAL_873 : _EVAL_380;
  assign _EVAL_304 = _EVAL_309 ? 1'h0 : 1'h1;
  assign _EVAL_325 = _EVAL_781 ? {{1'd0}, _EVAL_725} : _EVAL_628;
  assign _EVAL_181 = _EVAL_48[2];
  assign _EVAL_431 = _EVAL_664 ? _EVAL_291 : _EVAL_743;
  assign _EVAL_416 = {_EVAL_668,_EVAL_78};
  assign _EVAL_609 = _EVAL_415 >= _EVAL_172;
  assign _EVAL_827 = _EVAL_301 ? _EVAL_669 : _EVAL_475;
  assign _EVAL_711 = {_EVAL_221,_EVAL_54};
  assign _EVAL_303 = _EVAL_503 ? _EVAL_332 : _EVAL_584;
  assign _EVAL_232 = {_EVAL_541,_EVAL_75};
  assign _EVAL_499 = {{1'd0}, _EVAL_139};
  assign _EVAL_650 = _EVAL_771 >= _EVAL_576;
  assign _EVAL_823 = _EVAL_642 ? {{1'd0}, _EVAL_819} : _EVAL_765;
  assign _EVAL_354 = _EVAL_48[122];
  assign _EVAL_754 = _EVAL_153 ? _EVAL_677 : _EVAL_144;
  assign _EVAL_509 = _EVAL_753 ? _EVAL_363 : _EVAL_174;
  assign _EVAL_153 = _EVAL_677 >= _EVAL_144;
  assign _EVAL_662 = _EVAL_48[116];
  assign _EVAL_702 = _EVAL_712 >= _EVAL_870;
  assign _EVAL_655 = _EVAL_478 ? {{1'd0}, _EVAL_430} : _EVAL_777;
  assign _EVAL_493 = _EVAL_48[25];
  assign _EVAL_193 = _EVAL_588 ? _EVAL_673 : _EVAL_561;
  assign _EVAL_768 = {_EVAL_143,_EVAL_47};
  assign _EVAL_784 = _EVAL_535 ? _EVAL_418 : _EVAL_582;
  assign _EVAL_406 = {_EVAL_335,_EVAL_16};
  assign _EVAL_379 = _EVAL_517 ? _EVAL_425 : _EVAL_837;
  assign _EVAL_680 = _EVAL_309 ? _EVAL_786 : _EVAL_185;
  assign _EVAL_220 = 4'h8 | _EVAL_612;
  assign _EVAL_174 = {_EVAL_459,_EVAL_51};
  assign _EVAL_439 = _EVAL_149 >= _EVAL_601;
  assign _EVAL_262 = 3'h4 | _EVAL_744;
  assign _EVAL_540 = {{1'd0}, _EVAL_338};
  assign _EVAL_826 = 5'h10 | _EVAL_685;
  assign _EVAL_204 = _EVAL_48[23];
  assign _EVAL_410 = _EVAL_48[77];
  assign _EVAL_480 = _EVAL_472 ? 1'h0 : 1'h1;
  assign _EVAL_872 = _EVAL_250 ? _EVAL_536 : _EVAL_450;
  assign _EVAL_138 = _EVAL_48[58];
  assign _EVAL_834 = _EVAL_348 >= _EVAL_156;
  assign _EVAL_375 = _EVAL_719 ? 1'h0 : 1'h1;
  assign _EVAL_157 = _EVAL_48[42];
  assign _EVAL_863 = _EVAL_48[115];
  assign _EVAL_700 = {_EVAL_215,_EVAL_34};
  assign _EVAL_677 = _EVAL_559 ? _EVAL_797 : _EVAL_553;
  assign _EVAL_865 = _EVAL_542 >= _EVAL_784;
  assign _EVAL_625 = _EVAL_609 ? 1'h0 : 1'h1;
  assign _EVAL_217 = _EVAL_48[85];
  assign _EVAL_218 = _EVAL_787 ? 1'h0 : 1'h1;
  assign _EVAL_704 = {_EVAL_547,_EVAL_115};
  assign _EVAL_286 = _EVAL_137 >= _EVAL_409;
  assign _EVAL_852 = _EVAL_231 ? {{1'd0}, _EVAL_847} : _EVAL_866;
  assign _EVAL_383 = {_EVAL_716,_EVAL_9};
  assign _EVAL_460 = _EVAL_465 ? 1'h0 : 1'h1;
  assign _EVAL_750 = _EVAL_183 ? _EVAL_281 : _EVAL_835;
  assign _EVAL_191 = {{1'd0}, _EVAL_201};
  assign _EVAL_645 = 3'h4 | _EVAL_315;
  assign _EVAL_718 = {{1'd0}, _EVAL_188};
  assign _EVAL_613 = _EVAL_209 ? _EVAL_672 : _EVAL_850;
  assign _EVAL_874 = _EVAL_286 ? {{1'd0}, _EVAL_571} : _EVAL_645;
  assign _EVAL_239 = {_EVAL_818,_EVAL_83};
  assign _EVAL_295 = {{1'd0}, _EVAL_382};
  assign _EVAL_362 = {{1'd0}, _EVAL_471};
  assign _EVAL_559 = _EVAL_797 >= _EVAL_553;
  assign _EVAL_600 = _EVAL_48[91];
  assign _EVAL_708 = _EVAL_742 ? 1'h0 : 1'h1;
  assign _EVAL_781 = _EVAL_399 >= _EVAL_794;
  assign _EVAL_771 = _EVAL_203 ? _EVAL_370 : _EVAL_757;
  assign _EVAL_684 = {{1'd0}, _EVAL_456};
  assign _EVAL_735 = 2'h2 | _EVAL_398;
  assign _EVAL_261 = _EVAL_506 >= _EVAL_512;
  assign _EVAL_149 = _EVAL_327 ? _EVAL_709 : _EVAL_838;
  assign _EVAL_709 = {_EVAL_621,_EVAL_58};
  assign _EVAL_134 = _EVAL_882 ? {{1'd0}, _EVAL_854} : _EVAL_695;
  assign _EVAL_679 = {_EVAL_687,_EVAL_1};
  assign _EVAL_347 = _EVAL_199 ? {{1'd0}, _EVAL_446} : _EVAL_675;
  assign _EVAL_550 = _EVAL_544 >= _EVAL_431;
  assign _EVAL_359 = _EVAL_483 >= _EVAL_441;
  assign _EVAL_585 = _EVAL_337 >= _EVAL_316;
  assign _EVAL_748 = _EVAL_48[103];
  assign _EVAL_421 = {_EVAL_228,_EVAL_21};
  assign _EVAL_534 = _EVAL_48[27];
  assign _EVAL_794 = _EVAL_609 ? _EVAL_415 : _EVAL_172;
  assign _EVAL_411 = {{1'd0}, _EVAL_449};
  assign _EVAL_454 = _EVAL_664 ? {{1'd0}, _EVAL_607} : _EVAL_171;
  assign _EVAL_206 = {_EVAL_531,_EVAL_113};
  assign _EVAL_436 = _EVAL_297 ? _EVAL_529 : _EVAL_193;
  assign _EVAL_821 = _EVAL_439 ? {{1'd0}, _EVAL_751} : _EVAL_599;
  assign _EVAL_701 = _EVAL_585 ? 1'h0 : 1'h1;
  assign _EVAL_274 = _EVAL_168 ? _EVAL_458 : _EVAL_596;
  assign _EVAL_881 = _EVAL_535 ? {{1'd0}, _EVAL_480} : _EVAL_355;
  assign _EVAL_714 = _EVAL_153 ? {{1'd0}, _EVAL_133} : _EVAL_443;
  assign _EVAL_617 = 2'h2 | _EVAL_474;
  assign _EVAL_423 = _EVAL_385 ? 1'h0 : 1'h1;
  assign _EVAL_879 = _EVAL_244 >= _EVAL_275;
  assign _EVAL_376 = _EVAL_280 ? 1'h0 : 1'h1;
  assign _EVAL_197 = _EVAL_282 ? 1'h0 : 1'h1;
  assign _EVAL_596 = {_EVAL_523,_EVAL_56};
  assign _EVAL_240 = _EVAL_436 >= _EVAL_265;
  assign _EVAL_326 = {_EVAL_776,_EVAL_96};
  assign _EVAL_180 = _EVAL_829 >= _EVAL_145;
  assign _EVAL_760 = _EVAL_318 ? {{1'd0}, _EVAL_134} : _EVAL_629;
  assign _EVAL_615 = {{1'd0}, _EVAL_369};
  assign _EVAL_192 = {_EVAL_131,_EVAL_119};
  assign _EVAL_418 = _EVAL_472 ? _EVAL_528 : _EVAL_779;
  assign _EVAL_599 = 2'h2 | _EVAL_229;
  assign _EVAL_150 = 3'h4 | _EVAL_577;
  assign _EVAL_563 = {_EVAL_656,_EVAL_108};
  assign _EVAL_847 = _EVAL_516 ? 1'h0 : 1'h1;
  assign _EVAL_775 = _EVAL_722 ? {{1'd0}, _EVAL_224} : _EVAL_262;
  assign _EVAL_86 = _EVAL_681 ? {{1'd0}, _EVAL_697} : _EVAL_353;
  assign _EVAL_275 = {_EVAL_181,_EVAL_50};
  assign _EVAL_839 = _EVAL_168 ? 1'h0 : 1'h1;
  assign _EVAL_384 = {_EVAL_511,_EVAL_104};
  assign _EVAL_497 = _EVAL_817 ? _EVAL_154 : _EVAL_344;
  assign _EVAL_161 = _EVAL_627 ? 1'h0 : 1'h1;
  assign _EVAL_687 = _EVAL_48[47];
  assign _EVAL_578 = {_EVAL_288,_EVAL_41};
  assign _EVAL_401 = _EVAL_240 ? _EVAL_436 : _EVAL_265;
  assign _EVAL_452 = _EVAL_489 ? _EVAL_177 : _EVAL_293;
  assign _EVAL_446 = _EVAL_402 ? {{1'd0}, _EVAL_761} : _EVAL_147;
  assign _EVAL_644 = _EVAL_883 ? 1'h0 : 1'h1;
  assign _EVAL_252 = {_EVAL_640,_EVAL_74};
  assign _EVAL_791 = _EVAL_306 >= _EVAL_869;
  assign _EVAL_413 = {_EVAL_340,_EVAL_20};
  assign _EVAL_733 = _EVAL_381 ? _EVAL_679 : _EVAL_647;
  assign _EVAL_285 = _EVAL_692 >= _EVAL_391;
  assign _EVAL_259 = _EVAL_732 ? _EVAL_825 : _EVAL_680;
  assign _EVAL_305 = 2'h2 | _EVAL_624;
  assign _EVAL_513 = _EVAL_728 >= _EVAL_802;
  assign _EVAL_257 = _EVAL_858 ? _EVAL_350 : _EVAL_356;
  assign _EVAL_678 = _EVAL_740 ? _EVAL_590 : _EVAL_707;
  assign _EVAL_137 = _EVAL_302 ? _EVAL_810 : _EVAL_639;
  assign _EVAL_247 = {_EVAL_792,_EVAL_81};
  assign _EVAL_822 = {_EVAL_875,_EVAL_45};
  assign _EVAL_345 = _EVAL_225 ? _EVAL_538 : _EVAL_292;
  assign _EVAL_255 = _EVAL_48[73];
  assign _EVAL_857 = _EVAL_48[92];
  assign _EVAL_266 = {_EVAL_515,_EVAL_25};
  assign _EVAL_363 = {_EVAL_438,_EVAL_61};
  assign _EVAL_699 = {_EVAL_400,_EVAL_2};
  assign _EVAL_391 = _EVAL_395 ? _EVAL_713 : _EVAL_406;
  assign _EVAL_151 = _EVAL_842 ? _EVAL_864 : _EVAL_135;
  assign _EVAL_483 = {_EVAL_658,_EVAL_110};
  assign _EVAL_437 = _EVAL_455 ? {{1'd0}, _EVAL_311} : _EVAL_828;
  assign _EVAL_225 = _EVAL_538 >= _EVAL_292;
  assign _EVAL_245 = 3'h4 | _EVAL_407;
  assign _EVAL_287 = _EVAL_733 >= _EVAL_392;
  assign _EVAL_199 = _EVAL_739 >= _EVAL_271;
  assign _EVAL_572 = {_EVAL_778,_EVAL_118};
  assign _EVAL_319 = _EVAL_550 ? {{1'd0}, _EVAL_886} : _EVAL_587;
  assign _EVAL_429 = _EVAL_239 >= _EVAL_482;
  assign _EVAL_336 = {_EVAL_256,_EVAL_24};
  assign _EVAL_301 = _EVAL_669 >= _EVAL_475;
  assign _EVAL_331 = 3'h4 | _EVAL_414;
  assign _EVAL_685 = {{1'd0}, _EVAL_226};
  assign _EVAL_264 = _EVAL_659 >= _EVAL_303;
  assign _EVAL_297 = _EVAL_529 >= _EVAL_193;
  assign _EVAL_555 = {_EVAL_498,_EVAL_57};
  assign _EVAL_531 = _EVAL_48[79];
  assign _EVAL_294 = {_EVAL_272,_EVAL_27};
  assign _EVAL_170 = _EVAL_689 ? _EVAL_807 : _EVAL_237;
  assign _EVAL_339 = _EVAL_48[98];
  assign _EVAL_522 = _EVAL_845 ? _EVAL_384 : _EVAL_711;
  assign _EVAL_210 = _EVAL_48[124];
  assign _EVAL_491 = _EVAL_879 ? 1'h0 : 1'h1;
  assign _EVAL_470 = _EVAL_48[59];
  assign _EVAL_526 = _EVAL_48[14];
  assign _EVAL_606 = {_EVAL_492,_EVAL_59};
  assign _EVAL_878 = _EVAL_543 >= _EVAL_435;
  assign _EVAL_601 = _EVAL_759 ? _EVAL_461 : _EVAL_768;
  assign _EVAL_130 = _EVAL_572 >= _EVAL_326;
  assign _EVAL_322 = _EVAL_798 ? {{1'd0}, _EVAL_773} : _EVAL_360;
  assign _EVAL_390 = _EVAL_48[95];
  assign _EVAL_782 = _EVAL_756 ? 1'h0 : 1'h1;
  assign _EVAL_251 = _EVAL_702 ? _EVAL_712 : _EVAL_870;
  assign _EVAL_498 = _EVAL_48[49];
  assign _EVAL_160 = {{1'd0}, _EVAL_432};
  assign _EVAL_156 = {_EVAL_339,_EVAL_62};
  assign _EVAL_667 = {{1'd0}, _EVAL_520};
  assign _EVAL_141 = 2'h2 | _EVAL_641;
  assign _EVAL_681 = _EVAL_401 >= _EVAL_497;
  assign _EVAL_590 = _EVAL_261 ? _EVAL_506 : _EVAL_512;
  assign _EVAL_459 = _EVAL_48[62];
  assign _EVAL_469 = _EVAL_203 ? 1'h0 : 1'h1;
  assign _EVAL_267 = _EVAL_48[112];
  assign _EVAL_328 = _EVAL_873 >= _EVAL_380;
  assign _EVAL_490 = _EVAL_570 ? 1'h0 : 1'h1;
  assign _EVAL_885 = _EVAL_214 ? _EVAL_567 : _EVAL_234;
  assign _EVAL_804 = _EVAL_872 >= _EVAL_257;
  assign _EVAL_652 = {_EVAL_410,_EVAL_4};
  assign _EVAL_817 = _EVAL_154 >= _EVAL_344;
  assign _EVAL_365 = _EVAL_48[44];
  assign _EVAL_840 = {{1'd0}, _EVAL_233};
  assign _EVAL_424 = {{1'd0}, _EVAL_533};
  assign _EVAL_693 = _EVAL_48[71];
  assign _EVAL_183 = _EVAL_281 >= _EVAL_835;
  assign _EVAL_158 = _EVAL_689 ? {{1'd0}, _EVAL_731} : _EVAL_317;
  assign _EVAL_867 = _EVAL_824 ? 1'h0 : 1'h1;
  assign _EVAL_484 = _EVAL_830 ? {{1'd0}, _EVAL_665} : _EVAL_208;
  assign _EVAL_450 = _EVAL_795 ? _EVAL_151 : _EVAL_166;
  assign _EVAL_230 = {_EVAL_470,_EVAL_97};
  assign _EVAL_260 = 3'h4 | _EVAL_241;
  assign _EVAL_772 = {_EVAL_626,_EVAL_73};
  assign _EVAL_783 = _EVAL_48[9];
  assign _EVAL_551 = {{1'd0}, _EVAL_852};
  assign _EVAL_178 = {{1'd0}, _EVAL_491};
  assign _EVAL_547 = _EVAL_48[10];
  assign _EVAL_855 = {_EVAL_693,_EVAL_121};
  assign _EVAL_683 = _EVAL_754 >= _EVAL_473;
  assign _EVAL_371 = {{1'd0}, _EVAL_184};
  assign _EVAL_330 = _EVAL_558 ? _EVAL_162 : _EVAL_525;
  assign _EVAL_575 = _EVAL_48[53];
  assign _EVAL_449 = _EVAL_404 ? 1'h0 : 1'h1;
  assign _EVAL_621 = _EVAL_48[123];
  assign _EVAL_716 = _EVAL_48[80];
  assign _EVAL_494 = {_EVAL_694,_EVAL_6};
  assign _EVAL_836 = _EVAL_308 ? 1'h0 : 1'h1;
  assign _EVAL_739 = _EVAL_402 ? _EVAL_884 : _EVAL_186;
  assign _EVAL_321 = 2'h2 | _EVAL_191;
  assign _EVAL_536 = _EVAL_343 ? _EVAL_476 : _EVAL_885;
  assign _EVAL_629 = 4'h8 | _EVAL_632;
  assign _EVAL_624 = {{1'd0}, _EVAL_736};
  assign _EVAL_568 = _EVAL_48[30];
  assign _EVAL_728 = {_EVAL_600,_EVAL_88};
  assign _EVAL_327 = _EVAL_709 >= _EVAL_838;
  assign _EVAL_414 = {{1'd0}, _EVAL_881};
  assign _EVAL_558 = _EVAL_162 >= _EVAL_525;
  assign _EVAL_462 = _EVAL_266 >= _EVAL_633;
  assign _EVAL_740 = _EVAL_590 >= _EVAL_707;
  assign _EVAL_179 = 2'h2 | _EVAL_745;
  assign _EVAL_706 = 3'h4 | _EVAL_499;
  assign _EVAL_833 = _EVAL_564 ? 1'h0 : 1'h1;
  assign _EVAL_859 = _EVAL_263 >= _EVAL_213;
  assign _EVAL_815 = _EVAL_634 ? _EVAL_583 : _EVAL_440;
  assign _EVAL_516 = _EVAL_861 >= _EVAL_721;
  assign _EVAL_713 = {_EVAL_614,_EVAL_94};
  assign _EVAL_309 = _EVAL_786 >= _EVAL_185;
  assign _EVAL_719 = _EVAL_766 >= _EVAL_704;
  assign _EVAL_343 = _EVAL_476 >= _EVAL_885;
  assign _EVAL_221 = _EVAL_48[16];
  assign _EVAL_175 = _EVAL_732 ? {{1'd0}, _EVAL_444} : _EVAL_880;
  assign _EVAL_539 = _EVAL_48[7];
  assign _EVAL_223 = _EVAL_48[50];
  assign _EVAL_672 = {_EVAL_622,_EVAL_10};
  assign _EVAL_761 = _EVAL_860 ? {{1'd0}, _EVAL_376} : _EVAL_486;
  assign _EVAL_594 = {{1'd0}, _EVAL_698};
  assign _EVAL_378 = _EVAL_48[4];
  assign _EVAL_777 = 2'h2 | _EVAL_718;
  assign _EVAL_428 = _EVAL_48[84];
  assign _EVAL_626 = _EVAL_48[99];
  assign _EVAL_269 = {_EVAL_831,_EVAL_117};
  assign _EVAL_65 = _EVAL_648[2:0];
  assign _EVAL_357 = _EVAL_48[31];
  assign _EVAL_487 = {_EVAL_366,_EVAL_112};
  assign _EVAL_519 = _EVAL_48[36];
  assign _EVAL_273 = _EVAL_48[32];
  assign _EVAL_825 = _EVAL_510 ? _EVAL_269 : _EVAL_451;
  assign _EVAL_249 = _EVAL_48[97];
  assign _EVAL_864 = _EVAL_756 ? _EVAL_589 : _EVAL_192;
  assign _EVAL_189 = _EVAL_719 ? _EVAL_766 : _EVAL_704;
  assign _EVAL_767 = _EVAL_264 ? {{1'd0}, _EVAL_490} : _EVAL_549;
  assign _EVAL_875 = _EVAL_48[6];
  assign _EVAL_456 = _EVAL_795 ? {{1'd0}, _EVAL_397} : _EVAL_774;
  assign _EVAL_868 = _EVAL_258 ? _EVAL_598 : _EVAL_373;
  assign _EVAL_837 = {_EVAL_298,_EVAL_30};
  assign _EVAL_244 = {_EVAL_434,_EVAL_76};
  assign _EVAL_492 = _EVAL_48[28];
  assign _EVAL_387 = 4'h8 | _EVAL_540;
  assign _EVAL_579 = _EVAL_394 >= _EVAL_342;
  assign _EVAL_690 = {{1'd0}, _EVAL_720};
  assign _EVAL_250 = _EVAL_536 >= _EVAL_450;
  assign _EVAL_712 = _EVAL_507 ? _EVAL_422 : _EVAL_846;
  assign _EVAL_803 = _EVAL_48[22];
  assign _EVAL_741 = _EVAL_845 ? 1'h0 : 1'h1;
  assign _EVAL_404 = _EVAL_738 >= _EVAL_187;
  assign _EVAL_806 = _EVAL_742 ? _EVAL_230 : _EVAL_232;
  assign _EVAL_368 = 2'h2 | _EVAL_729;
  assign _EVAL_651 = _EVAL_504 ? 1'h0 : 1'h1;
  assign _EVAL_448 = _EVAL_48[24];
  assign _EVAL_209 = _EVAL_672 >= _EVAL_850;
  assign _EVAL_861 = {_EVAL_405,_EVAL_103};
  assign _EVAL_524 = _EVAL_48[34];
  assign _EVAL_461 = {_EVAL_799,_EVAL_99};
  assign _EVAL_661 = {{1'd0}, _EVAL_812};
  assign _EVAL_457 = {{1'd0}, _EVAL_325};
  assign _EVAL_515 = _EVAL_48[3];
  assign _EVAL_694 = _EVAL_48[66];
  assign _EVAL_464 = {_EVAL_604,_EVAL_37};
  assign _EVAL_888 = {{1'd0}, _EVAL_849};
  assign _EVAL_308 = _EVAL_699 >= _EVAL_494;
  assign _EVAL_882 = _EVAL_330 >= _EVAL_248;
  assign _EVAL_858 = _EVAL_350 >= _EVAL_356;
  assign _EVAL_471 = _EVAL_130 ? 1'h0 : 1'h1;
  assign _EVAL_426 = {{1'd0}, _EVAL_836};
  assign _EVAL_759 = _EVAL_461 >= _EVAL_768;
  assign _EVAL_807 = _EVAL_453 ? _EVAL_251 : _EVAL_508;
  assign _EVAL_587 = 3'h4 | _EVAL_727;
  assign _EVAL_797 = _EVAL_637 ? _EVAL_416 : _EVAL_278;
  assign _EVAL_720 = _EVAL_858 ? {{1'd0}, _EVAL_823} : _EVAL_848;
  assign _EVAL_465 = _EVAL_206 >= _EVAL_383;
  assign _EVAL_310 = _EVAL_817 ? {{1'd0}, _EVAL_670} : _EVAL_417;
  assign _EVAL_201 = _EVAL_359 ? 1'h0 : 1'h1;
  assign _EVAL_142 = _EVAL_715 ? {{1'd0}, _EVAL_484} : _EVAL_663;
  assign _EVAL_614 = _EVAL_48[89];
  assign _EVAL_453 = _EVAL_251 >= _EVAL_508;
  assign _EVAL_565 = _EVAL_560 >= _EVAL_606;
  assign _EVAL_364 = _EVAL_242 >= _EVAL_346;
  assign _EVAL_148 = _EVAL_48[35];
  assign _EVAL_871 = _EVAL_48[82];
  assign _EVAL_393 = _EVAL_48[81];
  assign _EVAL_352 = 3'h4 | _EVAL_671;
  assign _EVAL_355 = 2'h2 | _EVAL_888;
  assign _EVAL_341 = {{1'd0}, _EVAL_644};
  assign _EVAL_412 = {{1'd0}, _EVAL_605};
  assign _EVAL_466 = _EVAL_48[29];
  assign _EVAL_212 = _EVAL_207 ? _EVAL_247 : _EVAL_595;
  assign _EVAL_605 = _EVAL_865 ? {{1'd0}, _EVAL_290} : _EVAL_331;
  assign _EVAL_302 = _EVAL_810 >= _EVAL_639;
  assign _EVAL_254 = _EVAL_381 ? 1'h0 : 1'h1;
  assign _EVAL_620 = _EVAL_246 ? _EVAL_329 : _EVAL_212;
  assign _EVAL_743 = _EVAL_878 ? _EVAL_543 : _EVAL_435;
  assign _EVAL_780 = {_EVAL_255,_EVAL_87};
  assign _EVAL_508 = _EVAL_264 ? _EVAL_659 : _EVAL_303;
  assign _EVAL_789 = 2'h2 | _EVAL_661;
  assign _EVAL_532 = _EVAL_132 ? _EVAL_652 : _EVAL_563;
  assign _EVAL_318 = _EVAL_314 >= _EVAL_796;
  assign _EVAL_382 = _EVAL_588 ? {{1'd0}, _EVAL_319} : _EVAL_220;
  assign _EVAL_808 = _EVAL_170 >= _EVAL_546;
  assign _EVAL_850 = {_EVAL_705,_EVAL_84};
  assign _EVAL_389 = _EVAL_562 >= _EVAL_294;
  assign _EVAL_400 = _EVAL_48[65];
  assign _EVAL_334 = _EVAL_517 ? 1'h0 : 1'h1;
  assign _EVAL_280 = _EVAL_276 >= _EVAL_190;
  assign _EVAL_692 = _EVAL_787 ? _EVAL_578 : _EVAL_313;
  assign _EVAL_415 = {_EVAL_548,_EVAL_36};
  assign _EVAL_527 = {_EVAL_138,_EVAL};
  assign _EVAL_643 = _EVAL_48[119];
  assign _EVAL_675 = 4'h8 | _EVAL_371;
  assign _EVAL_589 = {_EVAL_696,_EVAL_85};
  assign _EVAL_598 = {_EVAL_217,_EVAL_68};
  assign _EVAL_581 = {{1'd0}, _EVAL_310};
  assign _EVAL_549 = 2'h2 | _EVAL_615;
  assign _EVAL_472 = _EVAL_528 >= _EVAL_779;
  assign _EVAL_873 = {_EVAL_863,_EVAL_91};
  assign _EVAL_419 = _EVAL_258 ? 1'h0 : 1'h1;
  assign _EVAL_689 = _EVAL_807 >= _EVAL_237;
  assign _EVAL_637 = _EVAL_416 >= _EVAL_278;
  assign _EVAL_182 = 3'h4 | _EVAL_569;
  assign _EVAL_860 = _EVAL_299 >= _EVAL_717;
  assign _EVAL_765 = 3'h4 | _EVAL_222;
  assign _EVAL_812 = _EVAL_207 ? 1'h0 : 1'h1;
  assign _EVAL_653 = _EVAL_48[102];
  assign _EVAL_851 = _EVAL_48[63];
  assign _EVAL_258 = _EVAL_598 >= _EVAL_373;
  assign _EVAL_346 = {_EVAL_377,_EVAL_52};
  assign _EVAL_146 = 5'h10 | _EVAL_295;
  assign _EVAL_495 = _EVAL_788 ? _EVAL_592 : _EVAL_762;
  assign _EVAL_474 = {{1'd0}, _EVAL_556};
  assign _EVAL_523 = _EVAL_48[8];
  assign _EVAL_445 = _EVAL_132 ? 1'h0 : 1'h1;
  assign _EVAL_154 = _EVAL_841 ? _EVAL_611 : _EVAL_678;
  assign _EVAL_669 = {_EVAL_493,_EVAL_12};
  assign _EVAL_496 = _EVAL_495 >= _EVAL_532;
  assign _EVAL_133 = _EVAL_559 ? {{1'd0}, _EVAL_195} : _EVAL_876;
  assign _EVAL_583 = {_EVAL_467,_EVAL_125};
  assign _EVAL_288 = _EVAL_48[87];
  assign _EVAL_744 = {{1'd0}, _EVAL_821};
  assign _EVAL_676 = {{1'd0}, _EVAL_423};
  assign _EVAL_845 = _EVAL_384 >= _EVAL_711;
  assign _EVAL_542 = _EVAL_180 ? _EVAL_829 : _EVAL_145;
  assign _EVAL_340 = _EVAL_48[57];
  assign _EVAL_366 = _EVAL_48[46];
  assign _EVAL_290 = _EVAL_180 ? {{1'd0}, _EVAL_701} : _EVAL_617;
  assign _EVAL_228 = _EVAL_48[114];
  assign _EVAL_350 = _EVAL_642 ? _EVAL_485 : _EVAL_631;
  assign _EVAL_314 = _EVAL_882 ? _EVAL_330 : _EVAL_248;
  assign _EVAL_727 = {{1'd0}, _EVAL_454};
  assign _EVAL_353 = 7'h40 | _EVAL_581;
  assign _EVAL_482 = {_EVAL_243,_EVAL_69};
  assign _EVAL_283 = _EVAL_788 ? 1'h0 : 1'h1;
  assign _EVAL_538 = _EVAL_565 ? _EVAL_560 : _EVAL_606;
  assign _EVAL_143 = _EVAL_48[126];
  assign _EVAL_489 = _EVAL_177 >= _EVAL_293;
  assign _EVAL_196 = {{1'd0}, _EVAL_651};
  assign _EVAL_778 = _EVAL_48[17];
  assign _EVAL_548 = _EVAL_48[117];
  assign _EVAL_805 = {{1'd0}, _EVAL_586};
  assign _EVAL_243 = _EVAL_48[68];
  assign _EVAL_300 = _EVAL_274 >= _EVAL_189;
  assign _EVAL_380 = {_EVAL_662,_EVAL_44};
  assign _EVAL_349 = 2'h2 | _EVAL_424;
  assign _EVAL_172 = {_EVAL_755,_EVAL_60};
  assign _EVAL_793 = _EVAL_683 ? {{1'd0}, _EVAL_714} : _EVAL_501;
  assign _EVAL_546 = _EVAL_683 ? _EVAL_754 : _EVAL_473;
  assign _EVAL_377 = _EVAL_48[120];
  assign _EVAL_811 = 2'h2 | _EVAL_649;
  assign _EVAL_790 = _EVAL_48[12];
  assign _EVAL_738 = {_EVAL_393,_EVAL_126};
  assign _EVAL_788 = _EVAL_592 >= _EVAL_762;
  assign _EVAL_633 = {_EVAL_378,_EVAL_5};
  assign _EVAL_584 = {_EVAL_653,_EVAL_42};
  assign _EVAL_838 = {_EVAL_210,_EVAL_55};
  assign _EVAL_619 = 4'h8 | _EVAL_684;
  assign _EVAL_306 = {_EVAL_763,_EVAL_102};
  assign _EVAL_409 = _EVAL_887 ? _EVAL_806 : _EVAL_509;
  assign _EVAL_703 = {{1'd0}, _EVAL_874};
  assign _EVAL_507 = _EVAL_422 >= _EVAL_846;
  assign _EVAL_798 = _EVAL_813 >= _EVAL_868;
  assign _EVAL_226 = _EVAL_740 ? {{1'd0}, _EVAL_163} : _EVAL_387;
  assign _EVAL_688 = _EVAL_855 >= _EVAL_566;
  assign _EVAL_569 = {{1'd0}, _EVAL_479};
  assign _EVAL_348 = {_EVAL_249,_EVAL_63};
  assign _EVAL_485 = _EVAL_287 ? _EVAL_733 : _EVAL_392;
  assign _EVAL_502 = _EVAL_297 ? {{1'd0}, _EVAL_760} : _EVAL_146;
  assign _EVAL_809 = 2'h2 | _EVAL_312;
  assign _EVAL_132 = _EVAL_652 >= _EVAL_563;
  assign _EVAL_208 = 2'h2 | _EVAL_667;
  assign _EVAL_646 = {_EVAL_374,_EVAL_127};
  assign _EVAL_730 = {{1'd0}, _EVAL_793};
  assign _EVAL_479 = _EVAL_214 ? {{1'd0}, _EVAL_235} : _EVAL_321;
  assign _EVAL_543 = {_EVAL_129,_EVAL_66};
  assign _EVAL_749 = 6'h20 | _EVAL_805;
  assign _EVAL_567 = _EVAL_173 ? _EVAL_333 : _EVAL_420;
  assign _EVAL_648 = _EVAL_681 ? _EVAL_401 : _EVAL_497;
  assign _EVAL_521 = _EVAL_747 ? {{1'd0}, _EVAL_388} : _EVAL_349;
  assign _EVAL_514 = _EVAL_403 >= _EVAL_259;
  assign _EVAL_440 = {_EVAL_758,_EVAL_120};
  assign _EVAL_427 = _EVAL_834 ? 1'h0 : 1'h1;
  assign _EVAL_520 = _EVAL_301 ? 1'h0 : 1'h1;
  assign _EVAL_751 = _EVAL_327 ? 1'h0 : 1'h1;
  assign _EVAL_670 = _EVAL_841 ? {{1'd0}, _EVAL_347} : _EVAL_826;
  assign _EVAL_582 = _EVAL_579 ? _EVAL_394 : _EVAL_342;
  assign _EVAL_796 = _EVAL_514 ? _EVAL_403 : _EVAL_259;
  assign _EVAL_216 = {_EVAL_223,_EVAL_80};
  assign _EVAL_779 = {_EVAL_623,_EVAL_22};
  assign _EVAL_500 = _EVAL_404 ? _EVAL_738 : _EVAL_187;
  assign _EVAL_604 = _EVAL_48[33];
  assign _EVAL_666 = _EVAL_522 >= _EVAL_505;
  assign _EVAL_441 = {_EVAL_463,_EVAL_33};
  assign _EVAL_877 = _EVAL_753 ? 1'h0 : 1'h1;
  assign _EVAL_203 = _EVAL_370 >= _EVAL_757;
  assign _EVAL_278 = {_EVAL_267,_EVAL_105};
  assign _EVAL_603 = _EVAL_48[19];
  assign _EVAL_574 = _EVAL_48[109];
  assign _EVAL_556 = _EVAL_610 ? 1'h0 : 1'h1;
  assign _EVAL_324 = _EVAL_48[105];
  assign _EVAL_139 = _EVAL_246 ? {{1'd0}, _EVAL_442} : _EVAL_789;
  assign _EVAL_475 = {_EVAL_816,_EVAL_72};
  assign _EVAL_135 = _EVAL_627 ? _EVAL_635 : _EVAL_660;
  assign _EVAL_732 = _EVAL_825 >= _EVAL_680;
  assign _EVAL_311 = _EVAL_634 ? 1'h0 : 1'h1;
  assign _EVAL_866 = 2'h2 | _EVAL_196;
  assign _EVAL_611 = _EVAL_199 ? _EVAL_739 : _EVAL_271;
  assign _EVAL_291 = _EVAL_358 ? _EVAL_320 : _EVAL_646;
  assign _EVAL_164 = {_EVAL_568,_EVAL_70};
  assign _EVAL_395 = _EVAL_713 >= _EVAL_406;
  assign _EVAL_715 = _EVAL_433 >= _EVAL_345;
  assign _EVAL_420 = {_EVAL_519,_EVAL_122};
  assign _EVAL_560 = {_EVAL_534,_EVAL_128};
  assign _EVAL_691 = _EVAL_452 >= _EVAL_573;
  assign _EVAL_673 = _EVAL_550 ? _EVAL_544 : _EVAL_431;
  assign _EVAL_810 = _EVAL_389 ? _EVAL_562 : _EVAL_294;
  assign _EVAL_332 = {_EVAL_636,_EVAL_89};
  assign _EVAL_554 = _EVAL_285 ? {{1'd0}, _EVAL_218} : _EVAL_856;
  assign _EVAL_458 = {_EVAL_539,_EVAL_19};
  assign _EVAL_402 = _EVAL_884 >= _EVAL_186;
  assign _EVAL_504 = _EVAL_654 >= _EVAL_487;
  assign _EVAL_722 = _EVAL_176 >= _EVAL_630;
  assign _EVAL_766 = {_EVAL_783,_EVAL_29};
  assign _EVAL_668 = _EVAL_48[111];
  assign _EVAL_312 = {{1'd0}, _EVAL_833};
  assign _EVAL_435 = {_EVAL_803,_EVAL_14};
  assign _EVAL_729 = {{1'd0}, _EVAL_375};
  assign _EVAL_351 = _EVAL_48[0];
  assign _EVAL_200 = _EVAL_462 ? _EVAL_266 : _EVAL_633;
  assign _EVAL_282 = _EVAL_464 >= _EVAL_593;
  assign _EVAL_576 = _EVAL_282 ? _EVAL_464 : _EVAL_593;
  assign _EVAL_155 = _EVAL_225 ? {{1'd0}, _EVAL_746} : _EVAL_305;
  assign _EVAL_289 = {{1'd0}, _EVAL_775};
  assign _EVAL_649 = {{1'd0}, _EVAL_197};
  assign _EVAL_397 = _EVAL_842 ? {{1'd0}, _EVAL_782} : _EVAL_801;
  assign _EVAL_233 = _EVAL_808 ? {{1'd0}, _EVAL_158} : _EVAL_608;
  assign _EVAL_595 = {_EVAL_545,_EVAL_7};
  assign _EVAL_385 = _EVAL_336 >= _EVAL_421;
  assign _EVAL_533 = _EVAL_140 ? 1'h0 : 1'h1;
  assign _EVAL_165 = _EVAL_48[104];
  assign _EVAL_663 = 3'h4 | _EVAL_814;
  assign _EVAL_634 = _EVAL_583 >= _EVAL_440;
  assign _EVAL_256 = _EVAL_48[113];
  assign _EVAL_844 = {{1'd0}, _EVAL_521};
  assign _EVAL_299 = _EVAL_280 ? _EVAL_276 : _EVAL_190;
  assign _EVAL_173 = _EVAL_333 >= _EVAL_420;
  assign _EVAL_707 = _EVAL_723 ? _EVAL_530 : _EVAL_620;
  assign _EVAL_639 = _EVAL_883 ? _EVAL_413 : _EVAL_527;
  assign _EVAL_166 = _EVAL_231 ? _EVAL_557 : _EVAL_236;
  assign _EVAL_236 = _EVAL_504 ? _EVAL_654 : _EVAL_487;
  assign _EVAL_682 = _EVAL_202 ? 1'h0 : 1'h1;
  assign _EVAL_846 = {_EVAL_396,_EVAL_17};
  assign _EVAL_573 = _EVAL_496 ? _EVAL_495 : _EVAL_532;
  assign _EVAL_444 = _EVAL_510 ? 1'h0 : 1'h1;
  assign _EVAL_525 = _EVAL_879 ? _EVAL_244 : _EVAL_275;
  assign _EVAL_762 = {_EVAL_284,_EVAL_32};
  assign _EVAL_167 = {{1'd0}, _EVAL_334};
  assign _EVAL_654 = {_EVAL_270,_EVAL_107};
  assign _EVAL_829 = _EVAL_585 ? _EVAL_337 : _EVAL_316;
  assign _EVAL_802 = {_EVAL_857,_EVAL_109};
  assign _EVAL_281 = {_EVAL_204,_EVAL_46};
  assign _EVAL_510 = _EVAL_269 >= _EVAL_451;
  assign _EVAL_530 = _EVAL_285 ? _EVAL_692 : _EVAL_391;
  assign _EVAL_144 = _EVAL_781 ? _EVAL_399 : _EVAL_794;
  assign _EVAL_814 = {{1'd0}, _EVAL_155};
  assign _EVAL_843 = _EVAL_514 ? {{1'd0}, _EVAL_468} : _EVAL_245;
  assign _EVAL_638 = _EVAL_759 ? 1'h0 : 1'h1;
  assign _EVAL_320 = {_EVAL_603,_EVAL_111};
  assign _EVAL_272 = _EVAL_48[56];
  assign _EVAL_284 = _EVAL_48[76];
  assign _EVAL_747 = _EVAL_200 >= _EVAL_674;
  assign _EVAL_816 = _EVAL_48[26];
  assign _EVAL_335 = _EVAL_48[90];
  assign _EVAL_786 = {_EVAL_227,_EVAL_38};
  assign _EVAL_842 = _EVAL_864 >= _EVAL_135;
  assign _EVAL_776 = _EVAL_48[18];
  assign _EVAL_588 = _EVAL_673 >= _EVAL_561;
  assign _EVAL_394 = {_EVAL_574,_EVAL_64};
  assign _EVAL_518 = _EVAL_48[86];
  assign _EVAL_607 = _EVAL_358 ? 1'h0 : 1'h1;
  assign _EVAL_323 = _EVAL_702 ? {{1'd0}, _EVAL_136} : _EVAL_179;
  assign _EVAL_195 = _EVAL_637 ? 1'h0 : 1'h1;
  assign _EVAL_792 = _EVAL_48[93];
  assign _EVAL_403 = _EVAL_300 ? _EVAL_274 : _EVAL_189;
  assign _EVAL_373 = {_EVAL_518,_EVAL_43};
  assign _EVAL_253 = _EVAL_395 ? 1'h0 : 1'h1;
  assign _EVAL_405 = _EVAL_48[43];
  assign _EVAL_734 = 2'h2 | _EVAL_178;
  assign _EVAL_506 = _EVAL_800 ? _EVAL_597 : _EVAL_500;
  assign _EVAL_710 = {{1'd0}, _EVAL_867};
  assign _EVAL_848 = 4'h8 | _EVAL_703;
  assign _EVAL_317 = 4'h8 | _EVAL_412;
  assign _EVAL_213 = _EVAL_564 ? _EVAL_770 : _EVAL_268;
  assign _EVAL_202 = 4'h8 >= _EVAL_724;
  assign _EVAL_647 = {_EVAL_238,_EVAL_98};
  assign _EVAL_190 = {_EVAL_481,_EVAL_31};
  assign _EVAL_279 = _EVAL_48[110];
  assign _EVAL_545 = _EVAL_48[94];
  assign _EVAL_356 = _EVAL_286 ? _EVAL_137 : _EVAL_409;
  assign _EVAL_425 = {_EVAL_575,_EVAL_11};
  assign _EVAL_430 = _EVAL_429 ? 1'h0 : 1'h1;
  assign _EVAL_769 = {{1'd0}, _EVAL_253};
  assign _EVAL_313 = {_EVAL_361,_EVAL_71};
  assign _EVAL_541 = _EVAL_48[60];
  assign _EVAL_535 = _EVAL_418 >= _EVAL_582;
  assign _EVAL_696 = _EVAL_48[39];
  assign _EVAL_432 = _EVAL_686 ? 1'h0 : 1'h1;
  assign _EVAL_725 = _EVAL_328 ? 1'h0 : 1'h1;
  assign _EVAL_820 = 2'h2 | _EVAL_411;
  assign _EVAL_248 = _EVAL_747 ? _EVAL_200 : _EVAL_674;
  assign _EVAL_659 = _EVAL_570 ? _EVAL_772 : _EVAL_700;
  assign _EVAL_695 = 3'h4 | _EVAL_844;
  assign _EVAL_198 = 2'h2 | _EVAL_362;
  assign _EVAL_211 = _EVAL_887 ? {{1'd0}, _EVAL_708} : _EVAL_735;
  assign _EVAL_597 = _EVAL_465 ? _EVAL_206 : _EVAL_383;
  assign _EVAL_544 = _EVAL_666 ? _EVAL_522 : _EVAL_505;
  assign _EVAL_764 = _EVAL_48[75];
  assign _EVAL_358 = _EVAL_320 >= _EVAL_646;
  assign _EVAL_571 = _EVAL_302 ? {{1'd0}, _EVAL_737} : _EVAL_537;
  assign _EVAL_467 = _EVAL_48[51];
  assign _EVAL_388 = _EVAL_462 ? 1'h0 : 1'h1;
  assign _EVAL_593 = {_EVAL_524,_EVAL_95};
  assign _EVAL_386 = {_EVAL_466,_EVAL_49};
  assign _EVAL_552 = {_EVAL_324,_EVAL_100};
  assign _EVAL_442 = _EVAL_513 ? 1'h0 : 1'h1;
  assign _EVAL_503 = _EVAL_332 >= _EVAL_584;
  assign _EVAL_486 = 2'h2 | _EVAL_426;
  assign _EVAL_185 = {_EVAL_526,_EVAL_18};
  assign _EVAL_176 = _EVAL_859 ? _EVAL_263 : _EVAL_213;
  assign _EVAL_374 = _EVAL_48[20];
  assign _EVAL_612 = {{1'd0}, _EVAL_142};
  assign _EVAL_162 = _EVAL_202 ? 4'h8 : _EVAL_724;
  assign _EVAL_705 = _EVAL_48[70];
  assign _EVAL_517 = _EVAL_425 >= _EVAL_837;
  assign _EVAL_869 = {_EVAL_428,_EVAL_106};
  assign _EVAL_580 = _EVAL_800 ? {{1'd0}, _EVAL_460} : _EVAL_820;
  assign _EVAL_329 = _EVAL_513 ? _EVAL_728 : _EVAL_802;
  assign _EVAL_745 = {{1'd0}, _EVAL_427};
  assign _EVAL_187 = {_EVAL_871,_EVAL_124};
  assign _EVAL_169 = _EVAL_48[121];
  assign _EVAL_184 = _EVAL_691 ? {{1'd0}, _EVAL_488} : _EVAL_352;
  assign _EVAL_129 = _EVAL_48[21];
  assign _EVAL_627 = _EVAL_635 >= _EVAL_660;
  assign _EVAL_338 = _EVAL_723 ? {{1'd0}, _EVAL_554} : _EVAL_706;
  assign _EVAL_292 = _EVAL_367 ? _EVAL_386 : _EVAL_164;
  assign _EVAL_631 = _EVAL_455 ? _EVAL_815 : _EVAL_379;
  assign _EVAL_407 = {{1'd0}, _EVAL_175};
  assign _EVAL_476 = _EVAL_650 ? _EVAL_771 : _EVAL_576;
  assign _EVAL_229 = {{1'd0}, _EVAL_638};
  assign _EVAL_447 = _EVAL_48[107];
  assign _EVAL_529 = _EVAL_318 ? _EVAL_314 : _EVAL_796;
  assign _EVAL_658 = _EVAL_48[37];
  assign _EVAL_824 = _EVAL_555 >= _EVAL_216;
  assign _EVAL_307 = _EVAL_688 ? 1'h0 : 1'h1;
  assign _EVAL_214 = _EVAL_567 >= _EVAL_234;
  assign _EVAL_293 = _EVAL_686 ? _EVAL_780 : _EVAL_616;
  assign _EVAL_433 = _EVAL_830 ? _EVAL_750 : _EVAL_827;
  assign _EVAL_697 = _EVAL_240 ? {{1'd0}, _EVAL_502} : _EVAL_749;
  assign _EVAL_205 = _EVAL_48[5];
  assign _EVAL_392 = _EVAL_824 ? _EVAL_555 : _EVAL_216;
  assign _EVAL_417 = 6'h20 | _EVAL_840;
  assign _EVAL_553 = _EVAL_385 ? _EVAL_336 : _EVAL_421;
  assign _EVAL_752 = 2'h2 | _EVAL_710;
  assign _EVAL_737 = _EVAL_389 ? 1'h0 : 1'h1;
  assign _EVAL_818 = _EVAL_48[67];
  assign _EVAL_369 = _EVAL_503 ? 1'h0 : 1'h1;
  assign _EVAL_488 = _EVAL_489 ? {{1'd0}, _EVAL_307} : _EVAL_832;
  assign _EVAL_136 = _EVAL_507 ? 1'h0 : 1'h1;
  assign _EVAL_337 = {_EVAL_748,_EVAL_53};
  assign _EVAL_528 = {_EVAL_447,_EVAL_0};
  assign _EVAL_664 = _EVAL_291 >= _EVAL_743;
  assign _EVAL_566 = {_EVAL_408,_EVAL_23};
  assign _EVAL_660 = {_EVAL_157,_EVAL_67};
  assign _EVAL_755 = _EVAL_48[118];
  assign _EVAL_830 = _EVAL_750 >= _EVAL_827;
  assign _EVAL_835 = {_EVAL_448,_EVAL_35};
  assign _EVAL_763 = _EVAL_48[83];
  assign _EVAL_152 = _EVAL_250 ? {{1'd0}, _EVAL_853} : _EVAL_619;
  assign _EVAL_561 = _EVAL_715 ? _EVAL_433 : _EVAL_345;
  assign _EVAL_398 = {{1'd0}, _EVAL_877};
  assign _EVAL_854 = _EVAL_558 ? {{1'd0}, _EVAL_682} : _EVAL_734;
  assign _EVAL_468 = _EVAL_300 ? {{1'd0}, _EVAL_839} : _EVAL_368;
  assign _EVAL_238 = _EVAL_48[48];
  assign _EVAL_640 = _EVAL_48[106];
  assign _EVAL_271 = _EVAL_691 ? _EVAL_452 : _EVAL_573;
  assign _EVAL_186 = _EVAL_478 ? _EVAL_219 : _EVAL_613;
  assign _EVAL_140 = _EVAL_296 >= _EVAL_822;
  assign _EVAL_451 = {_EVAL_790,_EVAL_93};
  assign _EVAL_880 = 2'h2 | _EVAL_477;
  assign _EVAL_586 = _EVAL_804 ? {{1'd0}, _EVAL_152} : _EVAL_602;
  assign _EVAL_632 = {{1'd0}, _EVAL_843};
  assign _EVAL_674 = _EVAL_140 ? _EVAL_296 : _EVAL_822;
  assign _EVAL_636 = _EVAL_48[101];
  assign _EVAL_876 = 2'h2 | _EVAL_676;
  assign _EVAL_224 = _EVAL_859 ? {{1'd0}, _EVAL_372} : _EVAL_809;
  assign _EVAL_623 = _EVAL_48[108];
  assign _EVAL_564 = _EVAL_770 >= _EVAL_268;
  assign _EVAL_537 = 2'h2 | _EVAL_341;
  assign _EVAL_381 = _EVAL_679 >= _EVAL_647;
  assign _EVAL_616 = {_EVAL_618,_EVAL_15};
  assign _EVAL_438 = _EVAL_48[61];
  assign _EVAL_753 = _EVAL_363 >= _EVAL_174;
  assign _EVAL_316 = {_EVAL_165,_EVAL_3};
  assign _EVAL_557 = _EVAL_516 ? _EVAL_861 : _EVAL_721;
  assign _EVAL_481 = _EVAL_48[64];
  assign _EVAL_235 = _EVAL_173 ? 1'h0 : 1'h1;
  assign _EVAL_159 = _EVAL_496 ? {{1'd0}, _EVAL_283} : _EVAL_141;
  assign _EVAL_758 = _EVAL_48[52];
  assign _EVAL_726 = _EVAL_48[41];
  assign _EVAL_270 = _EVAL_48[45];
  assign _EVAL_577 = {{1'd0}, _EVAL_322};
  assign _EVAL_785 = {{1'd0}, _EVAL_625};
  assign _EVAL_268 = {_EVAL_354,_EVAL_92};
  assign _EVAL_207 = _EVAL_247 >= _EVAL_595;
  assign _EVAL_591 = {{1'd0}, _EVAL_161};
  assign _EVAL_756 = _EVAL_589 >= _EVAL_192;
  assign _EVAL_887 = _EVAL_806 >= _EVAL_509;
  assign _EVAL_163 = _EVAL_261 ? {{1'd0}, _EVAL_580} : _EVAL_150;
  assign _EVAL_657 = _EVAL_650 ? {{1'd0}, _EVAL_469} : _EVAL_811;
  assign _EVAL_241 = {{1'd0}, _EVAL_767};
  assign _EVAL_628 = 2'h2 | _EVAL_785;
  assign _EVAL_227 = _EVAL_48[13];
  assign _EVAL_265 = _EVAL_804 ? _EVAL_872 : _EVAL_257;
  assign _EVAL_342 = {_EVAL_279,_EVAL_77};
  assign _EVAL_717 = _EVAL_308 ? _EVAL_699 : _EVAL_494;
  assign _EVAL_463 = _EVAL_48[38];
  assign _EVAL_841 = _EVAL_611 >= _EVAL_678;
  assign _EVAL_131 = _EVAL_48[40];
  assign _EVAL_641 = {{1'd0}, _EVAL_445};
  assign _EVAL_231 = _EVAL_557 >= _EVAL_236;
  assign _EVAL_742 = _EVAL_230 >= _EVAL_232;
  assign _EVAL_298 = _EVAL_48[54];
  assign _EVAL_222 = {{1'd0}, _EVAL_437};
  assign _EVAL_801 = 2'h2 | _EVAL_591;
  assign _EVAL_333 = {_EVAL_148,_EVAL_13};
  assign _EVAL_171 = 2'h2 | _EVAL_594;
  assign _EVAL_635 = {_EVAL_726,_EVAL_101};
  assign _EVAL_505 = _EVAL_130 ? _EVAL_572 : _EVAL_326;
  assign _EVAL_724 = {_EVAL_351,_EVAL_116};
  assign _EVAL_242 = {_EVAL_643,_EVAL_26};
  assign _EVAL_602 = 5'h10 | _EVAL_690;
  assign _EVAL_246 = _EVAL_329 >= _EVAL_212;
  assign _EVAL_642 = _EVAL_485 >= _EVAL_631;
  assign _EVAL_360 = 2'h2 | _EVAL_862;
  assign _EVAL_177 = _EVAL_688 ? _EVAL_855 : _EVAL_566;
  assign _EVAL_276 = {_EVAL_851,_EVAL_114};
  assign _EVAL_455 = _EVAL_815 >= _EVAL_379;
  assign _EVAL_315 = {{1'd0}, _EVAL_211};
  assign _EVAL_849 = _EVAL_579 ? 1'h0 : 1'h1;
  assign _EVAL_367 = _EVAL_386 >= _EVAL_164;
  assign _EVAL_886 = _EVAL_666 ? {{1'd0}, _EVAL_741} : _EVAL_198;
  assign _EVAL_296 = {_EVAL_205,_EVAL_39};
  assign _EVAL_686 = _EVAL_780 >= _EVAL_616;
  assign _EVAL_370 = {_EVAL_357,_EVAL_79};
  assign _EVAL_234 = _EVAL_359 ? _EVAL_483 : _EVAL_441;
  assign _EVAL_408 = _EVAL_48[72];
  assign _EVAL_622 = _EVAL_48[69];
  assign _EVAL_361 = _EVAL_48[88];
  assign _EVAL_721 = {_EVAL_365,_EVAL_123};
  assign _EVAL_799 = _EVAL_48[125];
  assign _EVAL_723 = _EVAL_530 >= _EVAL_620;
  assign _EVAL_592 = {_EVAL_764,_EVAL_90};
  assign _EVAL_832 = 2'h2 | _EVAL_160;
  assign _EVAL_263 = _EVAL_364 ? _EVAL_242 : _EVAL_346;
  assign _EVAL_757 = {_EVAL_273,_EVAL_8};
  assign _EVAL_501 = 4'h8 | _EVAL_289;
  assign _EVAL_147 = 3'h4 | _EVAL_277;
  assign _EVAL_856 = 2'h2 | _EVAL_769;
  assign _EVAL_219 = _EVAL_429 ? _EVAL_239 : _EVAL_482;
  assign _EVAL_787 = _EVAL_578 >= _EVAL_313;
  assign _EVAL_477 = {{1'd0}, _EVAL_304};
  assign _EVAL_473 = _EVAL_722 ? _EVAL_176 : _EVAL_630;
  assign _EVAL_372 = _EVAL_364 ? 1'h0 : 1'h1;
  assign _EVAL_145 = _EVAL_610 ? _EVAL_552 : _EVAL_252;
  assign _EVAL_671 = {{1'd0}, _EVAL_159};
  assign _EVAL_883 = _EVAL_413 >= _EVAL_527;
  assign _EVAL_237 = _EVAL_865 ? _EVAL_542 : _EVAL_784;
  assign _EVAL_800 = _EVAL_597 >= _EVAL_500;
  assign _EVAL_434 = _EVAL_48[1];
  assign _EVAL_422 = {_EVAL_390,_EVAL_40};
  assign _EVAL_736 = _EVAL_367 ? 1'h0 : 1'h1;
  assign _EVAL_795 = _EVAL_151 >= _EVAL_166;
  assign _EVAL_698 = _EVAL_878 ? 1'h0 : 1'h1;
  assign _EVAL_656 = _EVAL_48[78];
  assign _EVAL_853 = _EVAL_343 ? {{1'd0}, _EVAL_657} : _EVAL_182;
  assign _EVAL_512 = _EVAL_798 ? _EVAL_813 : _EVAL_868;
  assign _EVAL_774 = 3'h4 | _EVAL_551;
endmodule
