//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_115(
  input         _EVAL,
  input  [29:0] _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input  [29:0] _EVAL_4,
  input  [31:0] _EVAL_5,
  output        _EVAL_6,
  output [1:0]  _EVAL_7,
  input  [2:0]  _EVAL_8,
  input  [31:0] _EVAL_9,
  output [4:0]  _EVAL_10,
  input         _EVAL_11,
  input  [31:0] _EVAL_12,
  input  [31:0] _EVAL_13,
  output [31:0] _EVAL_14,
  input         _EVAL_15,
  input  [31:0] _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18,
  output        _EVAL_19,
  output [31:0] _EVAL_20,
  input         _EVAL_21,
  input         _EVAL_22,
  input  [31:0] _EVAL_23,
  input  [1:0]  _EVAL_24,
  input         _EVAL_25,
  input  [1:0]  _EVAL_26,
  output        _EVAL_27,
  input  [31:0] _EVAL_28,
  input  [7:0]  _EVAL_29,
  input  [31:0] _EVAL_30,
  input  [29:0] _EVAL_31,
  input  [3:0]  _EVAL_32,
  input         _EVAL_33,
  input         _EVAL_34,
  input         _EVAL_35,
  input         _EVAL_36,
  input  [29:0] _EVAL_37,
  input  [31:0] _EVAL_38,
  output        _EVAL_39,
  input  [31:0] _EVAL_40,
  input         _EVAL_41,
  input         _EVAL_42,
  input  [4:0]  _EVAL_43,
  input  [29:0] _EVAL_44,
  input         _EVAL_45,
  input  [24:0] _EVAL_46,
  output        _EVAL_47,
  output        _EVAL_48,
  input         _EVAL_49,
  input         _EVAL_50,
  input  [31:0] _EVAL_51,
  input  [1:0]  _EVAL_52,
  input         _EVAL_53,
  input         _EVAL_54,
  input  [31:0] _EVAL_55,
  output        _EVAL_56,
  input         _EVAL_57,
  output [7:0]  _EVAL_58,
  input         _EVAL_59,
  input         _EVAL_60,
  input  [10:0] _EVAL_61,
  output [31:0] _EVAL_62,
  input  [1:0]  _EVAL_63,
  input         _EVAL_64,
  input         _EVAL_65,
  input         _EVAL_66,
  input         _EVAL_67,
  output        _EVAL_68,
  input  [31:0] _EVAL_69,
  input         _EVAL_70,
  input  [31:0] _EVAL_71,
  input  [3:0]  _EVAL_72,
  output [31:0] _EVAL_73,
  input  [2:0]  _EVAL_74,
  input         _EVAL_75,
  input  [29:0] _EVAL_76,
  input         _EVAL_77,
  input  [1:0]  _EVAL_78,
  input         _EVAL_79,
  input  [29:0] _EVAL_80,
  input         _EVAL_81,
  input         _EVAL_82,
  input         _EVAL_83,
  output [1:0]  _EVAL_84,
  input         _EVAL_85,
  output [10:0] _EVAL_86,
  input  [29:0] _EVAL_87,
  input         _EVAL_88,
  input         _EVAL_89,
  input  [1:0]  _EVAL_90,
  input         _EVAL_91,
  input  [31:0] _EVAL_92,
  input         _EVAL_93,
  input  [1:0]  _EVAL_94,
  input         _EVAL_95,
  input         _EVAL_96,
  input         _EVAL_97,
  output        _EVAL_98,
  output        _EVAL_99,
  input         _EVAL_100,
  output        _EVAL_101,
  input  [31:0] _EVAL_102,
  output [31:0] _EVAL_103,
  input         _EVAL_104,
  output [2:0]  _EVAL_105,
  input         _EVAL_106,
  input  [1:0]  _EVAL_107,
  input  [1:0]  _EVAL_108,
  input  [31:0] _EVAL_109,
  input  [1:0]  _EVAL_110,
  output        _EVAL_111,
  output        _EVAL_112,
  input         _EVAL_113,
  input         _EVAL_114,
  input  [1:0]  _EVAL_115,
  input         _EVAL_116,
  input         _EVAL_117,
  input         _EVAL_118,
  input         _EVAL_119,
  input         _EVAL_120
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] _EVAL_121;
  wire [1:0] _EVAL_122;
  wire  _EVAL_123;
  wire [20:0] _EVAL_124;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire [32:0] _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire [4:0] _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire [9:0] _EVAL_148;
  wire [1:0] _EVAL_149;
  wire  _EVAL_150;
  wire [32:0] _EVAL_151;
  wire [31:0] _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire [31:0] _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire [32:0] _EVAL_159;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire [33:0] _EVAL_163;
  wire [7:0] _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire [15:0] _EVAL_170;
  wire  _EVAL_171;
  wire [31:0] _EVAL_172;
  wire [1:0] _EVAL_173;
  wire [31:0] _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire [31:0] _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire [4:0] _EVAL_190;
  wire [15:0] _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire [31:0] _EVAL_197;
  wire [7:0] _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire [4:0] _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire [1:0] _EVAL_204;
  wire [4:0] _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_212;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire [20:0] _EVAL_217;
  reg  _EVAL_218;
  wire  _EVAL_219;
  wire [5:0] _EVAL_220;
  wire  _EVAL_221;
  wire [31:0] _EVAL_222;
  wire  _EVAL_223;
  wire [2:0] _EVAL_224;
  wire [31:0] _EVAL_225;
  wire [6:0] _EVAL_226;
  wire [4:0] _EVAL_227;
  wire  _EVAL_228;
  wire [32:0] _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_235;
  wire [31:0] _EVAL_236;
  wire  _EVAL_237;
  wire [32:0] _EVAL_239;
  wire [1:0] _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire [4:0] _EVAL_243;
  wire [31:0] _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire [15:0] _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_253;
  wire [3:0] _EVAL_254;
  wire  _EVAL_255;
  wire [31:0] _EVAL_256;
  wire [4:0] _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire [1:0] _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire [12:0] _EVAL_265;
  wire  _EVAL_266;
  wire [4:0] _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire [31:0] _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire [4:0] _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire [10:0] _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire  _EVAL_293;
  wire [32:0] _EVAL_294;
  wire [1:0] _EVAL_295;
  wire [1:0] _EVAL_296;
  wire [1:0] _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire [7:0] _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_307;
  wire [15:0] _EVAL_308;
  wire  _EVAL_309;
  wire  _EVAL_310;
  wire [6:0] _EVAL_311;
  wire  _EVAL_312;
  wire [4:0] _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_315;
  wire [15:0] _EVAL_317;
  wire [2:0] _EVAL_318;
  wire  _EVAL_319;
  wire [31:0] _EVAL_320;
  wire [32:0] _EVAL_321;
  wire  _EVAL_322;
  wire  _EVAL_323;
  wire [32:0] _EVAL_324;
  wire  _EVAL_325;
  wire  _EVAL_326;
  wire [15:0] _EVAL_327;
  wire  _EVAL_328;
  wire  _EVAL_329;
  wire [7:0] _EVAL_330;
  wire  _EVAL_331;
  wire  _EVAL_332;
  wire  _EVAL_333;
  wire  _EVAL_335;
  wire  _EVAL_336;
  wire  _EVAL_338;
  wire  _EVAL_339;
  wire  _EVAL_340;
  wire [31:0] _EVAL_344;
  wire  _EVAL_345;
  wire  _EVAL_346;
  wire  tlb__EVAL;
  wire  tlb__EVAL_0;
  wire  tlb__EVAL_1;
  wire [31:0] tlb__EVAL_2;
  wire [1:0] tlb__EVAL_3;
  wire [29:0] tlb__EVAL_4;
  wire  tlb__EVAL_5;
  wire [31:0] tlb__EVAL_6;
  wire  tlb__EVAL_7;
  wire [31:0] tlb__EVAL_8;
  wire  tlb__EVAL_9;
  wire [31:0] tlb__EVAL_10;
  wire  tlb__EVAL_11;
  wire  tlb__EVAL_12;
  wire  tlb__EVAL_13;
  wire [31:0] tlb__EVAL_14;
  wire  tlb__EVAL_15;
  wire  tlb__EVAL_16;
  wire  tlb__EVAL_17;
  wire  tlb__EVAL_18;
  wire  tlb__EVAL_19;
  wire [1:0] tlb__EVAL_20;
  wire  tlb__EVAL_21;
  wire [29:0] tlb__EVAL_22;
  wire [1:0] tlb__EVAL_23;
  wire  tlb__EVAL_24;
  wire  tlb__EVAL_25;
  wire  tlb__EVAL_26;
  wire  tlb__EVAL_27;
  wire  tlb__EVAL_28;
  wire  tlb__EVAL_29;
  wire [29:0] tlb__EVAL_30;
  wire [29:0] tlb__EVAL_31;
  wire [1:0] tlb__EVAL_32;
  wire  tlb__EVAL_33;
  wire  tlb__EVAL_34;
  wire [31:0] tlb__EVAL_35;
  wire [1:0] tlb__EVAL_36;
  wire [29:0] tlb__EVAL_37;
  wire [1:0] tlb__EVAL_38;
  wire [31:0] tlb__EVAL_39;
  wire  tlb__EVAL_40;
  wire  tlb__EVAL_41;
  wire  tlb__EVAL_42;
  wire  tlb__EVAL_43;
  wire  tlb__EVAL_44;
  wire [31:0] tlb__EVAL_45;
  wire  tlb__EVAL_46;
  wire [31:0] tlb__EVAL_47;
  wire  tlb__EVAL_48;
  wire [1:0] tlb__EVAL_49;
  wire  tlb__EVAL_50;
  wire  tlb__EVAL_51;
  wire  tlb__EVAL_52;
  wire [1:0] tlb__EVAL_53;
  wire  tlb__EVAL_54;
  wire [31:0] tlb__EVAL_55;
  wire  tlb__EVAL_56;
  wire [1:0] tlb__EVAL_57;
  wire [29:0] tlb__EVAL_58;
  wire  tlb__EVAL_59;
  wire [29:0] tlb__EVAL_60;
  wire [29:0] tlb__EVAL_61;
  wire  _EVAL_347;
  wire  _EVAL_348;
  wire  _EVAL_349;
  wire  _EVAL_350;
  wire [31:0] _EVAL_351;
  wire [20:0] _EVAL_352;
  wire  _EVAL_353;
  wire [7:0] _EVAL_354;
  wire [2:0] _EVAL_355;
  wire  _EVAL_356;
  wire  _EVAL_357;
  wire  _EVAL_358;
  wire [1:0] _EVAL_359;
  wire  _EVAL_360;
  wire  _EVAL_361;
  wire  _EVAL_362;
  wire [31:0] _EVAL_363;
  wire  _EVAL_365;
  wire  _EVAL_366;
  wire  _EVAL_367;
  wire  _EVAL_368;
  wire  _EVAL_369;
  wire  _EVAL_370;
  wire [32:0] _EVAL_371;
  wire  _EVAL_372;
  wire [20:0] _EVAL_373;
  wire  _EVAL_374;
  wire  _EVAL_375;
  wire  _EVAL_376;
  wire  _EVAL_377;
  wire  _EVAL_378;
  wire  _EVAL_379;
  wire  _EVAL_380;
  wire  _EVAL_381;
  wire  _EVAL_382;
  wire  _EVAL_383;
  wire  _EVAL_384;
  wire  _EVAL_385;
  wire [10:0] _EVAL_386;
  wire [4:0] _EVAL_387;
  wire  _EVAL_388;
  wire [32:0] _EVAL_389;
  wire [15:0] _EVAL_390;
  wire [31:0] btb__EVAL;
  wire  btb__EVAL_0;
  wire  btb__EVAL_1;
  wire  btb__EVAL_2;
  wire [31:0] btb__EVAL_3;
  wire  btb__EVAL_4;
  wire  btb__EVAL_5;
  wire  btb__EVAL_6;
  wire [1:0] btb__EVAL_7;
  wire [1:0] btb__EVAL_8;
  wire [31:0] btb__EVAL_9;
  wire  btb__EVAL_10;
  wire  btb__EVAL_11;
  wire  btb__EVAL_12;
  wire [31:0] btb__EVAL_13;
  wire  btb__EVAL_14;
  wire [31:0] btb__EVAL_15;
  wire [7:0] btb__EVAL_16;
  wire  btb__EVAL_17;
  wire [4:0] btb__EVAL_18;
  wire  btb__EVAL_19;
  wire  btb__EVAL_20;
  wire [31:0] btb__EVAL_21;
  wire  btb__EVAL_22;
  wire  btb__EVAL_23;
  wire [4:0] btb__EVAL_24;
  wire [7:0] btb__EVAL_25;
  wire  btb__EVAL_26;
  wire [31:0] btb__EVAL_27;
  wire  btb__EVAL_28;
  wire  _EVAL_392;
  wire  _EVAL_393;
  wire [1:0] _EVAL_394;
  wire [31:0] _EVAL_396;
  wire  _EVAL_397;
  wire  _EVAL_398;
  wire  _EVAL_399;
  wire  _EVAL_400;
  wire  _EVAL_401;
  wire [31:0] _EVAL_402;
  wire [2:0] _EVAL_403;
  wire  _EVAL_404;
  wire  _EVAL_405;
  wire [4:0] _EVAL_406;
  wire  _EVAL_407;
  wire [31:0] _EVAL_408;
  wire [1:0] _EVAL_409;
  wire  _EVAL_411;
  wire  _EVAL_412;
  wire  _EVAL_413;
  wire [31:0] _EVAL_414;
  wire [32:0] _EVAL_415;
  wire [10:0] _EVAL_416;
  wire  _EVAL_417;
  wire  _EVAL_418;
  wire  _EVAL_419;
  wire  _EVAL_420;
  wire  _EVAL_421;
  wire [31:0] _EVAL_423;
  wire [1:0] _EVAL_424;
  wire [1:0] _EVAL_425;
  wire  _EVAL_426;
  wire [31:0] _EVAL_427;
  wire [1:0] fq__EVAL;
  wire  fq__EVAL_0;
  wire  fq__EVAL_1;
  wire  fq__EVAL_2;
  wire  fq__EVAL_3;
  wire  fq__EVAL_4;
  wire  fq__EVAL_5;
  wire  fq__EVAL_6;
  wire [31:0] fq__EVAL_7;
  wire [1:0] fq__EVAL_8;
  wire [7:0] fq__EVAL_9;
  wire [4:0] fq__EVAL_10;
  wire  fq__EVAL_11;
  wire  fq__EVAL_12;
  wire  fq__EVAL_13;
  wire  fq__EVAL_14;
  wire  fq__EVAL_15;
  wire [31:0] fq__EVAL_16;
  wire  fq__EVAL_17;
  wire [31:0] fq__EVAL_18;
  wire  fq__EVAL_19;
  wire [4:0] fq__EVAL_20;
  wire [31:0] fq__EVAL_21;
  wire [4:0] fq__EVAL_22;
  wire [7:0] fq__EVAL_23;
  wire  _EVAL_428;
  wire  _EVAL_429;
  wire [1:0] _EVAL_430;
  wire  _EVAL_431;
  wire  _EVAL_432;
  wire  _EVAL_433;
  wire  _EVAL_434;
  wire  _EVAL_435;
  wire [32:0] _EVAL_436;
  wire [3:0] _EVAL_437;
  wire  _EVAL_438;
  wire  _EVAL_439;
  wire  _EVAL_440;
  wire  _EVAL_441;
  wire [7:0] _EVAL_442;
  wire [12:0] _EVAL_443;
  wire [7:0] _EVAL_444;
  wire  _EVAL_445;
  wire [32:0] _EVAL_446;
  wire  _EVAL_447;
  wire [31:0] _EVAL_449;
  wire  _EVAL_450;
  wire  _EVAL_452;
  wire  _EVAL_453;
  wire  _EVAL_454;
  wire [4:0] _EVAL_455;
  wire [31:0] _EVAL_456;
  wire  _EVAL_457;
  wire  _EVAL_458;
  wire  _EVAL_459;
  wire [31:0] _EVAL_460;
  wire  _EVAL_461;
  wire  _EVAL_462;
  wire  _EVAL_463;
  wire  _EVAL_464;
  wire  icache__EVAL;
  wire  icache__EVAL_0;
  wire  icache__EVAL_1;
  wire  icache__EVAL_2;
  wire  icache__EVAL_3;
  wire  icache__EVAL_4;
  wire  icache__EVAL_5;
  wire  icache__EVAL_6;
  wire [31:0] icache__EVAL_7;
  wire [3:0] icache__EVAL_8;
  wire [1:0] icache__EVAL_9;
  wire  icache__EVAL_10;
  wire [10:0] icache__EVAL_11;
  wire  icache__EVAL_12;
  wire  icache__EVAL_13;
  wire [31:0] icache__EVAL_14;
  wire [31:0] icache__EVAL_15;
  wire  icache__EVAL_16;
  wire  icache__EVAL_17;
  wire  icache__EVAL_18;
  wire  icache__EVAL_19;
  wire [1:0] icache__EVAL_20;
  wire  icache__EVAL_21;
  wire  icache__EVAL_22;
  wire  icache__EVAL_23;
  wire [24:0] icache__EVAL_24;
  wire  icache__EVAL_25;
  wire [3:0] icache__EVAL_26;
  wire [31:0] icache__EVAL_27;
  wire [2:0] icache__EVAL_28;
  wire [10:0] icache__EVAL_29;
  wire [31:0] icache__EVAL_30;
  wire [2:0] icache__EVAL_31;
  wire [31:0] icache__EVAL_32;
  wire [31:0] icache__EVAL_33;
  wire  icache__EVAL_34;
  wire  icache__EVAL_35;
  wire [31:0] icache__EVAL_36;
  wire [2:0] icache__EVAL_37;
  wire [10:0] _EVAL_465;
  wire [3:0] _EVAL_466;
  wire  _EVAL_467;
  wire  _EVAL_468;
  wire  _EVAL_470;
  wire  _EVAL_471;
  wire  _EVAL_472;
  wire [31:0] _EVAL_473;
  wire  _EVAL_474;
  wire  _EVAL_475;
  wire [20:0] _EVAL_476;
  wire  _EVAL_477;
  wire  _EVAL_478;
  wire  _EVAL_479;
  wire [32:0] _EVAL_480;
  wire [7:0] _EVAL_481;
  wire  _EVAL_482;
  wire  _EVAL_483;
  wire  _EVAL_484;
  wire  _EVAL_485;
  wire  _EVAL_486;
  wire [32:0] _EVAL_487;
  wire [32:0] _EVAL_488;
  wire  _EVAL_489;
  wire [9:0] _EVAL_490;
  wire [31:0] _EVAL_491;
  wire  _EVAL_492;
  wire  _EVAL_493;
  wire  _EVAL_494;
  wire  _EVAL_495;
  wire [32:0] _EVAL_496;
  wire  _EVAL_497;
  wire [12:0] _EVAL_498;
  wire  _EVAL_499;
  wire [7:0] _EVAL_500;
  wire [32:0] _EVAL_501;
  wire [31:0] _EVAL_502;
  wire [31:0] _EVAL_503;
  wire  _EVAL_504;
  wire [1:0] _EVAL_505;
  wire  _EVAL_506;
  wire  _EVAL_507;
  wire [20:0] _EVAL_508;
  wire  _EVAL_509;
  wire [32:0] _EVAL_510;
  wire  _EVAL_511;
  wire [7:0] _EVAL_513;
  wire [32:0] _EVAL_514;
  wire [31:0] _EVAL_515;
  wire  _EVAL_516;
  wire  _EVAL_517;
  wire [5:0] _EVAL_518;
  wire [1:0] _EVAL_519;
  wire [12:0] _EVAL_521;
  wire [31:0] _EVAL_522;
  wire  _EVAL_524;
  wire  _EVAL_525;
  wire  _EVAL_526;
  wire  _EVAL_527;
  wire  _EVAL_528;
  wire  _EVAL_529;
  wire  _EVAL_530;
  wire  _EVAL_531;
  wire  _EVAL_532;
  wire  _EVAL_533;
  wire  _EVAL_534;
  wire  _EVAL_536;
  wire  _EVAL_537;
  wire  _EVAL_538;
  wire [32:0] _EVAL_539;
  wire [31:0] _EVAL_540;
  wire  _EVAL_541;
  wire  _EVAL_542;
  wire  _EVAL_543;
  wire  _EVAL_545;
  wire  _EVAL_546;
  wire  _EVAL_548;
  wire  _EVAL_549;
  wire  gated_clock_icache_clock_gate_in;
  wire  gated_clock_icache_clock_gate_test_en;
  wire  gated_clock_icache_clock_gate_en;
  wire  gated_clock_icache_clock_gate_out;
  reg  _EVAL_550;
  reg  _EVAL_551;
  reg  _EVAL_552;
  reg  _EVAL_553;
  reg [15:0] _EVAL_554;
  reg  _EVAL_555;
  reg  _EVAL_556;
  reg [31:0] _EVAL_557;
  reg [31:0] _EVAL_558;
  reg [7:0] _EVAL_559;
  reg  _EVAL_560;
  reg  _EVAL_561;
  reg  _EVAL_562;
  reg [4:0] _EVAL_563;
  reg  _EVAL_564;
  reg  _EVAL_565;
  reg  _EVAL_566;
  reg  _EVAL_567;
  wire [31:0] _EVAL_568;
  wire  _EVAL_570;
  wire  _EVAL_571;
  wire  _EVAL_572;
  wire  _EVAL_573;
  wire  _EVAL_574;
  wire [31:0] _EVAL_575;
  wire [3:0] _EVAL_576;
  _EVAL_113 tlb (
    ._EVAL(tlb__EVAL),
    ._EVAL_0(tlb__EVAL_0),
    ._EVAL_1(tlb__EVAL_1),
    ._EVAL_2(tlb__EVAL_2),
    ._EVAL_3(tlb__EVAL_3),
    ._EVAL_4(tlb__EVAL_4),
    ._EVAL_5(tlb__EVAL_5),
    ._EVAL_6(tlb__EVAL_6),
    ._EVAL_7(tlb__EVAL_7),
    ._EVAL_8(tlb__EVAL_8),
    ._EVAL_9(tlb__EVAL_9),
    ._EVAL_10(tlb__EVAL_10),
    ._EVAL_11(tlb__EVAL_11),
    ._EVAL_12(tlb__EVAL_12),
    ._EVAL_13(tlb__EVAL_13),
    ._EVAL_14(tlb__EVAL_14),
    ._EVAL_15(tlb__EVAL_15),
    ._EVAL_16(tlb__EVAL_16),
    ._EVAL_17(tlb__EVAL_17),
    ._EVAL_18(tlb__EVAL_18),
    ._EVAL_19(tlb__EVAL_19),
    ._EVAL_20(tlb__EVAL_20),
    ._EVAL_21(tlb__EVAL_21),
    ._EVAL_22(tlb__EVAL_22),
    ._EVAL_23(tlb__EVAL_23),
    ._EVAL_24(tlb__EVAL_24),
    ._EVAL_25(tlb__EVAL_25),
    ._EVAL_26(tlb__EVAL_26),
    ._EVAL_27(tlb__EVAL_27),
    ._EVAL_28(tlb__EVAL_28),
    ._EVAL_29(tlb__EVAL_29),
    ._EVAL_30(tlb__EVAL_30),
    ._EVAL_31(tlb__EVAL_31),
    ._EVAL_32(tlb__EVAL_32),
    ._EVAL_33(tlb__EVAL_33),
    ._EVAL_34(tlb__EVAL_34),
    ._EVAL_35(tlb__EVAL_35),
    ._EVAL_36(tlb__EVAL_36),
    ._EVAL_37(tlb__EVAL_37),
    ._EVAL_38(tlb__EVAL_38),
    ._EVAL_39(tlb__EVAL_39),
    ._EVAL_40(tlb__EVAL_40),
    ._EVAL_41(tlb__EVAL_41),
    ._EVAL_42(tlb__EVAL_42),
    ._EVAL_43(tlb__EVAL_43),
    ._EVAL_44(tlb__EVAL_44),
    ._EVAL_45(tlb__EVAL_45),
    ._EVAL_46(tlb__EVAL_46),
    ._EVAL_47(tlb__EVAL_47),
    ._EVAL_48(tlb__EVAL_48),
    ._EVAL_49(tlb__EVAL_49),
    ._EVAL_50(tlb__EVAL_50),
    ._EVAL_51(tlb__EVAL_51),
    ._EVAL_52(tlb__EVAL_52),
    ._EVAL_53(tlb__EVAL_53),
    ._EVAL_54(tlb__EVAL_54),
    ._EVAL_55(tlb__EVAL_55),
    ._EVAL_56(tlb__EVAL_56),
    ._EVAL_57(tlb__EVAL_57),
    ._EVAL_58(tlb__EVAL_58),
    ._EVAL_59(tlb__EVAL_59),
    ._EVAL_60(tlb__EVAL_60),
    ._EVAL_61(tlb__EVAL_61)
  );
  _EVAL_114 btb (
    ._EVAL(btb__EVAL),
    ._EVAL_0(btb__EVAL_0),
    ._EVAL_1(btb__EVAL_1),
    ._EVAL_2(btb__EVAL_2),
    ._EVAL_3(btb__EVAL_3),
    ._EVAL_4(btb__EVAL_4),
    ._EVAL_5(btb__EVAL_5),
    ._EVAL_6(btb__EVAL_6),
    ._EVAL_7(btb__EVAL_7),
    ._EVAL_8(btb__EVAL_8),
    ._EVAL_9(btb__EVAL_9),
    ._EVAL_10(btb__EVAL_10),
    ._EVAL_11(btb__EVAL_11),
    ._EVAL_12(btb__EVAL_12),
    ._EVAL_13(btb__EVAL_13),
    ._EVAL_14(btb__EVAL_14),
    ._EVAL_15(btb__EVAL_15),
    ._EVAL_16(btb__EVAL_16),
    ._EVAL_17(btb__EVAL_17),
    ._EVAL_18(btb__EVAL_18),
    ._EVAL_19(btb__EVAL_19),
    ._EVAL_20(btb__EVAL_20),
    ._EVAL_21(btb__EVAL_21),
    ._EVAL_22(btb__EVAL_22),
    ._EVAL_23(btb__EVAL_23),
    ._EVAL_24(btb__EVAL_24),
    ._EVAL_25(btb__EVAL_25),
    ._EVAL_26(btb__EVAL_26),
    ._EVAL_27(btb__EVAL_27),
    ._EVAL_28(btb__EVAL_28)
  );
  _EVAL_112 fq (
    ._EVAL(fq__EVAL),
    ._EVAL_0(fq__EVAL_0),
    ._EVAL_1(fq__EVAL_1),
    ._EVAL_2(fq__EVAL_2),
    ._EVAL_3(fq__EVAL_3),
    ._EVAL_4(fq__EVAL_4),
    ._EVAL_5(fq__EVAL_5),
    ._EVAL_6(fq__EVAL_6),
    ._EVAL_7(fq__EVAL_7),
    ._EVAL_8(fq__EVAL_8),
    ._EVAL_9(fq__EVAL_9),
    ._EVAL_10(fq__EVAL_10),
    ._EVAL_11(fq__EVAL_11),
    ._EVAL_12(fq__EVAL_12),
    ._EVAL_13(fq__EVAL_13),
    ._EVAL_14(fq__EVAL_14),
    ._EVAL_15(fq__EVAL_15),
    ._EVAL_16(fq__EVAL_16),
    ._EVAL_17(fq__EVAL_17),
    ._EVAL_18(fq__EVAL_18),
    ._EVAL_19(fq__EVAL_19),
    ._EVAL_20(fq__EVAL_20),
    ._EVAL_21(fq__EVAL_21),
    ._EVAL_22(fq__EVAL_22),
    ._EVAL_23(fq__EVAL_23)
  );
  _EVAL_111 icache (
    ._EVAL(icache__EVAL),
    ._EVAL_0(icache__EVAL_0),
    ._EVAL_1(icache__EVAL_1),
    ._EVAL_2(icache__EVAL_2),
    ._EVAL_3(icache__EVAL_3),
    ._EVAL_4(icache__EVAL_4),
    ._EVAL_5(icache__EVAL_5),
    ._EVAL_6(icache__EVAL_6),
    ._EVAL_7(icache__EVAL_7),
    ._EVAL_8(icache__EVAL_8),
    ._EVAL_9(icache__EVAL_9),
    ._EVAL_10(icache__EVAL_10),
    ._EVAL_11(icache__EVAL_11),
    ._EVAL_12(icache__EVAL_12),
    ._EVAL_13(icache__EVAL_13),
    ._EVAL_14(icache__EVAL_14),
    ._EVAL_15(icache__EVAL_15),
    ._EVAL_16(icache__EVAL_16),
    ._EVAL_17(icache__EVAL_17),
    ._EVAL_18(icache__EVAL_18),
    ._EVAL_19(icache__EVAL_19),
    ._EVAL_20(icache__EVAL_20),
    ._EVAL_21(icache__EVAL_21),
    ._EVAL_22(icache__EVAL_22),
    ._EVAL_23(icache__EVAL_23),
    ._EVAL_24(icache__EVAL_24),
    ._EVAL_25(icache__EVAL_25),
    ._EVAL_26(icache__EVAL_26),
    ._EVAL_27(icache__EVAL_27),
    ._EVAL_28(icache__EVAL_28),
    ._EVAL_29(icache__EVAL_29),
    ._EVAL_30(icache__EVAL_30),
    ._EVAL_31(icache__EVAL_31),
    ._EVAL_32(icache__EVAL_32),
    ._EVAL_33(icache__EVAL_33),
    ._EVAL_34(icache__EVAL_34),
    ._EVAL_35(icache__EVAL_35),
    ._EVAL_36(icache__EVAL_36),
    ._EVAL_37(icache__EVAL_37)
  );
  EICG_wrapper gated_clock_icache_clock_gate (
    .in(gated_clock_icache_clock_gate_in),
    .test_en(gated_clock_icache_clock_gate_test_en),
    .en(gated_clock_icache_clock_gate_en),
    .out(gated_clock_icache_clock_gate_out)
  );
  assign _EVAL_532 = _EVAL_327[8];
  assign _EVAL_465 = _EVAL_416;
  assign _EVAL_515 = _EVAL_484 ? btb__EVAL_3 : _EVAL_402;
  assign _EVAL_321 = $signed(_EVAL_197) + $signed(_EVAL_172);
  assign icache__EVAL_2 = _EVAL_464 | _EVAL_276;
  assign _EVAL_313 = _EVAL_363[19:15];
  assign _EVAL_519 = _EVAL_157 ? 2'h2 : {{1'd0}, _EVAL_196};
  assign _EVAL_279 = _EVAL_202 & _EVAL_541;
  assign _EVAL_528 = _EVAL_555 & _EVAL_556;
  assign _EVAL_241 = _EVAL_572 | _EVAL_564;
  assign tlb__EVAL_15 = _EVAL_82;
  assign _EVAL_331 = fq__EVAL_11 & fq__EVAL_5;
  assign _EVAL_311 = _EVAL_363[6:0];
  assign _EVAL_308 = _EVAL_327 & 16'he003;
  assign _EVAL_503 = _EVAL_522 | 32'h2;
  assign _EVAL_273 = _EVAL_251 & _EVAL_440;
  assign _EVAL_346 = btb__EVAL_19 & _EVAL_463;
  assign _EVAL_437 = _EVAL_363[11:8];
  assign tlb__EVAL_26 = _EVAL_11;
  assign _EVAL_573 = _EVAL_405;
  assign _EVAL_318 = _EVAL_390[5:3];
  assign _EVAL_325 = _EVAL_495 & _EVAL_420;
  assign _EVAL_298 = _EVAL_13[0];
  assign _EVAL_221 = ~_EVAL_421;
  assign _EVAL_138 = _EVAL_393 | _EVAL_484;
  assign tlb__EVAL_39 = _EVAL_558;
  assign tlb__EVAL_55 = _EVAL_12;
  assign _EVAL_359 = _EVAL_390[11:10];
  assign _EVAL_163 = $signed(_EVAL_436) + $signed(_EVAL_539);
  assign _EVAL_463 = _EVAL_279 | _EVAL_249;
  assign _EVAL_454 = _EVAL_555 & _EVAL_326;
  assign _EVAL_58 = fq__EVAL_23;
  assign _EVAL_249 = _EVAL_288 & _EVAL_474;
  assign _EVAL_227 = _EVAL_455 & 5'h1b;
  assign _EVAL_126 = _EVAL_299;
  assign _EVAL_295 = _EVAL_390[1:0];
  assign _EVAL_145 = _EVAL_571 & _EVAL_129;
  assign _EVAL_179 = ~_EVAL_69;
  assign _EVAL_291 = _EVAL_132 & _EVAL_322;
  assign _EVAL_175 = _EVAL_153 | _EVAL_367;
  assign tlb__EVAL_27 = _EVAL_91;
  assign tlb__EVAL_31 = _EVAL_31;
  assign _EVAL_350 = _EVAL_129 & _EVAL_479;
  assign _EVAL_369 = _EVAL_289 | _EVAL_181;
  assign tlb__EVAL_10 = _EVAL_30;
  assign _EVAL_194 = _EVAL_275 & _EVAL_561;
  assign _EVAL_518 = _EVAL_363[30:25];
  assign _EVAL_256 = _EVAL_321[31:0];
  assign _EVAL_413 = _EVAL_555 & _EVAL_346;
  assign tlb__EVAL_14 = _EVAL_28;
  assign _EVAL_224 = _EVAL_327[5:3];
  assign _EVAL_143 = _EVAL_168 | _EVAL_493;
  assign tlb__EVAL_56 = _EVAL_42;
  assign _EVAL_200 = _EVAL_363[7];
  assign _EVAL_276 = _EVAL_315 | _EVAL_550;
  assign _EVAL_404 = 16'h8002 == _EVAL_191;
  assign _EVAL_235 = _EVAL_137 & _EVAL_319;
  assign btb__EVAL_21 = _EVAL_558;
  assign _EVAL_478 = _EVAL_222[20];
  assign tlb__EVAL_45 = _EVAL_16;
  assign _EVAL_530 = _EVAL_390[8];
  assign _EVAL_137 = ~_EVAL_165;
  assign _EVAL_492 = _EVAL_323 & _EVAL_447;
  assign _EVAL_509 = _EVAL_129 & _EVAL_329;
  assign _EVAL_287 = _EVAL_182;
  assign _EVAL_124 = {_EVAL_148,_EVAL_532,_EVAL_424,_EVAL_312,_EVAL_365,_EVAL_259,_EVAL_144,_EVAL_224,1'h0};
  assign _EVAL_261 = _EVAL_188 | _EVAL_382;
  assign _EVAL_158 = _EVAL_245 | _EVAL_216;
  assign _EVAL_431 = _EVAL_188 ? _EVAL_570 : _EVAL_567;
  assign _EVAL_502 = _EVAL_237 ? $signed(_EVAL_460) : $signed(_EVAL_456);
  assign icache__EVAL_20 = _EVAL_94;
  assign icache__EVAL_34 = _EVAL_77;
  assign _EVAL_297 = _EVAL_390[4:3];
  assign _EVAL_216 = _EVAL_399 & _EVAL_417;
  assign tlb__EVAL_59 = _EVAL_114;
  assign fq__EVAL_22 = _EVAL_453 ? _EVAL_133 : _EVAL_563;
  assign tlb__EVAL_57 = _EVAL_110;
  assign _EVAL_277 = _EVAL_307 ? 5'h1f : 5'h0;
  assign tlb__EVAL_48 = _EVAL_93;
  assign _EVAL_373 = {_EVAL_490,_EVAL_530,_EVAL_149,_EVAL_426,_EVAL_362,_EVAL_208,_EVAL_283,_EVAL_318,1'h0};
  assign _EVAL_495 = _EVAL_562 & _EVAL_193;
  assign _EVAL_317 = _EVAL_327 & 16'hf003;
  assign _EVAL_155 = ~icache__EVAL_21;
  assign _EVAL_205 = _EVAL_390[11:7];
  assign _EVAL_387 = _EVAL_290 ? 5'h1f : 5'h0;
  assign _EVAL_127 = _EVAL_495 & _EVAL_400;
  assign _EVAL_212 = _EVAL_166 | _EVAL_511;
  assign _EVAL_576 = _EVAL_222[11:8];
  assign _EVAL_390 = fq__EVAL_18[31:16];
  assign _EVAL_56 = fq__EVAL_6;
  assign _EVAL_377 = _EVAL_295 != 2'h3;
  assign _EVAL_98 = icache__EVAL_1;
  assign _EVAL_540 = ~_EVAL_558;
  assign _EVAL_328 = _EVAL_555 & _EVAL_260;
  assign _EVAL_400 = _EVAL_226 == 7'h63;
  assign _EVAL_20 = icache__EVAL_27;
  assign _EVAL_214 = _EVAL_435 | _EVAL_154;
  assign _EVAL_452 = _EVAL_228 & _EVAL_266;
  assign _EVAL_438 = _EVAL_331 & _EVAL_525;
  assign _EVAL_355 = {_EVAL_409, 1'h0};
  assign _EVAL_420 = _EVAL_226 == 7'h6f;
  assign _EVAL_39 = _EVAL_218 | _EVAL_104;
  assign _EVAL_533 = ~_EVAL_276;
  assign _EVAL_432 = _EVAL_561 | _EVAL_298;
  assign _EVAL_471 = _EVAL_292 | _EVAL_291;
  assign _EVAL_27 = fq__EVAL_12;
  assign _EVAL_14 = fq__EVAL_7;
  assign fq__EVAL_21 = _EVAL_557;
  assign _EVAL_152 = {_EVAL_304,_EVAL_465,_EVAL_302,_EVAL_287,_EVAL_518,_EVAL_466,1'h0};
  assign btb__EVAL_26 = _EVAL_15;
  assign _EVAL_299 = _EVAL_363[31];
  assign _EVAL_510 = _EVAL_130 ? _EVAL_389 : {{1'd0}, _EVAL_515};
  assign _EVAL_171 = _EVAL_384 & _EVAL_310;
  assign tlb__EVAL_37 = _EVAL_80;
  assign _EVAL_165 = fq__EVAL_10[3];
  assign _EVAL_574 = _EVAL_478;
  assign icache__EVAL_12 = _EVAL_97;
  assign _EVAL_497 = _EVAL_231 | _EVAL_509;
  assign _EVAL_534 = _EVAL_226 == 7'h67;
  assign _EVAL_548 = ~_EVAL_405;
  assign _EVAL_294 = _EVAL_300 ? {{1'd0}, btb__EVAL} : _EVAL_487;
  assign _EVAL_507 = _EVAL_551 & _EVAL_555;
  assign _EVAL_326 = _EVAL_275 | _EVAL_284;
  assign _EVAL_259 = _EVAL_327[2];
  assign tlb__EVAL_52 = _EVAL_89;
  assign btb__EVAL_12 = _EVAL_301 | _EVAL_113;
  assign tlb__EVAL_51 = _EVAL_119;
  assign _EVAL_482 = _EVAL_447 & _EVAL_366;
  assign _EVAL_248 = _EVAL_390 & 16'he003;
  assign _EVAL_445 = ~_EVAL_331;
  assign _EVAL_258 = _EVAL_327[6:2];
  assign _EVAL_197 = _EVAL_174;
  assign _EVAL_201 = _EVAL_190 & 5'h1b;
  assign _EVAL_290 = _EVAL_390[12];
  assign _EVAL_370 = _EVAL_288 & _EVAL_458;
  assign _EVAL_304 = _EVAL_126;
  assign _EVAL_517 = _EVAL_325 | _EVAL_264;
  assign _EVAL_281 = ~_EVAL_464;
  assign tlb__EVAL_23 = _EVAL_78;
  assign _EVAL_169 = _EVAL_363[20];
  assign _EVAL_251 = _EVAL_314 & _EVAL_288;
  assign _EVAL_86 = icache__EVAL_29;
  assign _EVAL_111 = icache__EVAL_23;
  assign _EVAL_84 = icache__EVAL_9;
  assign _EVAL_378 = _EVAL_181 & _EVAL_161;
  assign _EVAL_159 = ~_EVAL_151;
  assign btb__EVAL_0 = _EVAL_106;
  assign tlb__EVAL_25 = _EVAL_49;
  assign _EVAL_262 = _EVAL_554[1:0];
  assign _EVAL_539 = _EVAL_495 ? $signed(_EVAL_415) : $signed({{12{_EVAL_476[20]}},_EVAL_476});
  assign _EVAL_132 = 16'h8002 == _EVAL_317;
  assign tlb__EVAL_4 = _EVAL_37;
  assign _EVAL_455 = _EVAL_327[11:7];
  assign _EVAL_484 = btb__EVAL_2 & btb__EVAL_22;
  assign _EVAL_424 = _EVAL_327[10:9];
  assign _EVAL_225 = {{29'd0}, _EVAL_355};
  assign _EVAL_527 = ~_EVAL_517;
  assign _EVAL_338 = _EVAL_207 | _EVAL_517;
  assign _EVAL_464 = _EVAL_453 ? _EVAL_142 : _EVAL_18;
  assign tlb__EVAL_58 = _EVAL_76;
  assign _EVAL_498 = {_EVAL_387,_EVAL_173,_EVAL_208,_EVAL_359,_EVAL_297,1'h0};
  assign _EVAL_543 = fq__EVAL_10[2];
  assign _EVAL_367 = _EVAL_273 | _EVAL_332;
  assign _EVAL_419 = _EVAL_534 | _EVAL_420;
  assign _EVAL_457 = _EVAL_483 | _EVAL_235;
  assign _EVAL_353 = _EVAL_392 | _EVAL_136;
  assign _EVAL_237 = _EVAL_363[3];
  assign _EVAL_468 = 5'h1 == _EVAL_243;
  assign _EVAL_264 = _EVAL_129 & _EVAL_185;
  assign _EVAL_180 = 16'hc001 == _EVAL_308;
  assign _EVAL_229 = _EVAL_18 ? {{1'd0}, _EVAL_109} : _EVAL_496;
  assign icache__EVAL_24 = _EVAL_46;
  assign _EVAL_349 = _EVAL_223;
  assign _EVAL_136 = 16'h2001 == _EVAL_248;
  assign _EVAL_572 = _EVAL_104 | icache__EVAL_16;
  assign fq__EVAL_0 = _EVAL_77 | _EVAL_18;
  assign _EVAL_536 = _EVAL_390[14];
  assign _EVAL_459 = _EVAL_495 ? _EVAL_526 : _EVAL_140;
  assign btb__EVAL_6 = _EVAL_570 ? _EVAL_482 : _EVAL_339;
  assign _EVAL_195 = _EVAL_526 | _EVAL_485;
  assign _EVAL_570 = ~_EVAL_516;
  assign _EVAL_542 = _EVAL_306 | _EVAL_346;
  assign btb__EVAL_10 = _EVAL_273 | _EVAL_336;
  assign _EVAL_244 = {_EVAL_461,_EVAL_280,_EVAL_442,_EVAL_412,_EVAL_220,_EVAL_576,1'h0};
  assign _EVAL_458 = _EVAL_472 | _EVAL_474;
  assign tlb__EVAL_3 = _EVAL_115;
  assign btb__EVAL_8 = _EVAL_301 ? btb__EVAL_7 : _EVAL_26;
  assign _EVAL_356 = ~_EVAL_556;
  assign tlb__EVAL_29 = _EVAL_67;
  assign tlb__EVAL_30 = _EVAL_44;
  assign btb__EVAL_20 = _EVAL_570 ? _EVAL_135 : _EVAL_492;
  assign _EVAL_351 = _EVAL_540 | 32'h3;
  assign _EVAL_429 = _EVAL_288 & _EVAL_570;
  assign _EVAL_198 = _EVAL_164;
  assign icache__EVAL_11 = _EVAL_61;
  assign _EVAL_433 = icache__EVAL_21 & icache__EVAL_25;
  assign tlb__EVAL_6 = _EVAL_55;
  assign _EVAL_307 = _EVAL_327[12];
  assign icache__EVAL_32 = _EVAL_103;
  assign _EVAL_529 = _EVAL_420 | _EVAL_534;
  assign _EVAL_246 = 16'hc001 == _EVAL_248;
  assign _EVAL_474 = _EVAL_348 & _EVAL_531;
  assign btb__EVAL_9 = _EVAL_301 ? _EVAL_449 : _EVAL_5;
  assign _EVAL_329 = _EVAL_140 | _EVAL_167;
  assign _EVAL_403 = 3'h3 << _EVAL_134;
  assign _EVAL_531 = 5'h1 == _EVAL_267;
  assign _EVAL_191 = _EVAL_390 & 16'hf003;
  assign _EVAL_538 = _EVAL_438 & _EVAL_206;
  assign tlb__EVAL_0 = _EVAL_33;
  assign _EVAL_265 = _EVAL_521;
  assign tlb__EVAL_43 = _EVAL_88;
  assign _EVAL_376 = _EVAL_171 ? 1'h0 : 1'h1;
  assign icache__EVAL_19 = _EVAL_3;
  assign _EVAL_135 = _EVAL_199 ? _EVAL_447 : _EVAL_492;
  assign _EVAL_344 = ~_EVAL_396;
  assign _EVAL_220 = _EVAL_222[30:25];
  assign _EVAL_226 = _EVAL_222[6:0];
  assign _EVAL_333 = _EVAL_447 & _EVAL_282;
  assign _EVAL_374 = _EVAL_233 & _EVAL_432;
  assign _EVAL_481 = {8{_EVAL_475}};
  assign _EVAL_415 = $signed(_EVAL_568) - 32'sh2;
  assign icache__EVAL_8 = _EVAL_32;
  assign tlb__EVAL_61 = _EVAL_0;
  assign _EVAL_409 = _EVAL_570 ? 2'h2 : 2'h1;
  assign _EVAL_441 = _EVAL_333 & _EVAL_183;
  assign _EVAL_335 = _EVAL_222[31];
  assign _EVAL_306 = _EVAL_194 | _EVAL_284;
  assign _EVAL_493 = _EVAL_184 & _EVAL_432;
  assign _EVAL_571 = _EVAL_528 & _EVAL_268;
  assign _EVAL_405 = _EVAL_222[7];
  assign _EVAL_479 = _EVAL_471 | _EVAL_374;
  assign btb__EVAL_27 = _EVAL_40;
  assign tlb__EVAL_22 = _EVAL_87;
  assign _EVAL_435 = _EVAL_381 & _EVAL_215;
  assign _EVAL_48 = fq__EVAL_1;
  assign _EVAL_222 = {_EVAL_327,_EVAL_554};
  assign _EVAL_358 = 16'he001 == _EVAL_308;
  assign tlb__EVAL_24 = _EVAL_35;
  assign _EVAL_360 = _EVAL_338 | _EVAL_178;
  assign tlb__EVAL_8 = _EVAL_9;
  assign _EVAL_491 = ~_EVAL_557;
  assign _EVAL_368 = fq__EVAL[0];
  assign _EVAL_427 = ~_EVAL_351;
  assign tlb__EVAL_46 = _EVAL_17;
  assign _EVAL_189 = _EVAL_457 | _EVAL_209;
  assign tlb__EVAL_44 = _EVAL_75;
  assign _EVAL_219 = ~_EVAL_555;
  assign _EVAL_223 = _EVAL_200;
  assign _EVAL_263 = icache__EVAL_13;
  assign _EVAL_363 = {_EVAL_390,_EVAL_327};
  assign _EVAL_575 = _EVAL_256;
  assign _EVAL_233 = _EVAL_180 | _EVAL_358;
  assign tlb__EVAL_50 = _EVAL_81;
  assign _EVAL_151 = _EVAL_488 | 33'h1;
  assign tlb__EVAL_17 = _EVAL_77;
  assign _EVAL_384 = _EVAL_495 ? _EVAL_400 : _EVAL_233;
  assign fq__EVAL_9 = _EVAL_559;
  assign _EVAL_526 = _EVAL_419 & _EVAL_405;
  assign _EVAL_320 = _EVAL_491 | 32'h3;
  assign tlb__EVAL_19 = _EVAL_34;
  assign tlb__EVAL_32 = _EVAL_107;
  assign _EVAL_231 = _EVAL_495 & _EVAL_195;
  assign _EVAL_546 = icache__EVAL_21 | _EVAL_263;
  assign _EVAL_496 = _EVAL_276 ? {{1'd0}, _EVAL_557} : _EVAL_294;
  assign tlb__EVAL_53 = _EVAL_52;
  assign _EVAL_177 = fq__EVAL_10[4];
  assign _EVAL_521 = {_EVAL_277,_EVAL_505,_EVAL_259,_EVAL_430,_EVAL_296,1'h0};
  assign _EVAL_314 = _EVAL_528 & _EVAL_567;
  assign _EVAL_426 = _EVAL_390[6];
  assign tlb__EVAL_1 = _EVAL_95;
  assign _EVAL_275 = _EVAL_432 & _EVAL_199;
  assign _EVAL_366 = _EVAL_385 | _EVAL_370;
  assign _EVAL_511 = _EVAL_356 & _EVAL_360;
  assign _EVAL_123 = _EVAL_555 & _EVAL_178;
  assign _EVAL_173 = _EVAL_390[6:5];
  assign _EVAL_271 = {_EVAL_304,_EVAL_465,_EVAL_444,_EVAL_349,_EVAL_518,_EVAL_437,1'h0};
  assign _EVAL_253 = _EVAL_353 | _EVAL_452;
  assign tlb__EVAL_42 = gated_clock_icache_clock_gate_out;
  assign _EVAL_270 = _EVAL_222[3];
  assign _EVAL_442 = _EVAL_481;
  assign _EVAL_312 = _EVAL_327[6];
  assign _EVAL_164 = _EVAL_513;
  assign icache__EVAL_0 = _EVAL_116;
  assign _EVAL_389 = _EVAL_446;
  assign _EVAL_289 = _EVAL_311 == 7'h6f;
  assign _EVAL_247 = ~_EVAL_537;
  assign _EVAL_489 = _EVAL_331 & _EVAL_516;
  assign _EVAL_255 = _EVAL_369 | _EVAL_230;
  assign _EVAL_379 = _EVAL_429 & _EVAL_440;
  assign _EVAL_322 = _EVAL_258 == 5'h0;
  assign _EVAL_444 = _EVAL_500;
  assign _EVAL_105 = icache__EVAL_37;
  assign fq__EVAL_2 = _EVAL_100;
  assign _EVAL_398 = _EVAL_489 & _EVAL_221;
  assign _EVAL_310 = ~_EVAL_298;
  assign _EVAL_280 = _EVAL_386;
  assign fq__EVAL_18 = icache__EVAL_15;
  assign _EVAL_203 = _EVAL_534 & _EVAL_548;
  assign _EVAL_181 = _EVAL_311 == 7'h67;
  assign btb__EVAL_11 = _EVAL_77;
  assign _EVAL_184 = _EVAL_246 | _EVAL_477;
  assign _EVAL_99 = icache__EVAL;
  assign _EVAL_122 = _EVAL_347 ? 2'h3 : _EVAL_519;
  assign _EVAL_396 = _EVAL_179 | 32'h1;
  assign _EVAL_456 = _EVAL_271;
  assign _EVAL_372 = _EVAL_494 & _EVAL_310;
  assign _EVAL_156 = _EVAL_244;
  assign _EVAL_485 = _EVAL_203 & _EVAL_286;
  assign _EVAL_407 = ~_EVAL_553;
  assign _EVAL_154 = _EVAL_245 | _EVAL_553;
  assign _EVAL_153 = _EVAL_285 & _EVAL_131;
  assign _EVAL_250 = 16'h9002 == _EVAL_317;
  assign _EVAL_393 = _EVAL_566 | _EVAL_328;
  assign _EVAL_134 = _EVAL_557[1];
  assign _EVAL_514 = _EVAL_454 ? {{1'd0}, _EVAL_414} : _EVAL_324;
  assign _EVAL_149 = _EVAL_390[10:9];
  assign tlb__EVAL_18 = _EVAL_85;
  assign _EVAL_147 = _EVAL_574;
  assign _EVAL_157 = _EVAL_202 ? _EVAL_305 : _EVAL_472;
  assign tlb__EVAL_20 = _EVAL_63;
  assign btb__EVAL_25 = _EVAL_29;
  assign _EVAL_170 = _EVAL_390 | 16'h3;
  assign _EVAL_385 = _EVAL_202 & _EVAL_499;
  assign _EVAL_447 = _EVAL_331 & _EVAL_407;
  assign _EVAL_412 = _EVAL_573;
  assign gated_clock_icache_clock_gate_in = _EVAL_100;
  assign _EVAL_7 = fq__EVAL_8;
  assign _EVAL_440 = ~_EVAL_377;
  assign btb__EVAL_14 = _EVAL_561;
  assign _EVAL_232 = ~_EVAL_202;
  assign tlb__EVAL_41 = _EVAL_36;
  assign _EVAL_272 = _EVAL_276 & _EVAL_247;
  assign _EVAL_193 = ~_EVAL_139;
  assign tlb__EVAL_38 = _EVAL_24;
  assign icache__EVAL_4 = _EVAL_2;
  assign _EVAL_196 = _EVAL_372 ? 1'h0 : 1'h1;
  assign _EVAL_340 = 16'h2001 == _EVAL_308;
  assign icache__EVAL_10 = _EVAL_218 | _EVAL_104;
  assign _EVAL_545 = _EVAL_495 & _EVAL_401;
  assign _EVAL_245 = _EVAL_145 & _EVAL_506;
  assign icache__EVAL_22 = _EVAL_83;
  assign _EVAL_401 = _EVAL_529 | _EVAL_309;
  assign _EVAL_462 = _EVAL_202 & _EVAL_255;
  assign _EVAL_62 = icache__EVAL_14;
  assign tlb__EVAL_7 = _EVAL_79;
  assign _EVAL_504 = _EVAL_327[14];
  assign _EVAL_425 = {_EVAL_570, 1'h0};
  assign icache__EVAL_26 = _EVAL_72;
  assign _EVAL_254 = _EVAL_222[24:21];
  assign _EVAL_362 = _EVAL_390[7];
  assign _EVAL_361 = _EVAL_250 & _EVAL_322;
  assign btb__EVAL_13 = _EVAL_128[31:0];
  assign _EVAL_266 = _EVAL_406 == 5'h0;
  assign fq__EVAL = _EVAL_403[1:0];
  assign _EVAL_354 = _EVAL_330;
  assign _EVAL_332 = _EVAL_453 ? _EVAL_214 : _EVAL_154;
  assign _EVAL_68 = fq__EVAL_14;
  assign _EVAL_486 = _EVAL_129 & _EVAL_233;
  assign _EVAL_133 = _EVAL_188 ? 5'h1c : _EVAL_563;
  assign btb__EVAL_1 = _EVAL_298 ? 1'h0 : _EVAL_64;
  assign _EVAL_324 = _EVAL_453 ? _EVAL_510 : {{1'd0}, _EVAL_515};
  assign _EVAL_472 = _EVAL_136 | _EVAL_452;
  assign btb__EVAL_15 = _EVAL_301 ? _EVAL_522 : _EVAL_23;
  assign _EVAL_348 = _EVAL_404 & _EVAL_266;
  assign tlb__EVAL_60 = _EVAL_4;
  assign _EVAL_284 = _EVAL_345 | _EVAL_303;
  assign _EVAL_488 = ~_EVAL_229;
  assign tlb__EVAL_16 = _EVAL_1;
  assign _EVAL_166 = _EVAL_356 & _EVAL_542;
  assign _EVAL_300 = _EVAL_570 ? _EVAL_434 : _EVAL_192;
  assign _EVAL_190 = _EVAL_222[19:15];
  assign tlb__EVAL_47 = _EVAL_71;
  assign _EVAL_207 = _EVAL_421 & _EVAL_561;
  assign _EVAL_19 = 1'h0;
  assign _EVAL_475 = _EVAL_335;
  assign btb__EVAL_7 = _EVAL_570 ? _EVAL_122 : _EVAL_240;
  assign _EVAL_449 = _EVAL_522 | _EVAL_236;
  assign _EVAL_131 = ~_EVAL_346;
  assign _EVAL_215 = ~_EVAL_178;
  assign _EVAL_288 = _EVAL_269 & _EVAL_232;
  assign _EVAL_423 = {_EVAL_461,_EVAL_280,_EVAL_198,_EVAL_147,_EVAL_220,_EVAL_254,1'h0};
  assign _EVAL_176 = _EVAL_162 & _EVAL_219;
  assign _EVAL_436 = {{1{_EVAL_473[31]}},_EVAL_473};
  assign _EVAL_506 = ~_EVAL_278;
  assign _EVAL_408 = _EVAL_371[31:0];
  assign _EVAL_399 = icache__EVAL_13 & _EVAL_155;
  assign _EVAL_202 = _EVAL_129 & _EVAL_506;
  assign _EVAL_296 = _EVAL_327[4:3];
  assign _EVAL_228 = 16'h9002 == _EVAL_191;
  assign _EVAL_278 = _EVAL_394 != 2'h3;
  assign _EVAL_421 = _EVAL_432 & _EVAL_323;
  assign _EVAL_537 = _EVAL_18 | _EVAL_189;
  assign _EVAL_365 = _EVAL_327[7];
  assign _EVAL_386 = {11{_EVAL_475}};
  assign _EVAL_268 = ~_EVAL_567;
  assign _EVAL_144 = _EVAL_327[11];
  assign _EVAL_524 = ~_EVAL_177;
  assign _EVAL_73 = fq__EVAL_16;
  assign _EVAL_467 = _EVAL_181 | _EVAL_289;
  assign btb__EVAL_5 = gated_clock_icache_clock_gate_out;
  assign _EVAL_204 = _EVAL_459 ? 2'h2 : {{1'd0}, _EVAL_376};
  assign _EVAL_121 = _EVAL_423;
  assign btb__EVAL_4 = _EVAL_301 ? _EVAL_441 : _EVAL_65;
  assign _EVAL_327 = fq__EVAL_18[15:0];
  assign _EVAL_309 = _EVAL_400 & _EVAL_432;
  assign _EVAL_230 = _EVAL_439 & _EVAL_432;
  assign _EVAL_282 = ~_EVAL_187;
  assign _EVAL_494 = _EVAL_202 ? _EVAL_439 : _EVAL_184;
  assign _EVAL_416 = {11{_EVAL_126}};
  assign _EVAL_188 = _EVAL_516 | _EVAL_525;
  assign _EVAL_239 = _EVAL_163[32:0];
  assign _EVAL_439 = _EVAL_311 == 7'h63;
  assign _EVAL_242 = _EVAL_495 ? _EVAL_485 : _EVAL_167;
  assign _EVAL_345 = _EVAL_202 & _EVAL_289;
  assign _EVAL_185 = _EVAL_383 | _EVAL_340;
  assign _EVAL_446 = _EVAL_239;
  assign _EVAL_315 = _EVAL_555 & _EVAL_445;
  assign _EVAL_192 = _EVAL_453 & _EVAL_123;
  assign _EVAL_541 = _EVAL_378 & _EVAL_468;
  assign _EVAL_501 = _EVAL_453 ? _EVAL_514 : _EVAL_324;
  assign _EVAL_267 = _EVAL_205 & 5'h1b;
  assign _EVAL_47 = icache__EVAL_3;
  assign _EVAL_301 = ~_EVAL_65;
  assign icache__EVAL_18 = _EVAL;
  assign tlb__EVAL_49 = _EVAL_108;
  assign _EVAL_428 = _EVAL_382 | _EVAL_188;
  assign _EVAL_381 = _EVAL_398 & _EVAL_527;
  assign _EVAL_522 = ~_EVAL_320;
  assign _EVAL_470 = _EVAL_241 | _EVAL_555;
  assign icache__EVAL_28 = _EVAL_8;
  assign _EVAL_392 = 16'ha001 == _EVAL_248;
  assign _EVAL_206 = ~_EVAL_275;
  assign _EVAL_148 = _EVAL_307 ? 10'h3ff : 10'h0;
  assign _EVAL_199 = _EVAL_186 | _EVAL_375;
  assign icache__EVAL_17 = gated_clock_icache_clock_gate_out;
  assign tlb__EVAL_33 = _EVAL_117;
  assign _EVAL_112 = fq__EVAL_17;
  assign _EVAL_336 = _EVAL_245 | _EVAL_25;
  assign _EVAL_128 = _EVAL_522 + _EVAL_225;
  assign _EVAL_453 = ~_EVAL_382;
  assign _EVAL_394 = _EVAL_327[1:0];
  assign _EVAL_375 = _EVAL_288 & _EVAL_184;
  assign tlb__EVAL_54 = _EVAL_22;
  assign _EVAL_174 = _EVAL_202 ? _EVAL_408 : _EVAL_503;
  assign _EVAL_10 = fq__EVAL_20;
  assign tlb__EVAL_5 = _EVAL_120;
  assign _EVAL_406 = _EVAL_390[6:2];
  assign _EVAL_352 = _EVAL_373;
  assign _EVAL_418 = _EVAL_421 | _EVAL_517;
  assign _EVAL_286 = 5'h1 == _EVAL_201;
  assign _EVAL_380 = _EVAL_495 & _EVAL_485;
  assign fq__EVAL_4 = _EVAL_453 ? _EVAL_431 : _EVAL_567;
  assign _EVAL_411 = _EVAL_331 | _EVAL_18;
  assign _EVAL_150 = 5'h1 == _EVAL_227;
  assign _EVAL_490 = _EVAL_290 ? 10'h3ff : 10'h0;
  assign tlb__EVAL_28 = _EVAL_50;
  assign icache__EVAL_13 = _EVAL_560 | _EVAL_552;
  assign _EVAL_303 = _EVAL_288 & _EVAL_353;
  assign _EVAL_483 = ~_EVAL_543;
  assign _EVAL_292 = _EVAL_185 | _EVAL_361;
  assign _EVAL_371 = _EVAL_503 - 32'h2;
  assign _EVAL_319 = _EVAL_162 | _EVAL_219;
  assign _EVAL_103 = _EVAL_159[31:0];
  assign _EVAL_285 = _EVAL_538 & _EVAL_397;
  assign _EVAL_187 = fq__EVAL_10[1];
  assign tlb__EVAL_11 = _EVAL_53;
  assign _EVAL_269 = fq__EVAL[1];
  assign _EVAL_466 = _EVAL_363[24:21];
  assign _EVAL_182 = _EVAL_169;
  assign _EVAL_480 = _EVAL_427 + 32'h4;
  assign fq__EVAL_3 = _EVAL_433 | _EVAL_552;
  assign _EVAL_186 = _EVAL_202 & _EVAL_439;
  assign tlb__EVAL_13 = _EVAL_59;
  assign _EVAL_167 = _EVAL_291 & _EVAL_150;
  assign btb__EVAL_17 = _EVAL_54;
  assign tlb__EVAL_34 = _EVAL_21;
  assign _EVAL_243 = _EVAL_313 & 5'h1b;
  assign _EVAL_508 = _EVAL_536 ? $signed({{8{_EVAL_443[12]}},_EVAL_443}) : $signed(_EVAL_352);
  assign icache__EVAL_36 = _EVAL_557;
  assign _EVAL_477 = 16'he001 == _EVAL_248;
  assign _EVAL_161 = ~_EVAL_200;
  assign gated_clock_icache_clock_gate_en = _EVAL_218 | _EVAL_104;
  assign _EVAL_397 = ~_EVAL_284;
  assign _EVAL_473 = _EVAL_522;
  assign icache__EVAL_30 = tlb__EVAL_2;
  assign _EVAL_382 = _EVAL_556 & _EVAL_565;
  assign _EVAL_525 = _EVAL_462 | _EVAL_274;
  assign _EVAL_434 = _EVAL_453 ? _EVAL_450 : _EVAL_192;
  assign _EVAL_460 = _EVAL_152;
  assign fq__EVAL_13 = _EVAL_273 | _EVAL_158;
  assign _EVAL_383 = 16'ha001 == _EVAL_308;
  assign _EVAL_500 = {8{_EVAL_126}};
  assign _EVAL_209 = _EVAL_524 & _EVAL_176;
  assign _EVAL_402 = _EVAL_480[31:0];
  assign _EVAL_183 = _EVAL_570 ? _EVAL_212 : _EVAL_511;
  assign _EVAL_305 = _EVAL_467 & _EVAL_200;
  assign _EVAL_450 = _EVAL_413 | _EVAL_192;
  assign _EVAL_388 = _EVAL_331 & _EVAL_428;
  assign _EVAL_236 = {{30'd0}, _EVAL_425};
  assign btb__EVAL_24 = _EVAL_301 ? 5'h1c : _EVAL_43;
  assign _EVAL_549 = _EVAL_129 & _EVAL_167;
  assign _EVAL_168 = _EVAL_253 | _EVAL_348;
  assign _EVAL_217 = _EVAL_124;
  assign _EVAL_293 = _EVAL_533 & _EVAL_281;
  assign _EVAL_6 = _EVAL_66 & _EVAL_19;
  assign fq__EVAL_5 = _EVAL_507 & _EVAL_546;
  assign _EVAL_323 = _EVAL_127 | _EVAL_486;
  assign _EVAL_208 = _EVAL_390[2];
  assign icache__EVAL_7 = _EVAL_51;
  assign _EVAL_162 = ~_EVAL_564;
  assign _EVAL_513 = _EVAL_222[19:12];
  assign tlb__EVAL_21 = _EVAL_96;
  assign _EVAL_568 = _EVAL_270 ? $signed(_EVAL_121) : $signed(_EVAL_156);
  assign _EVAL_302 = _EVAL_354;
  assign _EVAL_283 = _EVAL_390[11];
  assign _EVAL_140 = _EVAL_340 | _EVAL_361;
  assign icache__EVAL_5 = _EVAL_18 | _EVAL_189;
  assign _EVAL_357 = ~_EVAL_495;
  assign icache__EVAL_33 = _EVAL_92;
  assign _EVAL_240 = _EVAL_242 ? 2'h3 : _EVAL_204;
  assign _EVAL_172 = _EVAL_202 ? $signed(_EVAL_502) : $signed({{11{_EVAL_508[20]}},_EVAL_508});
  assign _EVAL_430 = _EVAL_327[11:10];
  assign _EVAL_101 = icache__EVAL_6;
  assign tlb__EVAL_35 = _EVAL_38;
  assign _EVAL_274 = _EVAL_288 & _EVAL_143;
  assign _EVAL_178 = btb__EVAL_19 & _EVAL_146;
  assign _EVAL_260 = ~_EVAL_560;
  assign _EVAL_476 = _EVAL_504 ? $signed({{8{_EVAL_265[12]}},_EVAL_265}) : $signed(_EVAL_217);
  assign _EVAL_339 = _EVAL_447 & _EVAL_497;
  assign icache__EVAL_31 = _EVAL_74;
  assign _EVAL_142 = _EVAL_188 ? _EVAL_411 : _EVAL_18;
  assign _EVAL_443 = _EVAL_498;
  assign gated_clock_icache_clock_gate_test_en = _EVAL_70;
  assign _EVAL_129 = _EVAL_368 & _EVAL_357;
  assign tlb__EVAL_40 = _EVAL_60;
  assign _EVAL_414 = _EVAL_575;
  assign _EVAL_461 = _EVAL_475;
  assign _EVAL_417 = ~_EVAL_552;
  assign tlb__EVAL = _EVAL_41;
  assign fq__EVAL_15 = _EVAL_453 ? _EVAL_261 : _EVAL_382;
  assign _EVAL_487 = _EVAL_570 ? _EVAL_501 : _EVAL_324;
  assign tlb__EVAL_36 = _EVAL_90;
  assign _EVAL_130 = _EVAL_555 & _EVAL_418;
  assign _EVAL_146 = _EVAL_380 | _EVAL_549;
  assign tlb__EVAL_9 = _EVAL_57;
  assign _EVAL_330 = _EVAL_363[19:12];
  assign _EVAL_139 = _EVAL_262 != 2'h3;
  assign fq__EVAL_19 = _EVAL_45;
  assign _EVAL_347 = _EVAL_202 ? _EVAL_541 : _EVAL_474;
  assign _EVAL_516 = _EVAL_545 | _EVAL_350;
  assign _EVAL_499 = _EVAL_305 | _EVAL_541;
  assign _EVAL_505 = _EVAL_327[6:5];
  always @(posedge _EVAL_100) begin
    _EVAL_218 <= _EVAL_470 | _EVAL_524;
  end
  always @(posedge gated_clock_icache_clock_gate_out) begin
    _EVAL_550 <= _EVAL_77 | _EVAL_272;
    _EVAL_551 <= _EVAL_564;
    if (_EVAL_533) begin
      _EVAL_552 <= tlb__EVAL_12;
    end
    if (_EVAL_77) begin
      _EVAL_553 <= 1'h0;
    end else if (_EVAL_18) begin
      _EVAL_553 <= 1'h0;
    end else if (_EVAL_570) begin
      if (_EVAL_453) begin
        _EVAL_553 <= _EVAL_175;
      end else begin
        _EVAL_553 <= _EVAL_367;
      end
    end else begin
      _EVAL_553 <= _EVAL_367;
    end
    if (_EVAL_331) begin
      if (_EVAL_379) begin
        _EVAL_554 <= _EVAL_170;
      end
    end
    if (_EVAL_77) begin
      _EVAL_555 <= 1'h0;
    end else begin
      _EVAL_555 <= _EVAL_293;
    end
    if (_EVAL_533) begin
      _EVAL_556 <= btb__EVAL_2;
    end
    if (_EVAL_77) begin
      _EVAL_557 <= _EVAL_344;
    end else if (_EVAL_533) begin
      _EVAL_557 <= _EVAL_558;
    end
    _EVAL_558 <= _EVAL_103;
    if (_EVAL_533) begin
      _EVAL_559 <= btb__EVAL_16;
    end
    if (_EVAL_77) begin
      _EVAL_560 <= 1'h0;
    end else if (_EVAL_533) begin
      _EVAL_560 <= _EVAL_566;
    end
    if (_EVAL_533) begin
      _EVAL_561 <= btb__EVAL_23;
    end
    if (_EVAL_77) begin
      _EVAL_562 <= 1'h0;
    end else if (_EVAL_464) begin
      _EVAL_562 <= 1'h0;
    end else if (_EVAL_388) begin
      _EVAL_562 <= 1'h0;
    end else if (_EVAL_331) begin
      _EVAL_562 <= _EVAL_379;
    end
    if (_EVAL_533) begin
      _EVAL_563 <= btb__EVAL_18;
    end
    _EVAL_564 <= _EVAL_18 | _EVAL_189;
    if (_EVAL_533) begin
      _EVAL_565 <= btb__EVAL_22;
    end
    if (_EVAL_18) begin
      _EVAL_566 <= _EVAL_118;
    end else if (_EVAL_276) begin
      _EVAL_566 <= _EVAL_560;
    end else begin
      _EVAL_566 <= _EVAL_138;
    end
    if (_EVAL_533) begin
      _EVAL_567 <= btb__EVAL_28;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_218 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_550 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_551 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_552 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_553 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_554 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_555 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_556 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_557 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_558 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_559 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_560 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_561 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_562 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_563 = _RAND_14[4:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_564 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_565 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _EVAL_566 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _EVAL_567 = _RAND_18[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
