//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_143(
  input   _EVAL,
  input   _EVAL_0,
  output  _EVAL_1
);
  wire  output_chain__EVAL;
  wire  output_chain__EVAL_0;
  wire  output_chain__EVAL_1;
  _EVAL_142 output_chain (
    ._EVAL(output_chain__EVAL),
    ._EVAL_0(output_chain__EVAL_0),
    ._EVAL_1(output_chain__EVAL_1)
  );
  assign output_chain__EVAL_0 = _EVAL_0;
  assign output_chain__EVAL_1 = _EVAL;
  assign _EVAL_1 = output_chain__EVAL;
endmodule
