//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_90_assert(
  input  [2:0]  _EVAL,
  input  [2:0]  _EVAL_0,
  input         _EVAL_1,
  input  [4:0]  _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [3:0]  _EVAL_9,
  input  [4:0]  _EVAL_10,
  input  [2:0]  _EVAL_11,
  input         _EVAL_12,
  input  [14:0] _EVAL_13,
  input  [2:0]  _EVAL_14
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_15;
  reg [4:0] _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire [3:0] _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire [1:0] _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire [31:0] _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire [3:0] _EVAL_46;
  wire  _EVAL_47;
  reg [14:0] _EVAL_48;
  wire  _EVAL_49;
  wire [31:0] _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire [2:0] _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire [1:0] _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire [5:0] _EVAL_74;
  reg [3:0] _EVAL_75;
  wire  _EVAL_76;
  wire [12:0] _EVAL_77;
  wire [12:0] _EVAL_78;
  wire  _EVAL_79;
  reg [3:0] _EVAL_80;
  wire [17:0] _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  reg [2:0] _EVAL_89;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire [17:0] _EVAL_96;
  wire  _EVAL_97;
  reg [3:0] _EVAL_98;
  wire [17:0] _EVAL_99;
  wire  _EVAL_100;
  wire [3:0] _EVAL_101;
  wire  _EVAL_102;
  wire [15:0] _EVAL_103;
  wire  _EVAL_104;
  wire [3:0] _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire [14:0] _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire [15:0] _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire [31:0] _EVAL_138;
  wire  _EVAL_139;
  wire [14:0] _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire [1:0] _EVAL_143;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire [31:0] _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire [17:0] _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  reg [3:0] _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire [5:0] _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire [31:0] _EVAL_174;
  wire [4:0] _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  reg [2:0] _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire [17:0] _EVAL_184;
  wire [4:0] _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire [15:0] _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire [17:0] _EVAL_198;
  wire [2:0] _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire [4:0] _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_207;
  wire [3:0] _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  reg [17:0] _EVAL_222;
  reg [2:0] _EVAL_223;
  wire [5:0] _EVAL_224;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire [5:0] _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire [3:0] _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire [14:0] _EVAL_238;
  wire [3:0] _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire [3:0] _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire [17:0] _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_256;
  wire [17:0] _EVAL_257;
  wire [1:0] _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire [4:0] _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  reg [4:0] _EVAL_264;
  wire  _EVAL_265;
  wire [3:0] _EVAL_266;
  reg [2:0] _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  reg [31:0] _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  reg [2:0] _EVAL_276;
  wire [32:0] _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire [3:0] _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_266 = _EVAL_9 & _EVAL_101;
  assign _EVAL_218 = _EVAL_69 & _EVAL_232;
  assign _EVAL_279 = ~_EVAL_62;
  assign _EVAL_137 = _EVAL_5 == 3'h0;
  assign _EVAL_221 = _EVAL == 3'h4;
  assign _EVAL_101 = ~_EVAL_239;
  assign _EVAL_177 = _EVAL_229 & _EVAL_62;
  assign _EVAL_167 = _EVAL_59 | _EVAL_183;
  assign _EVAL_242 = ~_EVAL_51;
  assign _EVAL_217 = _EVAL_151 & _EVAL_201;
  assign _EVAL_269 = _EVAL_3 & _EVAL_221;
  assign _EVAL_92 = _EVAL_7 & _EVAL_17;
  assign _EVAL_41 = _EVAL_3 & _EVAL_79;
  assign _EVAL_39 = _EVAL_14 == 3'h2;
  assign _EVAL_278 = _EVAL_273 | _EVAL_8;
  assign _EVAL_226 = _EVAL_10 == 5'h8;
  assign _EVAL_61 = 3'h6 == _EVAL_11;
  assign _EVAL_115 = _EVAL_131 | _EVAL_8;
  assign _EVAL_248 = _EVAL_37 | _EVAL_8;
  assign _EVAL_155 = ~_EVAL_259;
  assign _EVAL_273 = _EVAL_5 <= 3'h2;
  assign _EVAL_204 = _EVAL_102 | _EVAL_216;
  assign _EVAL_212 = _EVAL_7 & _EVAL_113;
  assign _EVAL_196 = ~_EVAL_100;
  assign _EVAL_25 = _EVAL_10[4:3];
  assign _EVAL_169 = _EVAL_3 & _EVAL_147;
  assign _EVAL_197 = _EVAL_32 & _EVAL_282;
  assign _EVAL_246 = _EVAL_14 == 3'h0;
  assign _EVAL_235 = ~_EVAL_281;
  assign _EVAL_262 = _EVAL_132 | _EVAL_146;
  assign _EVAL_108 = _EVAL == 3'h1;
  assign _EVAL_270 = _EVAL_11 == _EVAL_89;
  assign _EVAL_147 = _EVAL == 3'h6;
  assign _EVAL_113 = _EVAL_14 == 3'h3;
  assign _EVAL_208 = _EVAL_185[3:0];
  assign _EVAL_40 = ~_EVAL_8;
  assign _EVAL_257 = _EVAL_138[17:0];
  assign _EVAL_28 = _EVAL_2 == _EVAL_16;
  assign _EVAL_176 = _EVAL_53 | _EVAL_8;
  assign _EVAL_82 = _EVAL_262 | _EVAL_265;
  assign _EVAL_72 = _EVAL_119 & _EVAL_229;
  assign _EVAL_172 = _EVAL_266 == 4'h0;
  assign _EVAL_96 = ~_EVAL_257;
  assign _EVAL_20 = _EVAL_14[2];
  assign _EVAL_253 = _EVAL_153[17:0];
  assign _EVAL_117 = _EVAL_14 == _EVAL_276;
  assign _EVAL_27 = _EVAL_3 & _EVAL_236;
  assign _EVAL_146 = _EVAL_2 == 5'h10;
  assign _EVAL_34 = _EVAL_190 & _EVAL_279;
  assign _EVAL_240 = _EVAL_143 == 2'h0;
  assign _EVAL_111 = _EVAL_5 == _EVAL_268;
  assign _EVAL_64 = _EVAL_142 | _EVAL_8;
  assign _EVAL_280 = _EVAL_261[3:0];
  assign _EVAL_43 = _EVAL_172 | _EVAL_8;
  assign _EVAL_17 = _EVAL_14 == 3'h7;
  assign _EVAL_112 = $signed(_EVAL_103) & -16'sh1000;
  assign _EVAL_156 = _EVAL_14 == 3'h1;
  assign _EVAL_120 = _EVAL_19 | _EVAL_8;
  assign _EVAL_31 = _EVAL_69 & _EVAL_84;
  assign _EVAL_200 = _EVAL_157 | _EVAL_226;
  assign _EVAL_160 = _EVAL_173 | _EVAL_125;
  assign _EVAL_165 = _EVAL_204 | _EVAL_249;
  assign _EVAL_136 = ~_EVAL_115;
  assign _EVAL_95 = ~_EVAL_29;
  assign _EVAL_237 = _EVAL_104 | _EVAL_69;
  assign _EVAL_281 = _EVAL_68 | _EVAL_8;
  assign _EVAL_129 = ~_EVAL_73;
  assign _EVAL_103 = {1'b0,$signed(_EVAL_109)};
  assign _EVAL_219 = |_EVAL_222;
  assign _EVAL_265 = _EVAL_61 & _EVAL_149;
  assign _EVAL_245 = _EVAL_7 & _EVAL_39;
  assign _EVAL_85 = ~_EVAL_83;
  assign _EVAL_105 = _EVAL_203[3:0];
  assign _EVAL_106 = _EVAL_7 & _EVAL_207;
  assign _EVAL_164 = _EVAL_11 <= 3'h2;
  assign _EVAL_193 = _EVAL_31 & _EVAL_195;
  assign _EVAL_59 = _EVAL_253 != _EVAL_257;
  assign _EVAL_37 = _EVAL_0 == _EVAL_181;
  assign _EVAL_236 = _EVAL == 3'h5;
  assign _EVAL_189 = ~_EVAL_260;
  assign _EVAL_109 = _EVAL_13 ^ 15'h4000;
  assign _EVAL_241 = ~_EVAL_141;
  assign _EVAL_45 = _EVAL_117 | _EVAL_8;
  assign _EVAL_252 = _EVAL_200 | _EVAL_8;
  assign _EVAL_35 = ~_EVAL_278;
  assign _EVAL_127 = ~_EVAL_247;
  assign _EVAL_33 = _EVAL_204 | _EVAL_170;
  assign _EVAL_66 = _EVAL_194 | _EVAL_8;
  assign _EVAL_124 = _EVAL_271 | _EVAL_8;
  assign _EVAL_38 = _EVAL_238 == 15'h0;
  assign _EVAL_277 = _EVAL_272 + 32'h1;
  assign _EVAL_233 = |_EVAL_253;
  assign _EVAL_15 = _EVAL_145 | _EVAL_8;
  assign _EVAL_130 = _EVAL_14 == 3'h4;
  assign _EVAL_53 = _EVAL_9 == _EVAL_239;
  assign _EVAL_227 = ~_EVAL_248;
  assign _EVAL_224 = _EVAL_77[5:0];
  assign _EVAL_214 = ~_EVAL_18;
  assign _EVAL_71 = _EVAL_123 | _EVAL_8;
  assign _EVAL_201 = _EVAL_229 & _EVAL_279;
  assign _EVAL_44 = ~_EVAL_47;
  assign _EVAL_122 = _EVAL_7 & _EVAL_256;
  assign _EVAL_134 = _EVAL_5 <= 3'h4;
  assign _EVAL_234 = _EVAL_175[3:0];
  assign _EVAL_104 = _EVAL_12 & _EVAL_7;
  assign _EVAL_74 = _EVAL_78[5:0];
  assign _EVAL_260 = _EVAL_134 | _EVAL_8;
  assign _EVAL_140 = {{9'd0}, _EVAL_230};
  assign _EVAL_65 = 2'h1 << _EVAL_283;
  assign _EVAL_52 = _EVAL_7 & _EVAL_130;
  assign _EVAL_220 = _EVAL_187 | _EVAL_210;
  assign _EVAL_249 = _EVAL_151 & _EVAL_231;
  assign _EVAL_211 = _EVAL_57 <= 3'h6;
  assign _EVAL_42 = ~_EVAL_66;
  assign _EVAL_231 = _EVAL_190 & _EVAL_62;
  assign _EVAL_174 = 32'h1 << _EVAL_10;
  assign _EVAL_282 = $signed(_EVAL_188) == 16'sh0;
  assign _EVAL_173 = ~_EVAL_219;
  assign _EVAL_145 = _EVAL_0 >= 3'h2;
  assign _EVAL_76 = ~_EVAL_20;
  assign _EVAL_49 = _EVAL_272 < plusarg_reader_out;
  assign _EVAL_141 = _EVAL_167 | _EVAL_8;
  assign _EVAL_154 = _EVAL_178 | _EVAL_110;
  assign _EVAL_203 = _EVAL_80 - 4'h1;
  assign _EVAL_157 = _EVAL_154 | _EVAL_274;
  assign _EVAL_209 = _EVAL_244 | _EVAL_8;
  assign _EVAL_191 = _EVAL_187 | _EVAL_146;
  assign _EVAL_151 = _EVAL_258[0];
  assign _EVAL_163 = ~_EVAL_124;
  assign _EVAL_283 = _EVAL_11[0];
  assign _EVAL_47 = _EVAL_81[0];
  assign _EVAL_247 = _EVAL_197 | _EVAL_8;
  assign _EVAL_271 = _EVAL_5 <= 3'h3;
  assign _EVAL_195 = ~_EVAL_147;
  assign _EVAL_202 = _EVAL_3 & _EVAL_108;
  assign _EVAL_118 = ~_EVAL_232;
  assign _EVAL_68 = ~_EVAL_4;
  assign _EVAL_69 = _EVAL_6 & _EVAL_3;
  assign _EVAL_54 = _EVAL_10 == _EVAL_264;
  assign _EVAL_216 = _EVAL_119 & _EVAL_190;
  assign _EVAL_210 = _EVAL_240 & _EVAL_215;
  assign _EVAL_84 = _EVAL_80 == 4'h0;
  assign _EVAL_152 = _EVAL_7 & _EVAL_156;
  assign _EVAL_30 = _EVAL_270 | _EVAL_8;
  assign _EVAL_244 = _EVAL_13 == _EVAL_48;
  assign _EVAL_190 = ~_EVAL_229;
  assign _EVAL_261 = _EVAL_75 - 4'h1;
  assign _EVAL_36 = _EVAL_277[31:0];
  assign _EVAL_131 = _EVAL == _EVAL_223;
  assign _EVAL_81 = _EVAL_222 >> _EVAL_2;
  assign _EVAL_274 = _EVAL_60 & _EVAL_211;
  assign _EVAL_99 = _EVAL_198 >> _EVAL_10;
  assign _EVAL_24 = ~_EVAL_176;
  assign _EVAL_251 = ~_EVAL_64;
  assign _EVAL_179 = ~_EVAL_15;
  assign _EVAL_78 = 13'h3f << _EVAL_0;
  assign _EVAL_77 = 13'h3f << _EVAL_11;
  assign _EVAL_132 = _EVAL_164 & _EVAL_220;
  assign _EVAL_79 = _EVAL == 3'h2;
  assign _EVAL_123 = _EVAL_160 | _EVAL_49;
  assign _EVAL_254 = ~_EVAL_252;
  assign _EVAL_175 = _EVAL_162 - 4'h1;
  assign _EVAL_178 = _EVAL_10 == 5'h11;
  assign _EVAL_138 = _EVAL_193 ? _EVAL_174 : 32'h0;
  assign _EVAL_205 = _EVAL == 3'h0;
  assign _EVAL_238 = _EVAL_13 & _EVAL_140;
  assign _EVAL_70 = ~_EVAL_87;
  assign _EVAL_62 = _EVAL_13[0];
  assign _EVAL_168 = ~_EVAL_74;
  assign _EVAL_186 = _EVAL[0];
  assign _EVAL_207 = _EVAL_14 == 3'h6;
  assign _EVAL_187 = _EVAL_2 == 5'h11;
  assign _EVAL_86 = ~_EVAL_71;
  assign _EVAL_263 = ~_EVAL_192;
  assign _EVAL_182 = ~_EVAL_58;
  assign _EVAL_83 = _EVAL_44 | _EVAL_8;
  assign _EVAL_243 = ~_EVAL_9;
  assign _EVAL_159 = ~_EVAL_30;
  assign _EVAL_139 = _EVAL_171 | _EVAL_8;
  assign _EVAL_215 = _EVAL_199 <= 3'h6;
  assign _EVAL_198 = _EVAL_253 | _EVAL_222;
  assign _EVAL_88 = ~_EVAL_43;
  assign _EVAL_100 = _EVAL_28 | _EVAL_8;
  assign _EVAL_142 = _EVAL_243 == 4'h0;
  assign _EVAL_258 = _EVAL_65 | 2'h1;
  assign _EVAL_171 = _EVAL_99[0];
  assign _EVAL_116 = _EVAL_191 | _EVAL_210;
  assign _EVAL_22 = ~_EVAL_120;
  assign _EVAL_183 = ~_EVAL_233;
  assign _EVAL_239 = {_EVAL_180,_EVAL_161,_EVAL_165,_EVAL_33};
  assign _EVAL_58 = _EVAL_111 | _EVAL_8;
  assign _EVAL_50 = 32'h1 << _EVAL_2;
  assign _EVAL_184 = _EVAL_222 | _EVAL_253;
  assign _EVAL_150 = ~_EVAL_97;
  assign _EVAL_97 = _EVAL_38 | _EVAL_8;
  assign _EVAL_229 = _EVAL_13[1];
  assign _EVAL_166 = _EVAL_3 & _EVAL_118;
  assign _EVAL_153 = _EVAL_23 ? _EVAL_50 : 32'h0;
  assign _EVAL_192 = _EVAL_82 | _EVAL_8;
  assign _EVAL_55 = _EVAL_128 | _EVAL_8;
  assign _EVAL_57 = _EVAL_10[2:0];
  assign _EVAL_94 = ~_EVAL_209;
  assign _EVAL_91 = _EVAL_102 | _EVAL_72;
  assign _EVAL_232 = _EVAL_75 == 4'h0;
  assign _EVAL_29 = _EVAL_162 == 4'h0;
  assign _EVAL_23 = _EVAL_104 & _EVAL_67;
  assign _EVAL_180 = _EVAL_91 | _EVAL_26;
  assign _EVAL_125 = plusarg_reader_out == 32'h0;
  assign _EVAL_114 = _EVAL_3 & _EVAL_205;
  assign _EVAL_275 = ~_EVAL_45;
  assign _EVAL_185 = _EVAL_98 - 4'h1;
  assign _EVAL_126 = _EVAL_104 & _EVAL_29;
  assign _EVAL_135 = _EVAL_5 <= 3'h1;
  assign _EVAL_67 = _EVAL_98 == 4'h0;
  assign _EVAL_259 = _EVAL_137 | _EVAL_8;
  assign _EVAL_60 = _EVAL_25 == 2'h0;
  assign _EVAL_21 = _EVAL_168[5:2];
  assign _EVAL_128 = _EVAL_116 | _EVAL_149;
  assign _EVAL_110 = _EVAL_10 == 5'h10;
  assign _EVAL_161 = _EVAL_91 | _EVAL_217;
  assign _EVAL_46 = _EVAL_230[5:2];
  assign _EVAL_170 = _EVAL_151 & _EVAL_34;
  assign _EVAL_19 = _EVAL_262 & _EVAL_197;
  assign _EVAL_119 = _EVAL_258[1];
  assign _EVAL_194 = _EVAL <= 3'h6;
  assign _EVAL_87 = _EVAL_228 | _EVAL_8;
  assign _EVAL_143 = _EVAL_2[4:3];
  assign _EVAL_199 = _EVAL_2[2:0];
  assign _EVAL_73 = _EVAL_54 | _EVAL_8;
  assign _EVAL_148 = ~_EVAL_139;
  assign _EVAL_133 = _EVAL_7 & _EVAL_246;
  assign _EVAL_158 = _EVAL_184 & _EVAL_96;
  assign _EVAL_188 = _EVAL_112;
  assign _EVAL_26 = _EVAL_151 & _EVAL_177;
  assign _EVAL_230 = ~_EVAL_224;
  assign _EVAL_149 = _EVAL_2 == 5'h8;
  assign _EVAL_32 = _EVAL_11 <= 3'h6;
  assign _EVAL_18 = _EVAL_135 | _EVAL_8;
  assign _EVAL_63 = _EVAL_7 & _EVAL_95;
  assign _EVAL_102 = _EVAL_11 >= 3'h2;
  assign _EVAL_107 = ~_EVAL_55;
  assign _EVAL_51 = _EVAL_102 | _EVAL_8;
  assign _EVAL_256 = _EVAL_14 == 3'h5;
  assign _EVAL_228 = _EVAL_5 != 3'h0;
  always @(posedge _EVAL_1) begin
    if (_EVAL_126) begin
      _EVAL_16 <= _EVAL_2;
    end
    if (_EVAL_126) begin
      _EVAL_48 <= _EVAL_13;
    end
    if (_EVAL_8) begin
      _EVAL_75 <= 4'h0;
    end else if (_EVAL_69) begin
      if (_EVAL_232) begin
        if (_EVAL_186) begin
          _EVAL_75 <= _EVAL_21;
        end else begin
          _EVAL_75 <= 4'h0;
        end
      end else begin
        _EVAL_75 <= _EVAL_280;
      end
    end
    if (_EVAL_8) begin
      _EVAL_80 <= 4'h0;
    end else if (_EVAL_69) begin
      if (_EVAL_84) begin
        if (_EVAL_186) begin
          _EVAL_80 <= _EVAL_21;
        end else begin
          _EVAL_80 <= 4'h0;
        end
      end else begin
        _EVAL_80 <= _EVAL_105;
      end
    end
    if (_EVAL_126) begin
      _EVAL_89 <= _EVAL_11;
    end
    if (_EVAL_8) begin
      _EVAL_98 <= 4'h0;
    end else if (_EVAL_104) begin
      if (_EVAL_67) begin
        if (_EVAL_76) begin
          _EVAL_98 <= _EVAL_46;
        end else begin
          _EVAL_98 <= 4'h0;
        end
      end else begin
        _EVAL_98 <= _EVAL_208;
      end
    end
    if (_EVAL_8) begin
      _EVAL_162 <= 4'h0;
    end else if (_EVAL_104) begin
      if (_EVAL_29) begin
        if (_EVAL_76) begin
          _EVAL_162 <= _EVAL_46;
        end else begin
          _EVAL_162 <= 4'h0;
        end
      end else begin
        _EVAL_162 <= _EVAL_234;
      end
    end
    if (_EVAL_218) begin
      _EVAL_181 <= _EVAL_0;
    end
    if (_EVAL_8) begin
      _EVAL_222 <= 18'h0;
    end else begin
      _EVAL_222 <= _EVAL_158;
    end
    if (_EVAL_218) begin
      _EVAL_223 <= _EVAL;
    end
    if (_EVAL_218) begin
      _EVAL_264 <= _EVAL_10;
    end
    if (_EVAL_126) begin
      _EVAL_268 <= _EVAL_5;
    end
    if (_EVAL_8) begin
      _EVAL_272 <= 32'h0;
    end else if (_EVAL_237) begin
      _EVAL_272 <= 32'h0;
    end else begin
      _EVAL_272 <= _EVAL_36;
    end
    if (_EVAL_126) begin
      _EVAL_276 <= _EVAL_14;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbd9a7e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c31961f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3552a909)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(877a037)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1404e59c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(455c22b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c2dd6c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7d74ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91e2ee74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(564047e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(573b31e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e71d71e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abac0efc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b983ae8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9acc5a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbd9a7e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a704a24b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(160629bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11f271cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbdebe72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffb5157e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca074c93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ebe3882f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3de35d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_275) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e995a7fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(141bca40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45ea1eb6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2b1e751)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9226677)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfadc7ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e2142b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a150bd81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e38ffe8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd07f2b3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1833ea67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a35ad612)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_3 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a3a2f97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(218fdee7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(277ba35e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f3f459f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e649a9aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(697af2ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_23 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(362dbec1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c735a92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7686e1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1f853fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edb6e7a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_202 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c01c2f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b187cb36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ea9877)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f48df8ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_35) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94858b88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19770407)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e3cefc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_107) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2408b005)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(191531e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_107) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e476b745)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ee7b09d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8df111a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_275) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_24) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afca74db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bd8d7bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_227) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b082ac21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5cea072)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6b5dff4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b2a218a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_129) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc5a9419)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc93bcc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d20bc61f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7664c53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_41 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e62b2338)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b8ca31a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_166 & _EVAL_129) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c84ead5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_35) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9e295b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1bd1ba41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_24) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7409695)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be6556fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_16 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_48 = _RAND_1[14:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_75 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_80 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_89 = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_98 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_162 = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_181 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_222 = _RAND_8[17:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_223 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_264 = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_268 = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_272 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_276 = _RAND_13[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
