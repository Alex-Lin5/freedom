//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_23_assert(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input  [3:0]  _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [2:0]  _EVAL_9,
  input  [3:0]  _EVAL_10,
  input         _EVAL_11,
  input  [1:0]  _EVAL_12,
  input  [3:0]  _EVAL_13,
  input  [31:0] _EVAL_14
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_15;
  wire [32:0] _EVAL_16;
  wire [32:0] _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire [5:0] _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire [32:0] _EVAL_24;
  wire [32:0] _EVAL_25;
  wire  _EVAL_26;
  wire [7:0] _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  reg  _EVAL_30;
  wire [32:0] _EVAL_31;
  wire [31:0] _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_36;
  wire [3:0] _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_42;
  wire [31:0] _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire [22:0] _EVAL_46;
  wire [31:0] _EVAL_47;
  reg [31:0] _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire [32:0] _EVAL_57;
  wire  _EVAL_58;
  wire [32:0] _EVAL_59;
  wire [1:0] _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire [5:0] _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire [5:0] _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire [32:0] _EVAL_82;
  wire [1:0] _EVAL_83;
  wire [32:0] _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire [32:0] _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  reg [5:0] _EVAL_91;
  wire  _EVAL_92;
  reg [3:0] _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire [22:0] _EVAL_98;
  wire [7:0] _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire [32:0] _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  reg  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire [7:0] _EVAL_113;
  wire [5:0] _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire [31:0] _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  reg [2:0] _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire [32:0] _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire [32:0] _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  reg  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire [5:0] _EVAL_147;
  wire  _EVAL_148;
  wire [32:0] _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire [31:0] _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire [32:0] _EVAL_163;
  wire  _EVAL_164;
  wire [32:0] _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire [31:0] _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire [32:0] _EVAL_184;
  wire  _EVAL_185;
  wire [7:0] _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire [3:0] _EVAL_198;
  wire [6:0] _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire [6:0] _EVAL_203;
  wire  _EVAL_204;
  wire [3:0] _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire [1:0] _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  reg [3:0] _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire [32:0] _EVAL_218;
  wire  _EVAL_219;
  wire [32:0] _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire [31:0] _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire [31:0] _EVAL_228;
  wire [31:0] _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire [32:0] _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  reg [1:0] _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  reg [5:0] _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire [6:0] _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire [32:0] _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire [32:0] _EVAL_253;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire [31:0] _EVAL_263;
  wire  _EVAL_264;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_265;
  reg [5:0] _EVAL_266;
  wire  _EVAL_268;
  wire [6:0] _EVAL_269;
  wire [32:0] _EVAL_270;
  wire [3:0] _EVAL_271;
  wire [32:0] _EVAL_272;
  wire [32:0] _EVAL_273;
  wire  _EVAL_274;
  wire [5:0] _EVAL_275;
  wire  _EVAL_276;
  wire [1:0] _EVAL_277;
  wire  _EVAL_278;
  reg [5:0] _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_285;
  wire  _EVAL_286;
  reg [2:0] _EVAL_287;
  wire  _EVAL_288;
  reg [31:0] _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_295;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_17 = $signed(_EVAL_103) & -33'sh1000;
  assign _EVAL_19 = _EVAL_1 == _EVAL_106;
  assign _EVAL_109 = _EVAL_0 == 3'h5;
  assign _EVAL_150 = _EVAL_12 <= 2'h2;
  assign _EVAL_278 = _EVAL_182 | _EVAL;
  assign _EVAL_268 = _EVAL_8 & _EVAL_295;
  assign _EVAL_69 = ~_EVAL_230;
  assign _EVAL_257 = _EVAL_141 & _EVAL_80;
  assign _EVAL_171 = _EVAL_9 == 3'h4;
  assign _EVAL_212 = _EVAL_185 | _EVAL;
  assign _EVAL_55 = _EVAL_11 & _EVAL_154;
  assign _EVAL_293 = _EVAL_63 & _EVAL_191;
  assign _EVAL_28 = _EVAL_8 & _EVAL_53;
  assign _EVAL_208 = 2'h1 << _EVAL_259;
  assign _EVAL_44 = _EVAL_11 & _EVAL_109;
  assign _EVAL_119 = _EVAL_62 | _EVAL_73;
  assign _EVAL_152 = ~_EVAL_212;
  assign _EVAL_290 = ~_EVAL_197;
  assign _EVAL_221 = ~_EVAL_170;
  assign _EVAL_95 = _EVAL_131 | _EVAL_293;
  assign _EVAL_63 = _EVAL_83[1];
  assign _EVAL_149 = {1'b0,$signed(_EVAL_172)};
  assign _EVAL_64 = _EVAL_265 & _EVAL_258;
  assign _EVAL_138 = _EVAL_12 == 2'h0;
  assign _EVAL_244 = _EVAL_0 == 3'h1;
  assign _EVAL_190 = ~_EVAL_202;
  assign _EVAL_216 = _EVAL_63 & _EVAL_74;
  assign _EVAL_139 = _EVAL_9 == 3'h5;
  assign _EVAL_114 = _EVAL_27[7:2];
  assign _EVAL_22 = _EVAL_11 & _EVAL_187;
  assign _EVAL_258 = _EVAL_240 == 6'h0;
  assign _EVAL_276 = _EVAL_11 & _EVAL_251;
  assign _EVAL_178 = ~_EVAL_176;
  assign _EVAL_27 = ~_EVAL_186;
  assign _EVAL_51 = _EVAL_8 & _EVAL_122;
  assign _EVAL_193 = _EVAL_224 | _EVAL_5;
  assign _EVAL_115 = _EVAL_217 | _EVAL;
  assign _EVAL_136 = _EVAL_189 | _EVAL_54;
  assign _EVAL_103 = {1'b0,$signed(_EVAL_263)};
  assign _EVAL_231 = _EVAL_13 <= 4'h6;
  assign _EVAL_186 = _EVAL_98[7:0];
  assign _EVAL_133 = _EVAL_261 & _EVAL_39;
  assign _EVAL_213 = _EVAL_37 == 4'h0;
  assign _EVAL_141 = _EVAL_13 <= 4'h8;
  assign _EVAL_20 = _EVAL_199[5:0];
  assign _EVAL_202 = _EVAL_150 | _EVAL;
  assign _EVAL_187 = _EVAL_0 == 3'h2;
  assign _EVAL_220 = $signed(_EVAL_149) & -33'sh400000;
  assign _EVAL_67 = _EVAL_13 == _EVAL_214;
  assign _EVAL_163 = _EVAL_184;
  assign _EVAL_81 = _EVAL_11 & _EVAL_164;
  assign _EVAL_263 = _EVAL_14 ^ 32'h3000;
  assign _EVAL_57 = _EVAL_24;
  assign _EVAL_277 = _EVAL_129 ? 2'h1 : 2'h0;
  assign _EVAL_92 = |_EVAL_108;
  assign _EVAL_100 = ~_EVAL_113;
  assign _EVAL_140 = _EVAL_138 | _EVAL;
  assign _EVAL_53 = _EVAL_9 == 3'h6;
  assign _EVAL_234 = _EVAL_8 & _EVAL_171;
  assign _EVAL_272 = _EVAL_220;
  assign _EVAL_36 = ~_EVAL_101;
  assign _EVAL_188 = _EVAL_8 & _EVAL_239;
  assign _EVAL_70 = ~_EVAL_251;
  assign _EVAL_31 = $signed(_EVAL_218) & -33'sh4000;
  assign _EVAL_249 = _EVAL_279 == 6'h0;
  assign _EVAL_123 = _EVAL_8 & _EVAL_139;
  assign _EVAL_246 = ~_EVAL_219;
  assign _EVAL_86 = _EVAL_116 | _EVAL_286;
  assign _EVAL_210 = _EVAL_108 != _EVAL_227;
  assign _EVAL_76 = |_EVAL_30;
  assign _EVAL_248 = _EVAL_9 == _EVAL_287;
  assign _EVAL_189 = _EVAL_119 | _EVAL_126;
  assign _EVAL_160 = _EVAL_14 ^ 32'h80000000;
  assign _EVAL_151 = ~_EVAL_115;
  assign _EVAL_108 = _EVAL_61[0];
  assign _EVAL_274 = _EVAL_281 | _EVAL;
  assign _EVAL_222 = _EVAL_252 | _EVAL;
  assign _EVAL_62 = $signed(_EVAL_165) == 33'sh0;
  assign _EVAL_154 = _EVAL_0 == 3'h0;
  assign _EVAL_197 = _EVAL_262 | _EVAL;
  assign _EVAL_262 = _EVAL_210 | _EVAL_169;
  assign _EVAL_25 = _EVAL_17;
  assign _EVAL_180 = _EVAL_0 == 3'h4;
  assign _EVAL_229 = _EVAL_14 ^ 32'h40000000;
  assign _EVAL_68 = _EVAL_245[5:0];
  assign _EVAL_147 = _EVAL_100[7:2];
  assign _EVAL_144 = _EVAL_231 & _EVAL_209;
  assign _EVAL_46 = 23'hff << _EVAL_13;
  assign _EVAL_166 = _EVAL_77 & _EVAL_249;
  assign _EVAL_174 = _EVAL_86 | _EVAL_110;
  assign _EVAL_126 = $signed(_EVAL_57) == 33'sh0;
  assign _EVAL_77 = _EVAL_2 & _EVAL_11;
  assign _EVAL_170 = _EVAL_264 | _EVAL;
  assign _EVAL_157 = _EVAL_18 & _EVAL_52;
  assign _EVAL_295 = _EVAL_9 == 3'h7;
  assign _EVAL_291 = ~_EVAL_104;
  assign _EVAL_245 = _EVAL_266 - 6'h1;
  assign _EVAL_29 = ~_EVAL_274;
  assign _EVAL_285 = _EVAL_175 | _EVAL_42;
  assign _EVAL_38 = _EVAL_11 & _EVAL_180;
  assign _EVAL_280 = _EVAL_18 & _EVAL_183;
  assign _EVAL_206 = ~_EVAL_107;
  assign _EVAL_238 = ~_EVAL_241;
  assign _EVAL_130 = _EVAL_45 | _EVAL;
  assign _EVAL_217 = _EVAL_257 | _EVAL_194;
  assign _EVAL_270 = {1'b0,$signed(_EVAL_228)};
  assign _EVAL_65 = _EVAL_203[5:0];
  assign _EVAL_283 = _EVAL_102 | _EVAL;
  assign _EVAL_264 = _EVAL_47 == 32'h0;
  assign _EVAL_43 = _EVAL_14 ^ 32'h2000000;
  assign _EVAL_227 = _EVAL_277[0];
  assign _EVAL_45 = _EVAL_108 | _EVAL_30;
  assign _EVAL_75 = _EVAL_174 | _EVAL;
  assign _EVAL_256 = _EVAL_255 | _EVAL_280;
  assign _EVAL_125 = _EVAL_265 | _EVAL_77;
  assign _EVAL_122 = _EVAL_9 == 3'h3;
  assign _EVAL_113 = _EVAL_46[7:0];
  assign _EVAL_237 = ~_EVAL_233;
  assign _EVAL_85 = ~_EVAL;
  assign _EVAL_132 = _EVAL_48 + 32'h1;
  assign _EVAL_79 = ~_EVAL_90;
  assign _EVAL_90 = _EVAL_168 | _EVAL;
  assign _EVAL_198 = {_EVAL_134,_EVAL_40,_EVAL_256,_EVAL_192};
  assign _EVAL_173 = ~_EVAL_5;
  assign _EVAL_162 = _EVAL_0[0];
  assign _EVAL_47 = _EVAL_14 & _EVAL_121;
  assign _EVAL_82 = _EVAL_250;
  assign _EVAL_172 = _EVAL_14 ^ 32'hc000000;
  assign _EVAL_58 = ~_EVAL_112;
  assign _EVAL_204 = _EVAL_213 | _EVAL;
  assign _EVAL_121 = {{24'd0}, _EVAL_100};
  assign _EVAL_80 = $signed(_EVAL_25) == 33'sh0;
  assign _EVAL_201 = ~_EVAL_75;
  assign _EVAL_184 = $signed(_EVAL_270) & -33'sh2000;
  assign _EVAL_54 = $signed(_EVAL_272) == 33'sh0;
  assign _EVAL_40 = _EVAL_95 | _EVAL_157;
  assign _EVAL_146 = _EVAL_173 | _EVAL;
  assign _EVAL_72 = ~_EVAL_23;
  assign _EVAL_223 = _EVAL_14 ^ 32'h1800000;
  assign _EVAL_183 = _EVAL_74 & _EVAL_247;
  assign _EVAL_161 = ~_EVAL_30;
  assign _EVAL_235 = _EVAL_77 & _EVAL_21;
  assign _EVAL_194 = _EVAL_231 & _EVAL_128;
  assign _EVAL_110 = _EVAL_48 < plusarg_reader_out;
  assign _EVAL_247 = _EVAL_14[0];
  assign _EVAL_87 = $signed(_EVAL_273) & -33'sh2000;
  assign _EVAL_252 = _EVAL_14 == _EVAL_289;
  assign _EVAL_131 = _EVAL_13 >= 4'h2;
  assign _EVAL_232 = _EVAL_31;
  assign _EVAL_185 = _EVAL_0 <= 3'h6;
  assign _EVAL_225 = _EVAL_226 | _EVAL;
  assign _EVAL_105 = ~_EVAL_130;
  assign _EVAL_107 = _EVAL_19 | _EVAL;
  assign _EVAL_176 = _EVAL_288 | _EVAL;
  assign _EVAL_78 = ~_EVAL_181;
  assign _EVAL_195 = _EVAL_13 <= 4'h2;
  assign _EVAL_164 = ~_EVAL_249;
  assign _EVAL_243 = _EVAL_94 | _EVAL;
  assign _EVAL_128 = _EVAL_156 | _EVAL_26;
  assign _EVAL_102 = _EVAL_6 >= 4'h2;
  assign _EVAL_145 = _EVAL_136 | _EVAL_175;
  assign _EVAL_281 = _EVAL_0 == _EVAL_124;
  assign _EVAL_167 = _EVAL_271 == 4'h0;
  assign _EVAL_265 = _EVAL_7 & _EVAL_8;
  assign _EVAL_117 = _EVAL_161 | _EVAL;
  assign _EVAL_199 = _EVAL_240 - 6'h1;
  assign _EVAL_26 = $signed(_EVAL_232) == 33'sh0;
  assign _EVAL_228 = _EVAL_14 ^ 32'h20000000;
  assign _EVAL_286 = plusarg_reader_out == 32'h0;
  assign _EVAL_33 = _EVAL_11 & _EVAL_244;
  assign _EVAL_16 = $signed(_EVAL_253) & -33'sh5000;
  assign _EVAL_34 = ~_EVAL_204;
  assign _EVAL_169 = ~_EVAL_92;
  assign _EVAL_230 = _EVAL_9[2];
  assign _EVAL_226 = _EVAL_195 & _EVAL_217;
  assign _EVAL_271 = ~_EVAL_10;
  assign _EVAL_207 = _EVAL_10 == _EVAL_198;
  assign _EVAL_32 = _EVAL_132[31:0];
  assign _EVAL_273 = {1'b0,$signed(_EVAL_229)};
  assign _EVAL_288 = _EVAL_12 == _EVAL_236;
  assign _EVAL_233 = _EVAL_193 | _EVAL;
  assign _EVAL_61 = _EVAL_64 ? 2'h1 : 2'h0;
  assign _EVAL_269 = _EVAL_279 - 6'h1;
  assign _EVAL_241 = _EVAL_195 | _EVAL;
  assign _EVAL_260 = _EVAL_18 & _EVAL_148;
  assign _EVAL_239 = ~_EVAL_215;
  assign _EVAL_292 = _EVAL_8 & _EVAL_49;
  assign _EVAL_242 = ~_EVAL_196;
  assign _EVAL_18 = _EVAL_83[0];
  assign _EVAL_49 = _EVAL_9 == 3'h1;
  assign _EVAL_192 = _EVAL_255 | _EVAL_15;
  assign _EVAL_215 = _EVAL_91 == 6'h0;
  assign _EVAL_251 = _EVAL_0 == 3'h6;
  assign _EVAL_94 = _EVAL_257 | _EVAL_137;
  assign _EVAL_52 = _EVAL_191 & _EVAL_179;
  assign _EVAL_104 = _EVAL_97 | _EVAL;
  assign _EVAL_88 = ~_EVAL_140;
  assign _EVAL_224 = ~_EVAL_1;
  assign _EVAL_200 = _EVAL_224 | _EVAL;
  assign _EVAL_219 = _EVAL_211 | _EVAL;
  assign _EVAL_129 = _EVAL_235 & _EVAL_70;
  assign _EVAL_21 = _EVAL_266 == 6'h0;
  assign _EVAL_83 = _EVAL_208 | 2'h1;
  assign _EVAL_177 = _EVAL_8 & _EVAL_282;
  assign _EVAL_250 = $signed(_EVAL_59) & -33'sh4000;
  assign _EVAL_135 = _EVAL_87;
  assign _EVAL_84 = {1'b0,$signed(_EVAL_43)};
  assign _EVAL_37 = _EVAL_10 & _EVAL_205;
  assign _EVAL_159 = ~_EVAL_117;
  assign _EVAL_179 = ~_EVAL_247;
  assign _EVAL_23 = _EVAL_248 | _EVAL;
  assign _EVAL_116 = ~_EVAL_76;
  assign _EVAL_89 = ~_EVAL_146;
  assign _EVAL_259 = _EVAL_13[0];
  assign _EVAL_218 = {1'b0,$signed(_EVAL_160)};
  assign _EVAL_191 = _EVAL_14[1];
  assign _EVAL_196 = _EVAL_67 | _EVAL;
  assign _EVAL_282 = _EVAL_9 == 3'h0;
  assign _EVAL_127 = ~_EVAL_243;
  assign _EVAL_112 = _EVAL_131 | _EVAL;
  assign _EVAL_205 = ~_EVAL_198;
  assign _EVAL_261 = _EVAL_30 | _EVAL_108;
  assign _EVAL_24 = $signed(_EVAL_84) & -33'sh10000;
  assign _EVAL_66 = _EVAL_9 == 3'h2;
  assign _EVAL_158 = ~_EVAL_278;
  assign _EVAL_134 = _EVAL_95 | _EVAL_260;
  assign _EVAL_111 = ~_EVAL_200;
  assign _EVAL_175 = $signed(_EVAL_163) == 33'sh0;
  assign _EVAL_15 = _EVAL_18 & _EVAL_96;
  assign _EVAL_203 = _EVAL_91 - 6'h1;
  assign _EVAL_155 = ~_EVAL_225;
  assign _EVAL_101 = _EVAL_207 | _EVAL;
  assign _EVAL_96 = _EVAL_74 & _EVAL_179;
  assign _EVAL_97 = _EVAL_12 != 2'h2;
  assign _EVAL_211 = _EVAL_4 == _EVAL_143;
  assign _EVAL_165 = _EVAL_16;
  assign _EVAL_275 = _EVAL_269[5:0];
  assign _EVAL_98 = 23'hff << _EVAL_6;
  assign _EVAL_142 = _EVAL_265 & _EVAL_215;
  assign _EVAL_74 = ~_EVAL_191;
  assign _EVAL_168 = _EVAL_257 | _EVAL_144;
  assign _EVAL_209 = _EVAL_136 | _EVAL_26;
  assign _EVAL_255 = _EVAL_131 | _EVAL_216;
  assign _EVAL_153 = ~_EVAL_222;
  assign _EVAL_156 = _EVAL_145 | _EVAL_42;
  assign _EVAL_59 = {1'b0,$signed(_EVAL_223)};
  assign _EVAL_73 = $signed(_EVAL_82) == 33'sh0;
  assign _EVAL_50 = ~_EVAL_283;
  assign _EVAL_137 = _EVAL_231 & _EVAL_285;
  assign _EVAL_120 = _EVAL_8 & _EVAL_66;
  assign _EVAL_148 = _EVAL_191 & _EVAL_247;
  assign _EVAL_253 = {1'b0,$signed(_EVAL_14)};
  assign _EVAL_42 = $signed(_EVAL_135) == 33'sh0;
  assign _EVAL_182 = _EVAL_6 == _EVAL_93;
  assign _EVAL_181 = _EVAL_167 | _EVAL;
  assign _EVAL_39 = ~_EVAL_227;
  always @(posedge _EVAL_3) begin
    if (_EVAL) begin
      _EVAL_30 <= 1'h0;
    end else begin
      _EVAL_30 <= _EVAL_133;
    end
    if (_EVAL) begin
      _EVAL_48 <= 32'h0;
    end else if (_EVAL_125) begin
      _EVAL_48 <= 32'h0;
    end else begin
      _EVAL_48 <= _EVAL_32;
    end
    if (_EVAL) begin
      _EVAL_91 <= 6'h0;
    end else if (_EVAL_265) begin
      if (_EVAL_215) begin
        if (_EVAL_69) begin
          _EVAL_91 <= _EVAL_147;
        end else begin
          _EVAL_91 <= 6'h0;
        end
      end else begin
        _EVAL_91 <= _EVAL_65;
      end
    end
    if (_EVAL_166) begin
      _EVAL_93 <= _EVAL_6;
    end
    if (_EVAL_166) begin
      _EVAL_106 <= _EVAL_1;
    end
    if (_EVAL_166) begin
      _EVAL_124 <= _EVAL_0;
    end
    if (_EVAL_166) begin
      _EVAL_143 <= _EVAL_4;
    end
    if (_EVAL_142) begin
      _EVAL_214 <= _EVAL_13;
    end
    if (_EVAL_166) begin
      _EVAL_236 <= _EVAL_12;
    end
    if (_EVAL) begin
      _EVAL_240 <= 6'h0;
    end else if (_EVAL_265) begin
      if (_EVAL_258) begin
        if (_EVAL_69) begin
          _EVAL_240 <= _EVAL_147;
        end else begin
          _EVAL_240 <= 6'h0;
        end
      end else begin
        _EVAL_240 <= _EVAL_20;
      end
    end
    if (_EVAL) begin
      _EVAL_266 <= 6'h0;
    end else if (_EVAL_77) begin
      if (_EVAL_21) begin
        if (_EVAL_162) begin
          _EVAL_266 <= _EVAL_114;
        end else begin
          _EVAL_266 <= 6'h0;
        end
      end else begin
        _EVAL_266 <= _EVAL_68;
      end
    end
    if (_EVAL) begin
      _EVAL_279 <= 6'h0;
    end else if (_EVAL_77) begin
      if (_EVAL_249) begin
        if (_EVAL_162) begin
          _EVAL_279 <= _EVAL_114;
        end else begin
          _EVAL_279 <= 6'h0;
        end
      end else begin
        _EVAL_279 <= _EVAL_275;
      end
    end
    if (_EVAL_142) begin
      _EVAL_287 <= _EVAL_9;
    end
    if (_EVAL_142) begin
      _EVAL_289 <= _EVAL_14;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_237) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_34) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb38aa00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(196965b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_34) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c748d81a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5335eefc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e92c8cf5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0ebd37e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5834e05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2b62259)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_155) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb76526e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32149494)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab341295)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc5dd0f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97fa6dbe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da99645f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d1b0c5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa3beb73)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8cbae113)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(232e637a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7305a98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf631267)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45354780)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d367052)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_237) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(672cca0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37f92993)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_79) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(631227c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98f444df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d34d115)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6380074d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b5a0f06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52a1b109)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86a75040)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49a99fb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f8ea883)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ade29e72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_155) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(721b0970)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e1399af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c320226)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(faf1d23b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8973ef18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28913d3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4da24bb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_237) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b91eb5ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_129 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb8610b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5adf5346)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74da1502)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_177 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6810a024)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d1d23a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3f9c70e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63502a1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(311194)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7e0dd1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(678c28a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9eb8386d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_221) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f368e7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c183b117)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(594c31d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_221) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(714464bf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_85) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_79) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_88) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a78c67d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(881ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_242) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e96966)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_242) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_64 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_238) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72d98bda)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_88) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6502ece9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35aac0da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_268 & _EVAL_85) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4da24bb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_234 & _EVAL_238) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_237) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e374b611)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_188 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_30 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_48 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_91 = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_93 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_106 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_124 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_143 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_214 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_236 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_240 = _RAND_9[5:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_266 = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_279 = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_287 = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_289 = _RAND_13[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
