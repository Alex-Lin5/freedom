//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_110(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  output        _EVAL_2,
  output [31:0] _EVAL_3,
  output        _EVAL_4,
  output        _EVAL_5,
  input  [3:0]  _EVAL_6,
  input  [1:0]  _EVAL_7,
  input  [29:0] _EVAL_8,
  output [31:0] _EVAL_9,
  input         _EVAL_10,
  output        _EVAL_11,
  input         _EVAL_12,
  output        _EVAL_13,
  input  [1:0]  _EVAL_14,
  input         _EVAL_15,
  input  [31:0] _EVAL_16,
  input         _EVAL_17,
  output [2:0]  _EVAL_18,
  input         _EVAL_19,
  output        _EVAL_20,
  input  [1:0]  _EVAL_21,
  input  [31:0] _EVAL_22,
  input         _EVAL_23,
  output [6:0]  _EVAL_24,
  output        _EVAL_25,
  output        _EVAL_26,
  output        _EVAL_27,
  output        _EVAL_28,
  input         _EVAL_29,
  input         _EVAL_30,
  output        _EVAL_31,
  input         _EVAL_32,
  output        _EVAL_33,
  output        _EVAL_34,
  input  [2:0]  _EVAL_35,
  input         _EVAL_36,
  input  [29:0] _EVAL_37,
  output [31:0] _EVAL_38,
  input  [31:0] _EVAL_39,
  input         _EVAL_40,
  input         _EVAL_41,
  input  [31:0] _EVAL_42,
  input         _EVAL_43,
  input         _EVAL_44,
  input         _EVAL_45,
  input         _EVAL_46,
  input         _EVAL_47,
  input         _EVAL_48,
  input         _EVAL_49,
  output        _EVAL_50,
  input  [2:0]  _EVAL_51,
  input  [31:0] _EVAL_52,
  output        _EVAL_53,
  output [31:0] _EVAL_54,
  input  [1:0]  _EVAL_55,
  output        _EVAL_56,
  input  [31:0] _EVAL_57,
  input  [31:0] _EVAL_58,
  input  [29:0] _EVAL_59,
  input  [1:0]  _EVAL_60,
  input  [29:0] _EVAL_61,
  input         _EVAL_62,
  input         _EVAL_63,
  output [3:0]  _EVAL_64,
  input  [1:0]  _EVAL_65,
  input  [1:0]  _EVAL_66,
  input  [1:0]  _EVAL_67,
  input         _EVAL_68,
  output        _EVAL_69,
  output        _EVAL_70,
  input  [29:0] _EVAL_71,
  output        _EVAL_72,
  input         _EVAL_73,
  input         _EVAL_74,
  input         _EVAL_75,
  input  [31:0] _EVAL_76,
  input  [6:0]  _EVAL_77,
  input  [29:0] _EVAL_78,
  output [3:0]  _EVAL_79,
  input         _EVAL_80,
  input  [29:0] _EVAL_81,
  input  [1:0]  _EVAL_82,
  output        _EVAL_83,
  input         _EVAL_84,
  input  [31:0] _EVAL_85,
  output        _EVAL_86,
  input  [3:0]  _EVAL_87,
  input         _EVAL_88,
  output [1:0]  _EVAL_89,
  input  [31:0] _EVAL_90,
  input  [29:0] _EVAL_91,
  input  [31:0] _EVAL_92,
  input         _EVAL_93,
  input         _EVAL_94,
  output [3:0]  _EVAL_95,
  input  [1:0]  _EVAL_96,
  input         _EVAL_97,
  input  [4:0]  _EVAL_98,
  output        _EVAL_99,
  output [31:0] _EVAL_100,
  output        _EVAL_101,
  output        _EVAL_102,
  input         _EVAL_103,
  input         _EVAL_104,
  input         _EVAL_105,
  output [2:0]  _EVAL_106,
  output [1:0]  _EVAL_107,
  input         _EVAL_108,
  input         _EVAL_109,
  input         _EVAL_110,
  input  [1:0]  _EVAL_111,
  input         _EVAL_112,
  input         _EVAL_113,
  output [31:0] _EVAL_114,
  input  [3:0]  _EVAL_115,
  output        _EVAL_116,
  output        _EVAL_117,
  input         _EVAL_118,
  output [31:0] _EVAL_119,
  input         _EVAL_120,
  input         _EVAL_121,
  input  [1:0]  _EVAL_122,
  input         _EVAL_123,
  output [4:0]  _EVAL_124,
  input  [31:0] _EVAL_125,
  input         _EVAL_126,
  output [2:0]  _EVAL_127,
  output        _EVAL_128
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire [6:0] _EVAL_133;
  wire [31:0] _EVAL_134;
  wire  _EVAL_135;
  wire [13:0] _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire [3:0] _EVAL_139;
  wire [31:0] _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire [1:0] _EVAL_144;
  wire [1:0] _EVAL_145;
  wire  _EVAL_146;
  wire [1:0] _EVAL_147;
  wire  pma_checker_pmp__EVAL;
  wire [31:0] pma_checker_pmp__EVAL_0;
  wire [29:0] pma_checker_pmp__EVAL_1;
  wire  pma_checker_pmp__EVAL_2;
  wire  pma_checker_pmp__EVAL_3;
  wire  pma_checker_pmp__EVAL_4;
  wire [29:0] pma_checker_pmp__EVAL_5;
  wire  pma_checker_pmp__EVAL_6;
  wire [1:0] pma_checker_pmp__EVAL_7;
  wire  pma_checker_pmp__EVAL_8;
  wire  pma_checker_pmp__EVAL_9;
  wire [1:0] pma_checker_pmp__EVAL_10;
  wire [1:0] pma_checker_pmp__EVAL_11;
  wire [1:0] pma_checker_pmp__EVAL_12;
  wire  pma_checker_pmp__EVAL_13;
  wire  pma_checker_pmp__EVAL_14;
  wire  pma_checker_pmp__EVAL_15;
  wire [1:0] pma_checker_pmp__EVAL_16;
  wire  pma_checker_pmp__EVAL_17;
  wire  pma_checker_pmp__EVAL_18;
  wire  pma_checker_pmp__EVAL_19;
  wire [29:0] pma_checker_pmp__EVAL_20;
  wire  pma_checker_pmp__EVAL_21;
  wire  pma_checker_pmp__EVAL_22;
  wire  pma_checker_pmp__EVAL_23;
  wire [31:0] pma_checker_pmp__EVAL_24;
  wire  pma_checker_pmp__EVAL_25;
  wire  pma_checker_pmp__EVAL_26;
  wire [31:0] pma_checker_pmp__EVAL_27;
  wire [31:0] pma_checker_pmp__EVAL_28;
  wire [31:0] pma_checker_pmp__EVAL_29;
  wire  pma_checker_pmp__EVAL_30;
  wire [1:0] pma_checker_pmp__EVAL_31;
  wire [1:0] pma_checker_pmp__EVAL_32;
  wire [29:0] pma_checker_pmp__EVAL_33;
  wire [31:0] pma_checker_pmp__EVAL_34;
  wire  pma_checker_pmp__EVAL_35;
  wire  pma_checker_pmp__EVAL_36;
  wire  pma_checker_pmp__EVAL_37;
  wire [31:0] pma_checker_pmp__EVAL_38;
  wire [31:0] pma_checker_pmp__EVAL_39;
  wire [1:0] pma_checker_pmp__EVAL_40;
  wire [29:0] pma_checker_pmp__EVAL_41;
  wire [29:0] pma_checker_pmp__EVAL_42;
  wire  pma_checker_pmp__EVAL_43;
  wire  pma_checker_pmp__EVAL_44;
  wire [29:0] pma_checker_pmp__EVAL_45;
  wire [31:0] pma_checker_pmp__EVAL_46;
  wire [1:0] pma_checker_pmp__EVAL_47;
  wire  pma_checker_pmp__EVAL_48;
  wire  pma_checker_pmp__EVAL_49;
  wire  pma_checker_pmp__EVAL_50;
  wire  pma_checker_pmp__EVAL_51;
  wire  pma_checker_pmp__EVAL_52;
  wire [29:0] pma_checker_pmp__EVAL_53;
  wire  pma_checker_pmp__EVAL_54;
  wire  pma_checker_pmp__EVAL_55;
  wire  pma_checker_pmp__EVAL_56;
  wire  pma_checker_pmp__EVAL_57;
  wire  pma_checker_pmp__EVAL_58;
  wire  pma_checker_pmp__EVAL_59;
  wire  pma_checker_pmp__EVAL_60;
  wire  pma_checker_pmp__EVAL_61;
  wire [3:0] _EVAL_148;
  wire  _EVAL_149;
  wire [2:0] _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire [3:0] _EVAL_154;
  wire [5:0] _EVAL_155;
  wire  _EVAL_156;
  wire [32:0] _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire [2:0] _EVAL_160;
  wire [31:0] _EVAL_161;
  wire  _EVAL_163;
  wire [2:0] _EVAL_164;
  wire [1:0] _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire [13:0] _EVAL_168;
  wire  _EVAL_169;
  wire [31:0] _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire [3:0] _EVAL_174;
  wire  _EVAL_176;
  wire [6:0] _EVAL_177;
  wire [31:0] _EVAL_178;
  wire [31:0] _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_182;
  wire [6:0] _EVAL_183;
  wire  _EVAL_185;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire [6:0] _EVAL_189;
  wire [31:0] _EVAL_190;
  wire  _EVAL_191;
  wire [31:0] _EVAL_192;
  wire  _EVAL_193;
  wire [2:0] _EVAL_194;
  wire  _EVAL_195;
  wire [3:0] _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire [1:0] _EVAL_199;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire [2:0] _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_207;
  wire [32:0] _EVAL_208;
  wire [1:0] _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire [1:0] _EVAL_213;
  wire [15:0] _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire [2:0] _EVAL_219;
  wire [31:0] _EVAL_220;
  wire  _EVAL_221;
  wire [29:0] _EVAL_222;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire [13:0] _EVAL_227;
  wire [7:0] _EVAL_228;
  wire [6:0] _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire [31:0] _EVAL_234;
  wire [31:0] _EVAL_236;
  wire [3:0] _EVAL_237;
  wire  _EVAL_238;
  wire [31:0] _EVAL_239;
  wire [3:0] _EVAL_240;
  wire [2:0] _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire [15:0] _EVAL_248;
  wire  _EVAL_249;
  wire [1:0] _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire [13:0] _EVAL_256;
  wire [13:0] _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire [15:0] _EVAL_262;
  wire [31:0] _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire [32:0] _EVAL_267;
  wire  _EVAL_268;
  wire [31:0] _EVAL_269;
  wire [29:0] _EVAL_270;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire [13:0] _EVAL_274;
  wire [1:0] _EVAL_275;
  wire [1:0] _EVAL_276;
  wire [2:0] _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire [32:0] _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire [31:0] _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire [2:0] _EVAL_289;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire [32:0] _EVAL_293;
  wire [13:0] _EVAL_294;
  wire  _EVAL_295;
  wire  _EVAL_297;
  wire [7:0] _EVAL_298;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire [32:0] _EVAL_302;
  wire  _EVAL_303;
  wire [31:0] _EVAL_304;
  wire  _EVAL_305;
  wire [3:0] _EVAL_306;
  wire  _EVAL_307;
  wire [31:0] _EVAL_308;
  wire  _EVAL_309;
  wire [1:0] _EVAL_310;
  wire  _EVAL_311;
  wire  _EVAL_312;
  wire [31:0] _EVAL_313;
  wire [31:0] _EVAL_314;
  wire  _EVAL_316;
  wire [31:0] _EVAL_317;
  wire [11:0] _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_320;
  wire  data__EVAL;
  wire [3:0] data__EVAL_0;
  wire [13:0] data__EVAL_1;
  wire [31:0] data__EVAL_2;
  wire [31:0] data__EVAL_3;
  wire  data__EVAL_4;
  wire  data__EVAL_5;
  wire [31:0] _EVAL_321;
  wire  _EVAL_322;
  wire [3:0] _EVAL_323;
  wire  _EVAL_324;
  wire  _EVAL_326;
  wire [3:0] _EVAL_327;
  wire [3:0] _EVAL_328;
  wire  _EVAL_329;
  wire  _EVAL_331;
  wire  _EVAL_332;
  wire  _EVAL_333;
  wire [1:0] _EVAL_334;
  wire [32:0] _EVAL_335;
  wire  _EVAL_336;
  wire  _EVAL_337;
  wire  _EVAL_338;
  wire  _EVAL_339;
  wire [32:0] _EVAL_340;
  wire  _EVAL_341;
  wire  _EVAL_342;
  wire [5:0] _EVAL_343;
  wire [15:0] _EVAL_344;
  wire [1:0] _EVAL_345;
  wire [32:0] _EVAL_346;
  wire  _EVAL_347;
  wire [19:0] _EVAL_348;
  wire  _EVAL_349;
  wire  _EVAL_350;
  wire  _EVAL_351;
  wire [32:0] _EVAL_352;
  wire [31:0] _EVAL_353;
  wire [5:0] _EVAL_354;
  wire  _EVAL_356;
  wire [3:0] _EVAL_357;
  wire [6:0] _EVAL_358;
  wire [13:0] _EVAL_359;
  wire [31:0] _EVAL_361;
  wire [3:0] _EVAL_362;
  wire  _EVAL_363;
  wire [2:0] _EVAL_364;
  wire  _EVAL_365;
  wire  _EVAL_367;
  wire  _EVAL_368;
  wire [2:0] _EVAL_369;
  wire  _EVAL_370;
  wire  _EVAL_371;
  wire [32:0] _EVAL_372;
  wire [13:0] _EVAL_373;
  wire [13:0] _EVAL_374;
  wire  _EVAL_376;
  wire  _EVAL_377;
  wire [3:0] _EVAL_378;
  wire [31:0] _EVAL_379;
  wire [2:0] _EVAL_380;
  wire [1:0] _EVAL_381;
  wire [2:0] _EVAL_383;
  wire [7:0] _EVAL_384;
  wire [7:0] _EVAL_385;
  wire  _EVAL_386;
  wire  _EVAL_387;
  wire  _EVAL_388;
  wire  _EVAL_389;
  wire  _EVAL_390;
  wire [13:0] _EVAL_391;
  wire [32:0] _EVAL_392;
  wire  _EVAL_393;
  wire  _EVAL_394;
  wire  _EVAL_395;
  wire  _EVAL_396;
  wire [31:0] _EVAL_398;
  wire [31:0] _EVAL_400;
  wire [1:0] _EVAL_401;
  wire  _EVAL_402;
  wire  _EVAL_403;
  wire  _EVAL_404;
  wire [31:0] _EVAL_405;
  wire [1:0] _EVAL_406;
  wire  _EVAL_407;
  wire [3:0] _EVAL_408;
  wire  _EVAL_409;
  wire  _EVAL_410;
  wire [32:0] _EVAL_411;
  wire [11:0] _EVAL_412;
  wire [2:0] _EVAL_414;
  wire [13:0] _EVAL_415;
  wire  _EVAL_416;
  wire  _EVAL_417;
  wire  _EVAL_418;
  wire  _EVAL_419;
  wire  _EVAL_420;
  wire  _EVAL_421;
  wire  q__EVAL;
  wire [31:0] q__EVAL_0;
  wire [3:0] q__EVAL_1;
  wire [2:0] q__EVAL_2;
  wire  q__EVAL_3;
  wire [3:0] q__EVAL_4;
  wire  q__EVAL_5;
  wire [31:0] q__EVAL_6;
  wire  q__EVAL_7;
  wire [2:0] q__EVAL_8;
  wire  q__EVAL_9;
  wire  q__EVAL_10;
  wire  q__EVAL_11;
  wire  q__EVAL_12;
  wire  q__EVAL_13;
  wire  q__EVAL_14;
  wire [2:0] q__EVAL_15;
  wire  q__EVAL_16;
  wire [2:0] q__EVAL_17;
  wire  q__EVAL_18;
  wire [31:0] q__EVAL_19;
  wire [3:0] q__EVAL_20;
  wire [2:0] q__EVAL_21;
  wire  q__EVAL_22;
  wire [2:0] q__EVAL_23;
  wire  q__EVAL_24;
  wire [3:0] q__EVAL_25;
  wire [31:0] q__EVAL_26;
  wire  q__EVAL_27;
  wire [31:0] _EVAL_422;
  wire [32:0] _EVAL_423;
  wire  _EVAL_424;
  wire [31:0] _EVAL_425;
  wire [31:0] _EVAL_426;
  wire  _EVAL_427;
  wire  _EVAL_428;
  wire  _EVAL_429;
  wire [11:0] _EVAL_430;
  wire  _EVAL_431;
  wire  _EVAL_433;
  wire  _EVAL_434;
  wire  _EVAL_435;
  wire  _EVAL_437;
  wire  _EVAL_438;
  wire  _EVAL_439;
  wire  _EVAL_440;
  wire [31:0] _EVAL_441;
  wire  _EVAL_442;
  wire [6:0] _EVAL_443;
  wire [6:0] _EVAL_444;
  wire  _EVAL_445;
  wire  _EVAL_446;
  wire  _EVAL_447;
  wire [32:0] _EVAL_448;
  wire  _EVAL_450;
  wire [5:0] _EVAL_451;
  wire [7:0] _EVAL_452;
  wire [3:0] _EVAL_453;
  wire [32:0] _EVAL_454;
  wire [31:0] _EVAL_455;
  wire  _EVAL_456;
  wire [1:0] _EVAL_457;
  wire  _EVAL_458;
  wire [32:0] _EVAL_459;
  wire  _EVAL_460;
  wire [6:0] _EVAL_461;
  wire [1:0] _EVAL_462;
  wire [3:0] _EVAL_463;
  wire [7:0] _EVAL_464;
  wire  _EVAL_466;
  wire [6:0] _EVAL_467;
  wire  _EVAL_468;
  wire  _EVAL_470;
  wire  _EVAL_471;
  wire  _EVAL_472;
  wire [2:0] _EVAL_473;
  wire  _EVAL_475;
  wire [2:0] _EVAL_476;
  wire  _EVAL_477;
  wire [31:0] amoalu__EVAL;
  wire [31:0] amoalu__EVAL_0;
  wire [4:0] amoalu__EVAL_1;
  wire [31:0] amoalu__EVAL_2;
  wire  _EVAL_479;
  wire [7:0] _EVAL_480;
  wire  _EVAL_481;
  wire [13:0] _EVAL_482;
  wire  _EVAL_483;
  wire  _EVAL_484;
  wire [31:0] _EVAL_485;
  wire [1:0] _EVAL_486;
  wire  _EVAL_487;
  wire [2:0] _EVAL_488;
  wire [31:0] _EVAL_489;
  wire  _EVAL_490;
  wire  _EVAL_491;
  wire  _EVAL_492;
  wire [31:0] _EVAL_494;
  wire [31:0] _EVAL_495;
  wire [2:0] _EVAL_496;
  wire [13:0] _EVAL_497;
  wire [2:0] _EVAL_498;
  wire  _EVAL_499;
  wire [1:0] _EVAL_500;
  wire [1:0] _EVAL_501;
  wire  tlb_pmp__EVAL;
  wire [31:0] tlb_pmp__EVAL_0;
  wire [29:0] tlb_pmp__EVAL_1;
  wire  tlb_pmp__EVAL_2;
  wire  tlb_pmp__EVAL_3;
  wire  tlb_pmp__EVAL_4;
  wire [29:0] tlb_pmp__EVAL_5;
  wire  tlb_pmp__EVAL_6;
  wire [1:0] tlb_pmp__EVAL_7;
  wire  tlb_pmp__EVAL_8;
  wire  tlb_pmp__EVAL_9;
  wire [1:0] tlb_pmp__EVAL_10;
  wire [1:0] tlb_pmp__EVAL_11;
  wire [1:0] tlb_pmp__EVAL_12;
  wire  tlb_pmp__EVAL_13;
  wire  tlb_pmp__EVAL_14;
  wire  tlb_pmp__EVAL_15;
  wire [1:0] tlb_pmp__EVAL_16;
  wire  tlb_pmp__EVAL_17;
  wire  tlb_pmp__EVAL_18;
  wire  tlb_pmp__EVAL_19;
  wire [29:0] tlb_pmp__EVAL_20;
  wire  tlb_pmp__EVAL_21;
  wire  tlb_pmp__EVAL_22;
  wire  tlb_pmp__EVAL_23;
  wire [31:0] tlb_pmp__EVAL_24;
  wire  tlb_pmp__EVAL_25;
  wire  tlb_pmp__EVAL_26;
  wire [31:0] tlb_pmp__EVAL_27;
  wire [31:0] tlb_pmp__EVAL_28;
  wire [31:0] tlb_pmp__EVAL_29;
  wire  tlb_pmp__EVAL_30;
  wire [1:0] tlb_pmp__EVAL_31;
  wire [1:0] tlb_pmp__EVAL_32;
  wire [29:0] tlb_pmp__EVAL_33;
  wire [31:0] tlb_pmp__EVAL_34;
  wire  tlb_pmp__EVAL_35;
  wire  tlb_pmp__EVAL_36;
  wire  tlb_pmp__EVAL_37;
  wire [31:0] tlb_pmp__EVAL_38;
  wire [31:0] tlb_pmp__EVAL_39;
  wire [1:0] tlb_pmp__EVAL_40;
  wire [29:0] tlb_pmp__EVAL_41;
  wire [29:0] tlb_pmp__EVAL_42;
  wire  tlb_pmp__EVAL_43;
  wire  tlb_pmp__EVAL_44;
  wire [29:0] tlb_pmp__EVAL_45;
  wire [31:0] tlb_pmp__EVAL_46;
  wire [1:0] tlb_pmp__EVAL_47;
  wire  tlb_pmp__EVAL_48;
  wire  tlb_pmp__EVAL_49;
  wire  tlb_pmp__EVAL_50;
  wire  tlb_pmp__EVAL_51;
  wire  tlb_pmp__EVAL_52;
  wire [29:0] tlb_pmp__EVAL_53;
  wire  tlb_pmp__EVAL_54;
  wire  tlb_pmp__EVAL_55;
  wire  tlb_pmp__EVAL_56;
  wire  tlb_pmp__EVAL_57;
  wire  tlb_pmp__EVAL_58;
  wire  tlb_pmp__EVAL_59;
  wire  tlb_pmp__EVAL_60;
  wire  tlb_pmp__EVAL_61;
  wire  _EVAL_502;
  wire  _EVAL_503;
  wire [31:0] _EVAL_504;
  wire  _EVAL_505;
  wire  _EVAL_506;
  wire [13:0] _EVAL_509;
  wire  _EVAL_510;
  wire  _EVAL_511;
  wire  _EVAL_512;
  wire  _EVAL_513;
  wire  _EVAL_514;
  wire  _EVAL_515;
  wire [2:0] _EVAL_518;
  wire  _EVAL_519;
  wire  _EVAL_520;
  wire  _EVAL_521;
  wire  _EVAL_522;
  wire [1:0] _EVAL_523;
  wire [13:0] _EVAL_524;
  wire  _EVAL_525;
  wire  _EVAL_526;
  wire  _EVAL_528;
  wire [31:0] _EVAL_529;
  wire [2:0] _EVAL_530;
  wire [11:0] _EVAL_531;
  wire  _EVAL_532;
  wire  _EVAL_533;
  wire  _EVAL_535;
  wire [1:0] _EVAL_537;
  wire  _EVAL_538;
  wire  _EVAL_539;
  wire  _EVAL_540;
  wire  _EVAL_542;
  wire  _EVAL_543;
  wire  _EVAL_544;
  wire [13:0] _EVAL_545;
  wire  _EVAL_546;
  wire [2:0] _EVAL_547;
  wire  _EVAL_548;
  wire  _EVAL_549;
  wire  _EVAL_550;
  wire [13:0] _EVAL_551;
  wire [29:0] _EVAL_552;
  wire  _EVAL_555;
  wire [31:0] _EVAL_556;
  wire [32:0] _EVAL_557;
  wire [2:0] _EVAL_558;
  wire [7:0] _EVAL_559;
  wire  _EVAL_560;
  wire [2:0] _EVAL_561;
  wire  _EVAL_562;
  wire [3:0] _EVAL_563;
  wire [29:0] _EVAL_564;
  wire [7:0] _EVAL_565;
  wire [3:0] _EVAL_566;
  wire  _EVAL_567;
  wire  _EVAL_568;
  wire  _EVAL_569;
  wire  _EVAL_570;
  wire  _EVAL_571;
  wire  _EVAL_573;
  wire [13:0] _EVAL_574;
  wire  _EVAL_575;
  wire  _EVAL_576;
  wire [3:0] _EVAL_577;
  wire  _EVAL_578;
  wire [2:0] _EVAL_579;
  wire [2:0] _EVAL_580;
  wire  _EVAL_581;
  wire  _EVAL_582;
  wire  _EVAL_583;
  wire [1:0] _EVAL_584;
  wire [31:0] _EVAL_585;
  wire  _EVAL_586;
  wire  _EVAL_587;
  wire  _EVAL_588;
  wire [3:0] _EVAL_589;
  wire [31:0] _EVAL_590;
  wire [7:0] _EVAL_591;
  wire [7:0] _EVAL_592;
  wire  _EVAL_593;
  wire [13:0] _EVAL_594;
  wire  _EVAL_595;
  wire [1:0] _EVAL_596;
  wire  _EVAL_597;
  wire  _EVAL_599;
  wire  _EVAL_600;
  wire  _EVAL_601;
  wire [13:0] _EVAL_602;
  wire  _EVAL_603;
  wire  _EVAL_604;
  wire  _EVAL_605;
  wire [31:0] _EVAL_606;
  wire [1:0] _EVAL_607;
  wire  _EVAL_608;
  wire [32:0] _EVAL_609;
  wire  _EVAL_610;
  wire  _EVAL_611;
  wire [3:0] _EVAL_612;
  wire [7:0] _EVAL_615;
  wire  _EVAL_616;
  wire [31:0] _EVAL_617;
  wire  _EVAL_618;
  wire [15:0] _EVAL_619;
  wire  _EVAL_620;
  wire  _EVAL_621;
  wire  _EVAL_622;
  wire [5:0] _EVAL_623;
  wire  _EVAL_624;
  wire  _EVAL_625;
  wire  _EVAL_626;
  wire [2:0] _EVAL_627;
  wire [13:0] _EVAL_628;
  wire  _EVAL_629;
  wire  _EVAL_630;
  wire  _EVAL_631;
  wire [32:0] _EVAL_632;
  wire  _EVAL_633;
  wire  _EVAL_634;
  wire  _EVAL_635;
  wire [31:0] _EVAL_636;
  wire  _EVAL_638;
  wire [1:0] _EVAL_639;
  wire  _EVAL_640;
  wire [13:0] _EVAL_641;
  wire  _EVAL_642;
  wire  _EVAL_643;
  wire [13:0] _EVAL_644;
  wire  _EVAL_645;
  wire  _EVAL_646;
  wire [31:0] _EVAL_647;
  wire [7:0] _EVAL_648;
  wire [32:0] _EVAL_649;
  wire [3:0] _EVAL_650;
  wire  _EVAL_651;
  wire  _EVAL_652;
  wire  _EVAL_653;
  wire [3:0] _EVAL_654;
  wire [3:0] _EVAL_655;
  wire  _EVAL_656;
  wire  _EVAL_657;
  wire  _EVAL_658;
  wire [7:0] _EVAL_659;
  wire  _EVAL_661;
  wire  _EVAL_662;
  wire [7:0] _EVAL_663;
  wire  _EVAL_664;
  wire [5:0] _EVAL_665;
  wire  _EVAL_667;
  wire  _EVAL_668;
  wire  _EVAL_669;
  wire  _EVAL_670;
  wire  _EVAL_671;
  wire [6:0] _EVAL_672;
  wire  _EVAL_673;
  wire  _EVAL_674;
  wire [3:0] _EVAL_675;
  wire  _EVAL_677;
  wire  _EVAL_678;
  wire [3:0] _EVAL_679;
  wire [31:0] _EVAL_680;
  wire [3:0] _EVAL_681;
  wire [1:0] _EVAL_682;
  wire  _EVAL_683;
  wire  _EVAL_684;
  wire  _EVAL_685;
  wire  _EVAL_686;
  wire [2:0] _EVAL_687;
  wire [31:0] _EVAL_688;
  wire  _EVAL_689;
  wire  _EVAL_690;
  wire  _EVAL_691;
  wire  _EVAL_693;
  wire  _EVAL_694;
  wire  _EVAL_696;
  wire [32:0] _EVAL_697;
  wire  _EVAL_698;
  wire  _EVAL_699;
  wire  _EVAL_700;
  wire [13:0] _EVAL_701;
  wire  _EVAL_702;
  wire  _EVAL_703;
  wire [31:0] _EVAL_704;
  wire [2:0] _EVAL_706;
  wire  _EVAL_707;
  wire  _EVAL_708;
  wire  _EVAL_709;
  wire [32:0] _EVAL_711;
  wire [3:0] _EVAL_712;
  wire  _EVAL_713;
  wire  _EVAL_714;
  wire  _EVAL_715;
  wire [31:0] _EVAL_716;
  wire [13:0] _EVAL_718;
  wire [1:0] _EVAL_719;
  wire [31:0] _EVAL_720;
  wire  _EVAL_721;
  wire [3:0] _EVAL_722;
  wire  _EVAL_723;
  wire  _EVAL_725;
  wire  _EVAL_726;
  wire [29:0] _EVAL_727;
  wire [22:0] _EVAL_728;
  wire [4:0] _EVAL_729;
  wire  _EVAL_730;
  wire [3:0] _EVAL_731;
  wire [31:0] _EVAL_732;
  wire [3:0] _EVAL_733;
  wire  _EVAL_735;
  wire [29:0] _EVAL_736;
  wire  _EVAL_737;
  wire [3:0] _EVAL_738;
  wire  _EVAL_739;
  wire [31:0] _EVAL_740;
  wire  _EVAL_741;
  wire [31:0] _EVAL_742;
  wire  _EVAL_743;
  wire  _EVAL_745;
  wire  _EVAL_747;
  wire  _EVAL_748;
  wire  _EVAL_749;
  wire  _EVAL_750;
  wire  _EVAL_751;
  wire  _EVAL_752;
  wire [7:0] _EVAL_753;
  wire [3:0] _EVAL_754;
  wire [31:0] _EVAL_756;
  wire  _EVAL_757;
  wire [15:0] _EVAL_758;
  wire  _EVAL_759;
  wire [2:0] _EVAL_760;
  wire  _EVAL_761;
  wire  _EVAL_762;
  wire [1:0] _EVAL_763;
  wire [23:0] _EVAL_764;
  wire  _EVAL_765;
  wire  _EVAL_766;
  wire  _EVAL_767;
  wire  _EVAL_768;
  wire [7:0] _EVAL_769;
  wire  _EVAL_770;
  wire  _EVAL_771;
  wire  _EVAL_772;
  wire  _EVAL_773;
  wire [19:0] _EVAL_774;
  wire  _EVAL_775;
  wire  _EVAL_776;
  wire  _EVAL_777;
  wire [31:0] _EVAL_779;
  wire  _EVAL_780;
  wire  _EVAL_782;
  wire  _EVAL_783;
  wire [2:0] _EVAL_784;
  wire [2:0] _EVAL_785;
  wire [29:0] _EVAL_786;
  wire  _EVAL_787;
  wire  _EVAL_788;
  wire  _EVAL_789;
  wire  _EVAL_791;
  wire [2:0] _EVAL_792;
  wire  _EVAL_793;
  wire  _EVAL_795;
  wire  _EVAL_796;
  wire [2:0] _EVAL_797;
  wire  _EVAL_798;
  wire  _EVAL_799;
  wire [13:0] _EVAL_800;
  wire [3:0] _EVAL_801;
  wire [2:0] _EVAL_802;
  wire  _EVAL_803;
  wire  _EVAL_804;
  wire  _EVAL_805;
  wire  _EVAL_806;
  wire  _EVAL_807;
  wire  _EVAL_808;
  wire [31:0] _EVAL_809;
  wire  _EVAL_810;
  wire  _EVAL_811;
  wire  _EVAL_812;
  wire [1:0] _EVAL_813;
  wire  _EVAL_814;
  wire  _EVAL_815;
  wire  _EVAL_817;
  wire [22:0] _EVAL_818;
  wire [1:0] _EVAL_819;
  wire  _EVAL_820;
  wire [7:0] _EVAL_821;
  wire  _EVAL_822;
  wire  _EVAL_824;
  wire [3:0] _EVAL_825;
  wire [32:0] _EVAL_826;
  wire  _EVAL_827;
  wire  _EVAL_828;
  wire [1:0] _EVAL_829;
  wire [6:0] _EVAL_830;
  wire  _EVAL_831;
  wire  _EVAL_832;
  wire  _EVAL_833;
  wire [13:0] _EVAL_834;
  wire  _EVAL_835;
  wire [7:0] _EVAL_836;
  wire  _EVAL_838;
  wire  _EVAL_840;
  wire [3:0] _EVAL_841;
  wire [31:0] _EVAL_842;
  wire  _EVAL_843;
  wire  _EVAL_844;
  wire  _EVAL_845;
  wire  _EVAL_846;
  wire [31:0] _EVAL_847;
  wire [1:0] _EVAL_848;
  wire  _EVAL_849;
  wire [2:0] _EVAL_850;
  wire [31:0] _EVAL_851;
  wire  _EVAL_852;
  wire  _EVAL_853;
  wire  _EVAL_854;
  wire  _EVAL_855;
  wire  _EVAL_856;
  wire [3:0] _EVAL_858;
  wire [6:0] _EVAL_860;
  wire  _EVAL_861;
  wire [7:0] _EVAL_862;
  wire [3:0] _EVAL_863;
  wire  _EVAL_865;
  wire  _EVAL_866;
  wire [2:0] _EVAL_867;
  wire [23:0] _EVAL_868;
  wire  _EVAL_869;
  wire [31:0] _EVAL_870;
  wire  _EVAL_871;
  wire  _EVAL_872;
  wire  _EVAL_873;
  wire [31:0] _EVAL_874;
  wire  _EVAL_875;
  wire  _EVAL_877;
  wire  _EVAL_878;
  wire  _EVAL_879;
  wire [32:0] _EVAL_880;
  wire  _EVAL_881;
  wire [32:0] _EVAL_882;
  wire [31:0] _EVAL_884;
  wire [6:0] _EVAL_885;
  wire  _EVAL_886;
  wire [13:0] _EVAL_888;
  wire  _EVAL_889;
  wire  _EVAL_890;
  wire  _EVAL_891;
  wire [13:0] _EVAL_892;
  wire [32:0] _EVAL_893;
  wire  _EVAL_894;
  wire [31:0] _EVAL_895;
  wire  _EVAL_896;
  wire  _EVAL_897;
  wire  _EVAL_899;
  wire  _EVAL_900;
  wire  _EVAL_902;
  wire [1:0] _EVAL_903;
  wire [31:0] _EVAL_905;
  wire  _EVAL_906;
  wire [2:0] _EVAL_907;
  wire  _EVAL_909;
  wire [7:0] _EVAL_910;
  wire  _EVAL_912;
  wire  _EVAL_913;
  wire  _EVAL_914;
  wire [1:0] _EVAL_915;
  wire  _EVAL_918;
  wire  _EVAL_919;
  wire  _EVAL_920;
  wire  _EVAL_921;
  wire  _EVAL_922;
  wire [31:0] _EVAL_923;
  wire  _EVAL_924;
  wire  _EVAL_925;
  wire  _EVAL_926;
  wire [2:0] _EVAL_927;
  wire  _EVAL_929;
  wire [31:0] _EVAL_930;
  wire  _EVAL_931;
  wire  _EVAL_932;
  wire  _EVAL_933;
  wire  _EVAL_934;
  wire  _EVAL_935;
  wire  _EVAL_936;
  wire [32:0] _EVAL_937;
  wire [31:0] _EVAL_938;
  wire  lfsr_prng__EVAL;
  wire  lfsr_prng__EVAL_0;
  wire  lfsr_prng__EVAL_1;
  wire  lfsr_prng__EVAL_2;
  wire  lfsr_prng__EVAL_3;
  wire  lfsr_prng__EVAL_4;
  wire  lfsr_prng__EVAL_5;
  wire  lfsr_prng__EVAL_6;
  wire  lfsr_prng__EVAL_7;
  wire  lfsr_prng__EVAL_8;
  wire  lfsr_prng__EVAL_9;
  wire  lfsr_prng__EVAL_10;
  wire  lfsr_prng__EVAL_11;
  wire  lfsr_prng__EVAL_12;
  wire  lfsr_prng__EVAL_13;
  wire  lfsr_prng__EVAL_14;
  wire  lfsr_prng__EVAL_15;
  wire  lfsr_prng__EVAL_16;
  wire  lfsr_prng__EVAL_17;
  wire  _EVAL_940;
  wire [17:0] _EVAL_941;
  wire  _EVAL_942;
  wire [4:0] _EVAL_943;
  wire  _EVAL_945;
  wire  _EVAL_946;
  wire  _EVAL_947;
  wire  _EVAL_949;
  wire [7:0] _EVAL_950;
  wire  _EVAL_951;
  wire [3:0] _EVAL_952;
  wire [32:0] _EVAL_953;
  wire  _EVAL_954;
  wire [2:0] _EVAL_955;
  wire  _EVAL_956;
  wire  _EVAL_957;
  wire [1:0] _EVAL_958;
  wire [31:0] _EVAL_959;
  wire  _EVAL_960;
  wire [29:0] _EVAL_961;
  wire  _EVAL_963;
  wire  _EVAL_964;
  wire  _EVAL_965;
  wire [2:0] _EVAL_966;
  wire  _EVAL_967;
  wire  _EVAL_968;
  wire  _EVAL_969;
  wire  _EVAL_970;
  wire  _EVAL_971;
  wire [25:0] _EVAL_972;
  wire  _EVAL_973;
  wire [1:0] _EVAL_974;
  wire  _EVAL_975;
  wire [31:0] _EVAL_976;
  wire  _EVAL_979;
  wire  _EVAL_980;
  wire  _EVAL_981;
  wire  _EVAL_982;
  wire [1:0] _EVAL_983;
  wire [13:0] _EVAL_984;
  wire  _EVAL_985;
  wire  _EVAL_986;
  wire  _EVAL_987;
  wire [31:0] _EVAL_988;
  wire  _EVAL_989;
  wire  _EVAL_990;
  wire [31:0] _EVAL_991;
  wire  _EVAL_992;
  wire  _EVAL_993;
  wire  _EVAL_995;
  wire [1:0] _EVAL_996;
  wire  _EVAL_998;
  wire  _EVAL_1001;
  wire [31:0] _EVAL_1002;
  wire  _EVAL_1003;
  wire [32:0] _EVAL_1004;
  wire [31:0] _EVAL_1005;
  wire [29:0] _EVAL_1006;
  wire [3:0] _EVAL_1008;
  wire  _EVAL_1009;
  wire [13:0] _EVAL_1010;
  wire  _EVAL_1011;
  wire [1:0] _EVAL_1012;
  wire  _EVAL_1013;
  wire  _EVAL_1015;
  wire [3:0] _EVAL_1016;
  wire [5:0] _EVAL_1017;
  wire  _EVAL_1019;
  wire  _EVAL_1020;
  wire  _EVAL_1021;
  wire [18:0] _EVAL_1022;
  wire  _EVAL_1023;
  wire  _EVAL_1024;
  wire  _EVAL_1025;
  wire  _EVAL_1026;
  wire [1:0] _EVAL_1027;
  wire [6:0] _EVAL_1028;
  wire [32:0] _EVAL_1029;
  wire  _EVAL_1030;
  wire  _EVAL_1032;
  wire  _EVAL_1033;
  wire [1:0] _EVAL_1034;
  wire  _EVAL_1035;
  wire  _EVAL_1037;
  wire  _EVAL_1039;
  wire [31:0] _EVAL_1040;
  wire [13:0] _EVAL_1042;
  wire  _EVAL_1043;
  wire [3:0] _EVAL_1044;
  wire [1:0] _EVAL_1045;
  wire [13:0] _EVAL_1046;
  wire [6:0] _EVAL_1047;
  wire [31:0] _EVAL_1048;
  wire  _EVAL_1049;
  wire  _EVAL_1050;
  wire [31:0] _EVAL_1051;
  wire  _EVAL_1053;
  wire [31:0] _EVAL_1054;
  wire [13:0] _EVAL_1055;
  wire  _EVAL_1056;
  wire  _EVAL_1057;
  wire [32:0] _EVAL_1059;
  wire [6:0] _EVAL_1060;
  wire [17:0] _EVAL_1061;
  wire  _EVAL_1062;
  wire  _EVAL_1064;
  wire [7:0] _EVAL_1065;
  wire  _EVAL_1066;
  wire [31:0] _EVAL_1067;
  wire [31:0] _EVAL_1068;
  wire [1:0] _EVAL_1069;
  wire [17:0] _EVAL_1070;
  wire  _EVAL_1071;
  wire [1:0] _EVAL_1072;
  wire  _EVAL_1073;
  wire  _EVAL_1075;
  wire  _EVAL_1077;
  wire [31:0] _EVAL_1078;
  wire  _EVAL_1079;
  wire [15:0] _EVAL_1081;
  wire [31:0] _EVAL_1082;
  wire  _EVAL_1083;
  wire  _EVAL_1084;
  wire [2:0] _EVAL_1085;
  wire [31:0] _EVAL_1086;
  wire  _EVAL_1087;
  wire  _EVAL_1088;
  wire  _EVAL_1089;
  wire [31:0] _EVAL_1090;
  wire [32:0] _EVAL_1091;
  wire [31:0] _EVAL_1092;
  wire [13:0] _EVAL_1093;
  wire  _EVAL_1094;
  wire [15:0] _EVAL_1096;
  wire  _EVAL_1097;
  wire [1:0] _EVAL_1098;
  wire [31:0] _EVAL_1100;
  wire  _EVAL_1101;
  wire [4:0] _EVAL_1102;
  wire [13:0] _EVAL_1103;
  wire  _EVAL_1104;
  wire  _EVAL_1105;
  wire [2:0] _EVAL_1106;
  wire  _EVAL_1107;
  wire [31:0] _EVAL_1108;
  wire  _EVAL_1109;
  wire  _EVAL_1110;
  wire [7:0] _EVAL_1111;
  wire  _EVAL_1112;
  wire  _EVAL_1113;
  wire [13:0] _EVAL_1114;
  wire  _EVAL_1115;
  wire  _EVAL_1116;
  wire  _EVAL_1117;
  wire  _EVAL_1118;
  wire  _EVAL_1119;
  wire  _EVAL_1120;
  wire [32:0] _EVAL_1121;
  wire [32:0] _EVAL_1122;
  wire  _EVAL_1123;
  wire [13:0] _EVAL_1124;
  wire [11:0] _EVAL_1125;
  wire  _EVAL_1126;
  wire  _EVAL_1127;
  wire [3:0] _EVAL_1129;
  wire  _EVAL_1130;
  wire [1:0] _EVAL_1131;
  wire  _EVAL_1132;
  wire  _EVAL_1133;
  wire [3:0] _EVAL_1134;
  wire  _EVAL_1137;
  wire  _EVAL_1138;
  wire [7:0] _EVAL_1139;
  wire  _EVAL_1140;
  wire  _EVAL_1142;
  wire [2:0] _EVAL_1143;
  wire [31:0] _EVAL_1144;
  wire [23:0] _EVAL_1145;
  wire  _EVAL_1146;
  wire  _EVAL_1147;
  wire  _EVAL_1149;
  wire  _EVAL_1150;
  wire [3:0] _EVAL_1151;
  wire  _EVAL_1152;
  wire [31:0] _EVAL_1154;
  wire  _EVAL_1155;
  wire  _EVAL_1156;
  wire  _EVAL_1157;
  wire [31:0] _EVAL_1159;
  reg  _EVAL_1160;
  wire  _EVAL_1161;
  wire [32:0] _EVAL_1163;
  wire  _EVAL_1164;
  wire  _EVAL_1165;
  wire  _EVAL_1166;
  wire  _EVAL_1167;
  wire [32:0] _EVAL_1169;
  wire [1:0] _EVAL_1170;
  wire [6:0] _EVAL_1171;
  wire  _EVAL_1172;
  wire  _EVAL_1173;
  wire [6:0] _EVAL_1174;
  wire  _EVAL_1175;
  wire  _EVAL_1176;
  wire  _EVAL_1178;
  wire  _EVAL_1180;
  wire  _EVAL_1181;
  wire [19:0] _EVAL_1182;
  wire  _EVAL_1183;
  wire  _EVAL_1184;
  wire  _EVAL_1185;
  wire  _EVAL_1186;
  wire  _EVAL_1187;
  wire  _EVAL_1188;
  wire [32:0] _EVAL_1189;
  wire [31:0] _EVAL_1190;
  wire  _EVAL_1191;
  wire  _EVAL_1192;
  wire  _EVAL_1193;
  wire [6:0] _EVAL_1196;
  wire [13:0] _EVAL_1197;
  wire  _EVAL_1198;
  wire [1:0] _EVAL_1199;
  wire [32:0] _EVAL_1200;
  wire  _EVAL_1201;
  wire  _EVAL_1202;
  wire [1:0] _EVAL_1204;
  wire  _EVAL_1205;
  wire  _EVAL_1206;
  wire [31:0] _EVAL_1207;
  wire  _EVAL_1208;
  wire  _EVAL_1210;
  wire  _EVAL_1211;
  wire  _EVAL_1212;
  wire  _EVAL_1214;
  wire  _EVAL_1215;
  wire [32:0] _EVAL_1216;
  wire  _EVAL_1217;
  wire [7:0] _EVAL_1218;
  wire  _EVAL_1219;
  wire [1:0] _EVAL_1220;
  wire [3:0] _EVAL_1221;
  wire [2:0] _EVAL_1222;
  wire  _EVAL_1223;
  wire [32:0] _EVAL_1224;
  wire  _EVAL_1225;
  wire  _EVAL_1226;
  wire [2:0] _EVAL_1227;
  wire  _EVAL_1228;
  wire  _EVAL_1229;
  wire [1:0] _EVAL_1230;
  wire [1:0] _EVAL_1231;
  wire [31:0] _EVAL_1232;
  wire  _EVAL_1233;
  wire  _EVAL_1234;
  wire  _EVAL_1235;
  wire [2:0] _EVAL_1236;
  wire [7:0] _EVAL_1237;
  wire [31:0] _EVAL_1238;
  wire  _EVAL_1239;
  wire  _EVAL_1240;
  wire [13:0] _EVAL_1241;
  wire  _EVAL_1242;
  wire  _EVAL_1243;
  wire [3:0] _EVAL_1244;
  wire [32:0] _EVAL_1245;
  wire  _EVAL_1246;
  wire  _EVAL_1247;
  wire  _EVAL_1248;
  wire [6:0] _EVAL_1249;
  wire [1:0] _EVAL_1250;
  wire  _EVAL_1251;
  wire [1:0] _EVAL_1252;
  wire  _EVAL_1253;
  wire [6:0] _EVAL_1254;
  wire  _EVAL_1255;
  wire  _EVAL_1256;
  wire [3:0] _EVAL_1259;
  wire  _EVAL_1260;
  wire [1:0] _EVAL_1261;
  wire  gated_clock_dcache_clock_gate_in;
  wire  gated_clock_dcache_clock_gate_test_en;
  wire  gated_clock_dcache_clock_gate_en;
  wire  gated_clock_dcache_clock_gate_out;
  reg [1:0] _EVAL_1263;
  reg  _EVAL_1264;
  reg  _EVAL_1265;
  reg  _EVAL_1266;
  reg  _EVAL_1267;
  reg [6:0] _EVAL_1268;
  reg [31:0] _EVAL_1269;
  reg  _EVAL_1270;
  reg [31:0] _EVAL_1271;
  reg  _EVAL_1272;
  reg [5:0] _EVAL_1273;
  reg [31:0] _EVAL_1274;
  reg [1:0] _EVAL_1275;
  reg [31:0] _EVAL_1276;
  reg  _EVAL_1277;
  reg [4:0] _EVAL_1278;
  reg [6:0] _EVAL_1279;
  reg  _EVAL_1280;
  reg [1:0] _EVAL_1281;
  reg  _EVAL_1282;
  reg [1:0] _EVAL_1283;
  reg [3:0] _EVAL_1284;
  reg  _EVAL_1285;
  reg [31:0] _EVAL_1286;
  reg [4:0] _EVAL_1287;
  reg [1:0] _EVAL_1288;
  reg  _EVAL_1289;
  reg [1:0] _EVAL_1290;
  reg [7:0] _EVAL_1291;
  reg [4:0] _EVAL_1292;
  reg  _EVAL_1293;
  reg  _EVAL_1294;
  reg [31:0] _EVAL_1295;
  reg [5:0] _EVAL_1296;
  reg [31:0] _EVAL_1297;
  reg [1:0] _EVAL_1298;
  reg  _EVAL_1299;
  reg  _EVAL_1300;
  reg [6:0] _EVAL_1301;
  reg [1:0] _EVAL_1302;
  reg  _EVAL_1303;
  reg [7:0] _EVAL_1304;
  reg [7:0] _EVAL_1305;
  reg [3:0] _EVAL_1306;
  reg  _EVAL_1307;
  reg [31:0] _EVAL_1308;
  reg [6:0] _EVAL_1309;
  reg [1:0] _EVAL_1310;
  reg [31:0] _EVAL_1311;
  reg [31:0] _EVAL_1312;
  reg [6:0] _EVAL_1313;
  reg [6:0] _EVAL_1314;
  reg [1:0] _EVAL_1315;
  reg [31:0] _EVAL_1316;
  reg [1:0] _EVAL_1317;
  reg  _EVAL_1318;
  reg  _EVAL_1319;
  reg  _EVAL_1320;
  reg [6:0] _EVAL_1321;
  reg [31:0] _EVAL_1322;
  reg [6:0] _EVAL_1323;
  reg  _EVAL_1324;
  reg [6:0] _EVAL_1325;
  reg [1:0] _EVAL_1326;
  reg  _EVAL_1327;
  reg  _EVAL_1328;
  reg [31:0] _EVAL_1329;
  reg  _EVAL_1330;
  reg [31:0] _EVAL_1331;
  reg  _EVAL_1332;
  reg  _EVAL_1333;
  reg  _EVAL_1334;
  reg [7:0] _EVAL_1335;
  reg [3:0] _EVAL_1336;
  reg  _EVAL_1337;
  reg  _EVAL_1338;
  reg  _EVAL_1339;
  reg  _EVAL_1340;
  reg [6:0] _EVAL_1341;
  reg  _EVAL_1342;
  reg [31:0] _EVAL_1343;
  reg [1:0] _EVAL_1344;
  reg [3:0] _EVAL_1345;
  reg [2:0] _EVAL_1346;
  reg  _EVAL_1347;
  reg  _EVAL_1348;
  reg [31:0] _EVAL_1349;
  reg  _EVAL_1350;
  reg [4:0] _EVAL_1351;
  wire  _EVAL_1352;
  wire [3:0] _EVAL_1353;
  wire [7:0] _EVAL_1354;
  wire  _EVAL_1355;
  wire [5:0] _EVAL_1356;
  wire [3:0] _EVAL_1357;
  wire [31:0] _EVAL_1359;
  wire  _EVAL_1360;
  wire [1:0] _EVAL_1361;
  wire [1:0] _EVAL_1362;
  wire [32:0] _EVAL_1363;
  wire  _EVAL_1364;
  wire [7:0] _EVAL_1365;
  wire [31:0] _EVAL_1366;
  wire  _EVAL_1367;
  wire  _EVAL_1368;
  wire [32:0] _EVAL_1369;
  wire  _EVAL_1370;
  wire [13:0] _EVAL_1371;
  wire  _EVAL_1372;
  wire [3:0] _EVAL_1373;
  wire  _EVAL_1374;
  wire  _EVAL_1375;
  wire  _EVAL_1376;
  wire [32:0] _EVAL_1377;
  wire [15:0] _EVAL_1378;
  wire  _EVAL_1379;
  wire  _EVAL_1380;
  wire  _EVAL_1382;
  wire  _EVAL_1383;
  wire  _EVAL_1384;
  wire  _EVAL_1385;
  wire [7:0] _EVAL_1386;
  wire [2:0] _EVAL_1387;
  wire  _EVAL_1388;
  wire  _EVAL_1389;
  _EVAL_105 pma_checker_pmp (
    ._EVAL(pma_checker_pmp__EVAL),
    ._EVAL_0(pma_checker_pmp__EVAL_0),
    ._EVAL_1(pma_checker_pmp__EVAL_1),
    ._EVAL_2(pma_checker_pmp__EVAL_2),
    ._EVAL_3(pma_checker_pmp__EVAL_3),
    ._EVAL_4(pma_checker_pmp__EVAL_4),
    ._EVAL_5(pma_checker_pmp__EVAL_5),
    ._EVAL_6(pma_checker_pmp__EVAL_6),
    ._EVAL_7(pma_checker_pmp__EVAL_7),
    ._EVAL_8(pma_checker_pmp__EVAL_8),
    ._EVAL_9(pma_checker_pmp__EVAL_9),
    ._EVAL_10(pma_checker_pmp__EVAL_10),
    ._EVAL_11(pma_checker_pmp__EVAL_11),
    ._EVAL_12(pma_checker_pmp__EVAL_12),
    ._EVAL_13(pma_checker_pmp__EVAL_13),
    ._EVAL_14(pma_checker_pmp__EVAL_14),
    ._EVAL_15(pma_checker_pmp__EVAL_15),
    ._EVAL_16(pma_checker_pmp__EVAL_16),
    ._EVAL_17(pma_checker_pmp__EVAL_17),
    ._EVAL_18(pma_checker_pmp__EVAL_18),
    ._EVAL_19(pma_checker_pmp__EVAL_19),
    ._EVAL_20(pma_checker_pmp__EVAL_20),
    ._EVAL_21(pma_checker_pmp__EVAL_21),
    ._EVAL_22(pma_checker_pmp__EVAL_22),
    ._EVAL_23(pma_checker_pmp__EVAL_23),
    ._EVAL_24(pma_checker_pmp__EVAL_24),
    ._EVAL_25(pma_checker_pmp__EVAL_25),
    ._EVAL_26(pma_checker_pmp__EVAL_26),
    ._EVAL_27(pma_checker_pmp__EVAL_27),
    ._EVAL_28(pma_checker_pmp__EVAL_28),
    ._EVAL_29(pma_checker_pmp__EVAL_29),
    ._EVAL_30(pma_checker_pmp__EVAL_30),
    ._EVAL_31(pma_checker_pmp__EVAL_31),
    ._EVAL_32(pma_checker_pmp__EVAL_32),
    ._EVAL_33(pma_checker_pmp__EVAL_33),
    ._EVAL_34(pma_checker_pmp__EVAL_34),
    ._EVAL_35(pma_checker_pmp__EVAL_35),
    ._EVAL_36(pma_checker_pmp__EVAL_36),
    ._EVAL_37(pma_checker_pmp__EVAL_37),
    ._EVAL_38(pma_checker_pmp__EVAL_38),
    ._EVAL_39(pma_checker_pmp__EVAL_39),
    ._EVAL_40(pma_checker_pmp__EVAL_40),
    ._EVAL_41(pma_checker_pmp__EVAL_41),
    ._EVAL_42(pma_checker_pmp__EVAL_42),
    ._EVAL_43(pma_checker_pmp__EVAL_43),
    ._EVAL_44(pma_checker_pmp__EVAL_44),
    ._EVAL_45(pma_checker_pmp__EVAL_45),
    ._EVAL_46(pma_checker_pmp__EVAL_46),
    ._EVAL_47(pma_checker_pmp__EVAL_47),
    ._EVAL_48(pma_checker_pmp__EVAL_48),
    ._EVAL_49(pma_checker_pmp__EVAL_49),
    ._EVAL_50(pma_checker_pmp__EVAL_50),
    ._EVAL_51(pma_checker_pmp__EVAL_51),
    ._EVAL_52(pma_checker_pmp__EVAL_52),
    ._EVAL_53(pma_checker_pmp__EVAL_53),
    ._EVAL_54(pma_checker_pmp__EVAL_54),
    ._EVAL_55(pma_checker_pmp__EVAL_55),
    ._EVAL_56(pma_checker_pmp__EVAL_56),
    ._EVAL_57(pma_checker_pmp__EVAL_57),
    ._EVAL_58(pma_checker_pmp__EVAL_58),
    ._EVAL_59(pma_checker_pmp__EVAL_59),
    ._EVAL_60(pma_checker_pmp__EVAL_60),
    ._EVAL_61(pma_checker_pmp__EVAL_61)
  );
  _EVAL_107 data (
    ._EVAL(data__EVAL),
    ._EVAL_0(data__EVAL_0),
    ._EVAL_1(data__EVAL_1),
    ._EVAL_2(data__EVAL_2),
    ._EVAL_3(data__EVAL_3),
    ._EVAL_4(data__EVAL_4),
    ._EVAL_5(data__EVAL_5)
  );
  _EVAL_108 q (
    ._EVAL(q__EVAL),
    ._EVAL_0(q__EVAL_0),
    ._EVAL_1(q__EVAL_1),
    ._EVAL_2(q__EVAL_2),
    ._EVAL_3(q__EVAL_3),
    ._EVAL_4(q__EVAL_4),
    ._EVAL_5(q__EVAL_5),
    ._EVAL_6(q__EVAL_6),
    ._EVAL_7(q__EVAL_7),
    ._EVAL_8(q__EVAL_8),
    ._EVAL_9(q__EVAL_9),
    ._EVAL_10(q__EVAL_10),
    ._EVAL_11(q__EVAL_11),
    ._EVAL_12(q__EVAL_12),
    ._EVAL_13(q__EVAL_13),
    ._EVAL_14(q__EVAL_14),
    ._EVAL_15(q__EVAL_15),
    ._EVAL_16(q__EVAL_16),
    ._EVAL_17(q__EVAL_17),
    ._EVAL_18(q__EVAL_18),
    ._EVAL_19(q__EVAL_19),
    ._EVAL_20(q__EVAL_20),
    ._EVAL_21(q__EVAL_21),
    ._EVAL_22(q__EVAL_22),
    ._EVAL_23(q__EVAL_23),
    ._EVAL_24(q__EVAL_24),
    ._EVAL_25(q__EVAL_25),
    ._EVAL_26(q__EVAL_26),
    ._EVAL_27(q__EVAL_27)
  );
  _EVAL_109 amoalu (
    ._EVAL(amoalu__EVAL),
    ._EVAL_0(amoalu__EVAL_0),
    ._EVAL_1(amoalu__EVAL_1),
    ._EVAL_2(amoalu__EVAL_2)
  );
  _EVAL_105 tlb_pmp (
    ._EVAL(tlb_pmp__EVAL),
    ._EVAL_0(tlb_pmp__EVAL_0),
    ._EVAL_1(tlb_pmp__EVAL_1),
    ._EVAL_2(tlb_pmp__EVAL_2),
    ._EVAL_3(tlb_pmp__EVAL_3),
    ._EVAL_4(tlb_pmp__EVAL_4),
    ._EVAL_5(tlb_pmp__EVAL_5),
    ._EVAL_6(tlb_pmp__EVAL_6),
    ._EVAL_7(tlb_pmp__EVAL_7),
    ._EVAL_8(tlb_pmp__EVAL_8),
    ._EVAL_9(tlb_pmp__EVAL_9),
    ._EVAL_10(tlb_pmp__EVAL_10),
    ._EVAL_11(tlb_pmp__EVAL_11),
    ._EVAL_12(tlb_pmp__EVAL_12),
    ._EVAL_13(tlb_pmp__EVAL_13),
    ._EVAL_14(tlb_pmp__EVAL_14),
    ._EVAL_15(tlb_pmp__EVAL_15),
    ._EVAL_16(tlb_pmp__EVAL_16),
    ._EVAL_17(tlb_pmp__EVAL_17),
    ._EVAL_18(tlb_pmp__EVAL_18),
    ._EVAL_19(tlb_pmp__EVAL_19),
    ._EVAL_20(tlb_pmp__EVAL_20),
    ._EVAL_21(tlb_pmp__EVAL_21),
    ._EVAL_22(tlb_pmp__EVAL_22),
    ._EVAL_23(tlb_pmp__EVAL_23),
    ._EVAL_24(tlb_pmp__EVAL_24),
    ._EVAL_25(tlb_pmp__EVAL_25),
    ._EVAL_26(tlb_pmp__EVAL_26),
    ._EVAL_27(tlb_pmp__EVAL_27),
    ._EVAL_28(tlb_pmp__EVAL_28),
    ._EVAL_29(tlb_pmp__EVAL_29),
    ._EVAL_30(tlb_pmp__EVAL_30),
    ._EVAL_31(tlb_pmp__EVAL_31),
    ._EVAL_32(tlb_pmp__EVAL_32),
    ._EVAL_33(tlb_pmp__EVAL_33),
    ._EVAL_34(tlb_pmp__EVAL_34),
    ._EVAL_35(tlb_pmp__EVAL_35),
    ._EVAL_36(tlb_pmp__EVAL_36),
    ._EVAL_37(tlb_pmp__EVAL_37),
    ._EVAL_38(tlb_pmp__EVAL_38),
    ._EVAL_39(tlb_pmp__EVAL_39),
    ._EVAL_40(tlb_pmp__EVAL_40),
    ._EVAL_41(tlb_pmp__EVAL_41),
    ._EVAL_42(tlb_pmp__EVAL_42),
    ._EVAL_43(tlb_pmp__EVAL_43),
    ._EVAL_44(tlb_pmp__EVAL_44),
    ._EVAL_45(tlb_pmp__EVAL_45),
    ._EVAL_46(tlb_pmp__EVAL_46),
    ._EVAL_47(tlb_pmp__EVAL_47),
    ._EVAL_48(tlb_pmp__EVAL_48),
    ._EVAL_49(tlb_pmp__EVAL_49),
    ._EVAL_50(tlb_pmp__EVAL_50),
    ._EVAL_51(tlb_pmp__EVAL_51),
    ._EVAL_52(tlb_pmp__EVAL_52),
    ._EVAL_53(tlb_pmp__EVAL_53),
    ._EVAL_54(tlb_pmp__EVAL_54),
    ._EVAL_55(tlb_pmp__EVAL_55),
    ._EVAL_56(tlb_pmp__EVAL_56),
    ._EVAL_57(tlb_pmp__EVAL_57),
    ._EVAL_58(tlb_pmp__EVAL_58),
    ._EVAL_59(tlb_pmp__EVAL_59),
    ._EVAL_60(tlb_pmp__EVAL_60),
    ._EVAL_61(tlb_pmp__EVAL_61)
  );
  _EVAL_106 lfsr_prng (
    ._EVAL(lfsr_prng__EVAL),
    ._EVAL_0(lfsr_prng__EVAL_0),
    ._EVAL_1(lfsr_prng__EVAL_1),
    ._EVAL_2(lfsr_prng__EVAL_2),
    ._EVAL_3(lfsr_prng__EVAL_3),
    ._EVAL_4(lfsr_prng__EVAL_4),
    ._EVAL_5(lfsr_prng__EVAL_5),
    ._EVAL_6(lfsr_prng__EVAL_6),
    ._EVAL_7(lfsr_prng__EVAL_7),
    ._EVAL_8(lfsr_prng__EVAL_8),
    ._EVAL_9(lfsr_prng__EVAL_9),
    ._EVAL_10(lfsr_prng__EVAL_10),
    ._EVAL_11(lfsr_prng__EVAL_11),
    ._EVAL_12(lfsr_prng__EVAL_12),
    ._EVAL_13(lfsr_prng__EVAL_13),
    ._EVAL_14(lfsr_prng__EVAL_14),
    ._EVAL_15(lfsr_prng__EVAL_15),
    ._EVAL_16(lfsr_prng__EVAL_16),
    ._EVAL_17(lfsr_prng__EVAL_17)
  );
  EICG_wrapper gated_clock_dcache_clock_gate (
    .in(gated_clock_dcache_clock_gate_in),
    .test_en(gated_clock_dcache_clock_gate_test_en),
    .en(gated_clock_dcache_clock_gate_en),
    .out(gated_clock_dcache_clock_gate_out)
  );
  assign _EVAL_650 = _EVAL_513 ? _EVAL_323 : _EVAL_1357;
  assign _EVAL_203 = _EVAL_1164 | _EVAL_1167;
  assign _EVAL_543 = ~_EVAL_1152;
  assign _EVAL_524 = _EVAL_1239 ? _EVAL_1093 : 14'h0;
  assign lfsr_prng__EVAL_2 = _EVAL_776 & _EVAL_548;
  assign _EVAL_699 = _EVAL_492 ? 1'h0 : _EVAL_439;
  assign _EVAL_1072 = _EVAL_1220 | _EVAL_584;
  assign q__EVAL_26 = _EVAL_153 ? _EVAL_1329 : _EVAL_361;
  assign _EVAL_395 = _EVAL_1317[0];
  assign _EVAL_936 = _EVAL_1047[1];
  assign _EVAL_1069 = _EVAL_1072 | _EVAL_275;
  assign _EVAL_607 = _EVAL_60;
  assign tlb_pmp__EVAL_43 = _EVAL_625;
  assign _EVAL_31 = _EVAL_1265;
  assign _EVAL_289 = _EVAL_1247 ? _EVAL_1387 : _EVAL_760;
  assign _EVAL_642 = _EVAL_287 | _EVAL_1319;
  assign _EVAL_851 = _EVAL_606 ^ 32'h40000000;
  assign _EVAL_138 = _EVAL_1016[1];
  assign _EVAL_328 = ~_EVAL_196;
  assign _EVAL_934 = _EVAL_217 & _EVAL_445;
  assign _EVAL_133 = {_EVAL_1350,_EVAL_1330,_EVAL_1272,_EVAL_1303,_EVAL_1342,_EVAL_1318,_EVAL_1307};
  assign _EVAL_129 = _EVAL_48;
  assign data__EVAL = _EVAL_1212;
  assign _EVAL_1180 = _EVAL_1317 >= 2'h2;
  assign _EVAL_230 = _EVAL_278 ? 1'h0 : 1'h1;
  assign _EVAL_1171 = _EVAL_470 ? 7'h4f : 7'h0;
  assign _EVAL_663 = _EVAL_1112 ? 8'hff : 8'h0;
  assign _EVAL_836 = _EVAL_1308[23:16];
  assign _EVAL_748 = _EVAL_1333 & _EVAL_207;
  assign _EVAL_248 = {_EVAL_1354,_EVAL_659};
  assign _EVAL_691 = _EVAL_1302 == 2'h1;
  assign _EVAL_983 = _EVAL_526 ? _EVAL_1131 : 2'h0;
  assign _EVAL_1071 = _EVAL_492 & _EVAL_631;
  assign _EVAL_1091 = $signed(_EVAL_208) & -33'sh1000;
  assign _EVAL_946 = _EVAL_1188 & _EVAL_1256;
  assign _EVAL_460 = _EVAL_540 ? 1'h0 : _EVAL_284;
  assign _EVAL_698 = _EVAL_861 | _EVAL_709;
  assign _EVAL_406 = _EVAL_1069 | _EVAL_996;
  assign pma_checker_pmp__EVAL_18 = 1'h0;
  assign _EVAL_1261 = _EVAL_651 ? _EVAL_1317 : _EVAL_1302;
  assign _EVAL_1384 = _EVAL_1351 == 5'h4;
  assign _EVAL_627 = _EVAL_35;
  assign pma_checker_pmp__EVAL_6 = 1'h0;
  assign _EVAL_988 = _EVAL_606 ^ 32'h80000000;
  assign _EVAL_813 = _EVAL_608 ? 2'h3 : 2'h0;
  assign _EVAL_843 = _EVAL_771 | _EVAL_152;
  assign _EVAL_265 = _EVAL_1298 == _EVAL_457;
  assign _EVAL_153 = ~_EVAL_316;
  assign pma_checker_pmp__EVAL_10 = 2'h0;
  assign _EVAL_701 = _EVAL_641 & 14'h2000;
  assign _EVAL_725 = _EVAL_1110 & _EVAL_316;
  assign _EVAL_1256 = _EVAL_1285 | _EVAL_1347;
  assign tlb_pmp__EVAL_39 = _EVAL_809;
  assign _EVAL_812 = ~_EVAL_730;
  assign _EVAL_1386 = _EVAL_556[23:16];
  assign _EVAL_1371 = _EVAL_294 & 14'h2000;
  assign pma_checker_pmp__EVAL_30 = _EVAL_1214;
  assign _EVAL_1152 = _EVAL_32 & _EVAL_338;
  assign tlb_pmp__EVAL_58 = _EVAL_1146;
  assign tlb_pmp__EVAL_45 = _EVAL_1006;
  assign _EVAL_570 = _EVAL_435 | _EVAL_169;
  assign _EVAL_1089 = _EVAL_651 ? _EVAL_1300 : _EVAL_1265;
  assign _EVAL_1040 = q__EVAL_19;
  assign _EVAL_589 = q__EVAL_20;
  assign _EVAL_722 = {_EVAL_575,_EVAL_490,_EVAL_838,_EVAL_745};
  assign _EVAL_128 = _EVAL_1267 & _EVAL_1334;
  assign _EVAL_514 = _EVAL_1302 == 2'h0;
  assign _EVAL_278 = _EVAL_1271[0];
  assign tlb_pmp__EVAL_36 = _EVAL_1104;
  assign _EVAL_272 = _EVAL_135 | _EVAL_1043;
  assign _EVAL_1020 = _EVAL_216 & _EVAL_1073;
  assign _EVAL_131 = _EVAL_245 | _EVAL_992;
  assign _EVAL_912 = _EVAL_520 | _EVAL_652;
  assign _EVAL_856 = ~_EVAL_291;
  assign _EVAL_425 = {_EVAL_774,_EVAL_430};
  assign _EVAL_1118 = _EVAL_68;
  assign _EVAL_511 = _EVAL_1217 ? _EVAL_232 : _EVAL_1350;
  assign _EVAL_1029 = $signed(_EVAL_352) & -33'sh2000;
  assign amoalu__EVAL_0 = {_EVAL_344,_EVAL_1096};
  assign _EVAL_198 = _EVAL_70 & _EVAL_32;
  assign _EVAL_33 = _EVAL_1110 | _EVAL_1328;
  assign _EVAL_914 = ~_EVAL_920;
  assign _EVAL_160 = _EVAL_766 ? 3'h1 : _EVAL_277;
  assign _EVAL_581 = _EVAL_1278 == 5'h8;
  assign _EVAL_127 = _EVAL_1143;
  assign _EVAL_189 = _EVAL_1013 ? _EVAL_1309 : 7'h0;
  assign _EVAL_617 = _EVAL_959 | _EVAL_842;
  assign _EVAL_974 = _EVAL_180 ? 2'h3 : _EVAL_145;
  assign _EVAL_304 = _EVAL_201 ? _EVAL_1329 : _EVAL_1159;
  assign tlb_pmp__EVAL_20 = _EVAL_736;
  assign _EVAL_585 = _EVAL_914 ? _EVAL_1331 : _EVAL_161;
  assign pma_checker_pmp__EVAL_38 = 32'h0;
  assign _EVAL_229 = _EVAL_648[6:0];
  assign pma_checker_pmp__EVAL_24 = 32'h0;
  assign _EVAL_743 = _EVAL_488[0];
  assign _EVAL_1234 = _EVAL_902 | _EVAL_750;
  assign _EVAL_892 = _EVAL_256 & 14'h2000;
  assign _EVAL_913 = _EVAL_943 == 5'h4;
  assign _EVAL_1239 = _EVAL_900 | _EVAL_499;
  assign _EVAL_670 = q__EVAL_9;
  assign _EVAL_155 = _EVAL_1254[5:0];
  assign _EVAL_143 = _EVAL_23;
  assign _EVAL_952 = _EVAL_1333 ? _EVAL_1284 : _EVAL_1306;
  assign _EVAL_801 = _EVAL_1037 ? _EVAL_731 : _EVAL_612;
  assign _EVAL_351 = 4'h2 == _EVAL_733;
  assign _EVAL_866 = _EVAL_1298 > 2'h0;
  assign _EVAL_168 = _EVAL_1271[13:0];
  assign _EVAL_949 = _EVAL_952[1];
  assign _EVAL_1205 = _EVAL_173 | _EVAL_799;
  assign _EVAL_593 = _EVAL_780 & _EVAL_539;
  assign _EVAL_485 = _EVAL_494;
  assign _EVAL_386 = _EVAL_751 & _EVAL_1385;
  assign _EVAL_441 = _EVAL_156 ? _EVAL_1349 : 32'h0;
  assign q__EVAL_24 = gated_clock_dcache_clock_gate_out;
  assign gated_clock_dcache_clock_gate_in = _EVAL_112;
  assign _EVAL_385 = _EVAL_1067[31:24];
  assign _EVAL_1073 = _EVAL_1181 & _EVAL_1132;
  assign _EVAL_675 = _EVAL_655 & _EVAL_378;
  assign _EVAL_423 = $signed(_EVAL_208) & 33'shcb002000;
  assign _EVAL_107 = _EVAL_1302;
  assign _EVAL_1353 = _EVAL_1248 ? _EVAL_1129 : 4'hf;
  assign _EVAL_255 = _EVAL_1372 ? 1'h0 : _EVAL_460;
  assign _EVAL_772 = _EVAL_492 | _EVAL_1071;
  assign _EVAL_900 = _EVAL_1130 | _EVAL_1084;
  assign _EVAL_86 = _EVAL_1267 & _EVAL_1327;
  assign _EVAL_881 = _EVAL_943 == 5'h1;
  assign _EVAL_1163 = _EVAL_157;
  assign _EVAL_1186 = ~_EVAL_1116;
  assign gated_clock_dcache_clock_gate_test_en = _EVAL_19;
  assign tlb_pmp__EVAL_14 = _EVAL_224;
  assign _EVAL_1147 = $signed(_EVAL_632) == 33'sh0;
  assign _EVAL_945 = _EVAL_1284[2];
  assign _EVAL_1090 = {_EVAL_385,_EVAL_910,_EVAL_559,_EVAL_565};
  assign _EVAL_623 = {_EVAL_27,_EVAL_86,_EVAL_50,_EVAL_11,_EVAL_34,_EVAL_128};
  assign _EVAL_197 = _EVAL_1351 == 5'h7;
  assign _EVAL_764 = _EVAL_814 ? 24'hffffff : 24'h0;
  assign _EVAL_807 = _EVAL_1283 == 2'h1;
  assign _EVAL_500 = {_EVAL_515,_EVAL_137};
  assign _EVAL_1192 = _EVAL_98 == 5'hb;
  assign _EVAL_228 = _EVAL_1308[15:8];
  assign _EVAL_825 = _EVAL_956 ? _EVAL_1134 : _EVAL_1353;
  assign _EVAL_1054 = {_EVAL_1061,_EVAL_415};
  assign _EVAL_472 = _EVAL_98 == 5'h8;
  assign tlb_pmp__EVAL_47 = _EVAL_473[1:0];
  assign _EVAL_921 = _EVAL_266 & _EVAL_1293;
  assign pma_checker_pmp__EVAL_32 = 2'h0;
  assign _EVAL_982 = _EVAL_351 | _EVAL_990;
  assign _EVAL_727 = _EVAL_71;
  assign _EVAL_456 = q__EVAL_5;
  assign _EVAL_451 = _EVAL_860[5:0];
  assign _EVAL_680 = _EVAL_780 ? _EVAL_1297 : 32'h0;
  assign _EVAL_446 = |_EVAL_471;
  assign _EVAL_906 = _EVAL_1217 ? _EVAL_433 : _EVAL_1342;
  assign _EVAL_204 = _EVAL_233 ? 3'h5 : 3'h6;
  assign _EVAL_1191 = _EVAL_1278 == 5'h0;
  assign _EVAL_533 = _EVAL_1306[0];
  assign _EVAL_810 = _EVAL_49;
  assign _EVAL_542 = _EVAL_403 | _EVAL_770;
  assign _EVAL_767 = _EVAL_943 == 5'h0;
  assign _EVAL_495 = _EVAL_422 & _EVAL_489;
  assign _EVAL_867 = _EVAL_618 ? 3'h4 : _EVAL_364;
  assign _EVAL_192 = _EVAL_618 ? _EVAL_1331 : _EVAL_1232;
  assign _EVAL_648 = 8'h1 << _EVAL_1387;
  assign _EVAL_303 = 4'h4 == _EVAL_733;
  assign _EVAL_532 = _EVAL_428 | _EVAL_964;
  assign _EVAL_1170 = _EVAL_780 ? _EVAL_1288 : 2'h0;
  assign _EVAL_1165 = _EVAL_337 & _EVAL_1181;
  assign _EVAL_376 = _EVAL_1185 | _EVAL_1219;
  assign _EVAL_401 = _EVAL_351 ? 2'h2 : _EVAL_1250;
  assign _EVAL_20 = _EVAL_696;
  assign _EVAL_729 = _EVAL_651 ? _EVAL_1278 : _EVAL_1351;
  assign _EVAL_1083 = _EVAL_943 == 5'h5;
  assign _EVAL_963 = _EVAL_878 & _EVAL_367;
  assign _EVAL_1092 = {_EVAL_972,_EVAL_1356};
  assign _EVAL_845 = _EVAL_935 | _EVAL_319;
  assign _EVAL_262 = _EVAL_308[15:0];
  assign _EVAL_137 = |_EVAL_326;
  assign _EVAL_416 = _EVAL_998 & _EVAL_634;
  assign _EVAL_970 = _EVAL_412 == _EVAL_318;
  assign pma_checker_pmp__EVAL_31 = 2'h0;
  assign tlb_pmp__EVAL_30 = _EVAL_477;
  assign _EVAL_307 = _EVAL_1278 == 5'h17;
  assign _EVAL_283 = 4'he == _EVAL_733;
  assign pma_checker_pmp__EVAL_61 = 1'h0;
  assign _EVAL_1134 = {_EVAL_500,_EVAL_1045};
  assign _EVAL_332 = _EVAL_1351 == 5'hf;
  assign _EVAL_1008 = _EVAL_722 & _EVAL_378;
  assign _EVAL_619 = _EVAL_555 ? 16'hffff : 16'h0;
  assign _EVAL_565 = _EVAL_1067[7:0];
  assign _EVAL_311 = _EVAL_202 | _EVAL_418;
  assign _EVAL_317 = _EVAL_22;
  assign _EVAL_69 = ~_EVAL_349;
  assign _EVAL_518 = _EVAL_1352 ? 3'h1 : _EVAL_784;
  assign _EVAL_420 = |_EVAL_701;
  assign _EVAL_1144 = _EVAL_76;
  assign _EVAL_873 = _EVAL_758[15];
  assign pma_checker_pmp__EVAL_28 = 32'h0;
  assign _EVAL_835 = _EVAL_943 == 5'hc;
  assign _EVAL_1146 = _EVAL_29;
  assign _EVAL_388 = _EVAL_487 | _EVAL_1307;
  assign _EVAL_1132 = ~_EVAL_305;
  assign _EVAL_932 = _EVAL_1033 ? 1'h0 : _EVAL_971;
  assign _EVAL_647 = _EVAL_502 ? _EVAL_1054 : _EVAL_236;
  assign _EVAL_353 = {_EVAL_941,_EVAL_168};
  assign _EVAL_1064 = _EVAL_98 == 5'h9;
  assign _EVAL_969 = _EVAL_336 & _EVAL_993;
  assign _EVAL_161 = _EVAL_404 ? _EVAL_1331 : _EVAL_720;
  assign pma_checker_pmp__EVAL_53 = 30'h0;
  assign _EVAL_1151 = _EVAL_1247 ? _EVAL_323 : _EVAL_154;
  assign _EVAL_134 = ~_EVAL_1078;
  assign _EVAL_947 = _EVAL_503 | _EVAL_166;
  assign _EVAL_1199 = _EVAL_963 ? 2'h3 : 2'h0;
  assign _EVAL_731 = {_EVAL_253,_EVAL_1127,_EVAL_973,_EVAL_1229};
  assign _EVAL_1182 = _EVAL_422[31:12];
  assign _EVAL_902 = _EVAL_479 | _EVAL_450;
  assign _EVAL_1021 = ~_EVAL_1184;
  assign q__EVAL_25 = _EVAL_153 ? _EVAL_731 : _EVAL_754;
  assign _EVAL_774 = _EVAL_716[31:12];
  assign _EVAL_391 = _EVAL_1226 ? 14'h1fff : 14'h0;
  assign _EVAL_473 = {_EVAL_1389,_EVAL_607};
  assign _EVAL_240 = _EVAL_1284 & _EVAL_1016;
  assign _EVAL_193 = ~_EVAL_1339;
  assign _EVAL_894 = _EVAL_768 | _EVAL_307;
  assign _EVAL_768 = _EVAL_396 | _EVAL_324;
  assign _EVAL_99 = _EVAL_105 & _EVAL_101;
  assign _EVAL_95 = _EVAL_589;
  assign _EVAL_222 = _EVAL_37;
  assign _EVAL_1172 = 4'h0 == _EVAL_733;
  assign _EVAL_765 = _EVAL_350 | _EVAL_631;
  assign _EVAL_276 = _EVAL_488[1:0];
  assign _EVAL_915 = _EVAL_7;
  assign _EVAL_487 = _EVAL_229[0];
  assign _EVAL_421 = _EVAL_12;
  assign tlb_pmp__EVAL_51 = _EVAL_587;
  assign _EVAL_492 = _EVAL_118;
  assign _EVAL_285 = _EVAL_703 & _EVAL_686;
  assign _EVAL_702 = _EVAL_63;
  assign _EVAL_897 = _EVAL_1382 | _EVAL_513;
  assign _EVAL_852 = _EVAL_921 & _EVAL_1155;
  assign _EVAL_560 = _EVAL_1019 | _EVAL_255;
  assign _EVAL_212 = $signed(_EVAL_280) == 33'sh0;
  assign _EVAL_990 = _EVAL_394 | _EVAL_1150;
  assign _EVAL_595 = _EVAL_113;
  assign _EVAL_1093 = ~_EVAL_1055;
  assign _EVAL_632 = _EVAL_1091;
  assign _EVAL_796 = ~_EVAL_1320;
  assign _EVAL_214 = _EVAL_308[31:16];
  assign _EVAL_652 = _EVAL_1035 | _EVAL_1242;
  assign _EVAL_11 = _EVAL_1267 & _EVAL_1264;
  assign _EVAL_243 = _EVAL_1239 | _EVAL_141;
  assign _EVAL_986 = _EVAL_10;
  assign _EVAL_583 = _EVAL_1211 | _EVAL_759;
  assign pma_checker_pmp__EVAL_1 = 30'h0;
  assign _EVAL_640 = ~_EVAL_1110;
  assign _EVAL_117 = _EVAL_1205 & _EVAL_1217;
  assign _EVAL_1201 = _EVAL_472 | _EVAL_708;
  assign _EVAL_591 = _EVAL_919 ? 8'hff : 8'h0;
  assign _EVAL_232 = _EVAL_684 | _EVAL_1350;
  assign _EVAL_757 = _EVAL_1217 ? _EVAL_388 : _EVAL_1307;
  assign _EVAL_1369 = _EVAL_293;
  assign _EVAL_1363 = $signed(_EVAL_267) & 33'sheb004000;
  assign _EVAL_148 = _EVAL_404 ? _EVAL_323 : _EVAL_408;
  assign _EVAL_621 = _EVAL_108;
  assign _EVAL_270 = _EVAL_61;
  assign _EVAL_38 = _EVAL_1366;
  assign _EVAL_1106 = _EVAL_673 ? 3'h2 : _EVAL_1222;
  assign _EVAL_159 = _EVAL_946 ? _EVAL_1050 : _EVAL_1087;
  assign _EVAL_941 = _EVAL_1271[31:14];
  assign _EVAL_786 = _EVAL_78;
  assign _EVAL_682 = _EVAL_66;
  assign _EVAL_1122 = $signed(_EVAL_937) & -33'sh1000;
  assign _EVAL_782 = |_EVAL_133;
  assign _EVAL_655 = {_EVAL_656,_EVAL_1137,_EVAL_1187,_EVAL_1101};
  assign _EVAL_720 = _EVAL_1183 ? _EVAL_1331 : _EVAL_171;
  assign _EVAL_609 = {1'b0,$signed(_EVAL_988)};
  assign _EVAL_394 = 4'h1 == _EVAL_733;
  assign _EVAL_742 = _EVAL_766 ? _EVAL_1329 : _EVAL_321;
  assign _EVAL_819 = _EVAL_82;
  assign q__EVAL_18 = _EVAL_969 | _EVAL_653;
  assign _EVAL_584 = _EVAL_855 ? _EVAL_1310 : 2'h0;
  assign tlb_pmp__EVAL_32 = _EVAL_596;
  assign _EVAL_116 = _EVAL_1328;
  assign _EVAL_1244 = _EVAL_766 ? _EVAL_323 : _EVAL_712;
  assign _EVAL_871 = _EVAL_532 | _EVAL_1094;
  assign _EVAL_462 = _EVAL_1180 ? 2'h3 : 2'h0;
  assign _EVAL_490 = _EVAL_1259[2];
  assign _EVAL_1149 = 4'hc == _EVAL_733;
  assign _EVAL_797 = _EVAL_1057 ? _EVAL_1387 : 3'h0;
  assign _EVAL_1037 = 5'hb == _EVAL_1351;
  assign _EVAL_178 = _EVAL_606 ^ 32'h4000;
  assign _EVAL_1035 = _EVAL_542 | _EVAL_1192;
  assign tlb_pmp__EVAL_56 = _EVAL_252;
  assign _EVAL_187 = _EVAL_845 | _EVAL_215;
  assign _EVAL_1364 = _EVAL_739 | _EVAL_1147;
  assign _EVAL_664 = _EVAL_229[5];
  assign tlb_pmp__EVAL_19 = _EVAL_1118;
  assign _EVAL_1197 = _EVAL_522 ? _EVAL_1241 : 14'h0;
  assign _EVAL_604 = _EVAL_231 & tlb_pmp__EVAL_9;
  assign _EVAL_776 = _EVAL_568 & _EVAL_492;
  assign _EVAL_863 = q__EVAL_4;
  assign _EVAL_176 = _EVAL_943 == 5'hd;
  assign _EVAL_1145 = _EVAL_514 ? _EVAL_764 : _EVAL_868;
  assign _EVAL_559 = _EVAL_1067[15:8];
  assign _EVAL_341 = _EVAL_1215 | _EVAL_418;
  assign _EVAL_368 = _EVAL_881 | _EVAL_149;
  assign _EVAL_587 = _EVAL_103;
  assign _EVAL_766 = 5'hd == _EVAL_1351;
  assign _EVAL_872 = _EVAL_1278 == 5'h11;
  assign _EVAL_1065 = _EVAL_1279 - 7'h1;
  assign _EVAL_1026 = _EVAL_583 | _EVAL_1043;
  assign _EVAL_1075 = _EVAL_957 & _EVAL_305;
  assign q__EVAL_0 = _EVAL_153 ? 32'h0 : _EVAL_895;
  assign _EVAL_577 = _EVAL_201 ? _EVAL_731 : _EVAL_327;
  assign _EVAL_926 = _EVAL_871 ? _EVAL_1375 : _EVAL_662;
  assign _EVAL_1061 = _EVAL_16[31:14];
  assign _EVAL_646 = _EVAL_891 | _EVAL_726;
  assign _EVAL_173 = _EVAL_1296 == 6'h1;
  assign _EVAL_277 = _EVAL_673 ? 3'h0 : _EVAL_867;
  assign _EVAL_971 = 4'hb == _EVAL_1373;
  assign _EVAL_925 = _EVAL_331 | _EVAL_1120;
  assign data__EVAL_5 = gated_clock_dcache_clock_gate_out;
  assign _EVAL_649 = {1'b0,$signed(_EVAL_286)};
  assign _EVAL_606 = {_EVAL_348,_EVAL_1125};
  assign _EVAL_630 = _EVAL_371 & _EVAL_894;
  assign _EVAL_576 = _EVAL_912 & _EVAL_288;
  assign _EVAL_1059 = _EVAL_454;
  assign _EVAL_217 = _EVAL_266 & _EVAL_225;
  assign _EVAL_1010 = ~_EVAL_1241;
  assign _EVAL_751 = _EVAL_765 & _EVAL_918;
  assign _EVAL_639 = _EVAL_303 ? 2'h1 : _EVAL_144;
  assign _EVAL_854 = $signed(_EVAL_882) == 33'sh0;
  assign _EVAL_1230 = _EVAL_776 ? _EVAL_1362 : 2'h1;
  assign _EVAL_882 = _EVAL_1200;
  assign _EVAL_2 = _EVAL_934 & _EVAL_640;
  assign _EVAL_885 = _EVAL_1060 | _EVAL_189;
  assign tlb_pmp__EVAL_17 = _EVAL_1228;
  assign _EVAL_346 = _EVAL_340;
  assign tlb_pmp__EVAL_1 = _EVAL_552;
  assign lfsr_prng__EVAL_11 = gated_clock_dcache_clock_gate_out;
  assign _EVAL_665 = _EVAL_743 ? _EVAL_343 : 6'h0;
  assign _EVAL_806 = ~_EVAL_560;
  assign _EVAL_135 = _EVAL_333 | _EVAL_246;
  assign data__EVAL_0 = _EVAL_825;
  assign _EVAL_1101 = _EVAL_237[0];
  assign _EVAL_464 = ~_EVAL_1365;
  assign _EVAL_968 = _EVAL_1319 & _EVAL_193;
  assign _EVAL_233 = _EVAL_443[5];
  assign _EVAL_302 = _EVAL_1169;
  assign _EVAL_409 = _EVAL_943 == 5'h17;
  assign pma_checker_pmp__EVAL_59 = 1'h0;
  assign _EVAL_482 = _EVAL_16[13:0];
  assign _EVAL_1025 = q__EVAL_3;
  assign _EVAL_1033 = 4'h4 == _EVAL_1373;
  assign _EVAL_848 = _EVAL_1361 | _EVAL_1034;
  assign _EVAL_662 = |_EVAL_453;
  assign tlb_pmp__EVAL_11 = _EVAL_345;
  assign _EVAL_608 = _EVAL_231 & tlb_pmp__EVAL_54;
  assign tlb_pmp__EVAL_49 = _EVAL_599;
  assign _EVAL_210 = ~_EVAL_402;
  assign _EVAL_910 = _EVAL_1067[23:16];
  assign _EVAL_567 = _EVAL_229[2];
  assign tlb_pmp__EVAL_53 = _EVAL_786;
  assign tlb_pmp__EVAL_27 = _EVAL_504;
  assign pma_checker_pmp__EVAL_0 = 32'h0;
  assign _EVAL_1139 = 8'h1 << _EVAL_627;
  assign _EVAL_651 = _EVAL_1347 & _EVAL_685;
  assign _EVAL_18 = _EVAL_151;
  assign _EVAL_1243 = _EVAL_1278 == 5'h9;
  assign _EVAL_221 = _EVAL_668 & _EVAL_661;
  assign gated_clock_dcache_clock_gate_en = _EVAL_1160;
  assign _EVAL_537 = _EVAL_1190[1:0];
  assign _EVAL_992 = _EVAL_98 == 5'h6;
  assign _EVAL_940 = _EVAL_956 ? _EVAL_1087 : _EVAL_791;
  assign _EVAL_582 = q__EVAL_14;
  assign _EVAL_1086 = _EVAL_404 ? _EVAL_1329 : _EVAL_1207;
  assign _EVAL_847 = _EVAL_201 ? _EVAL_1331 : _EVAL_1238;
  assign _EVAL_933 = _EVAL_1333 == _EVAL_562;
  assign pma_checker_pmp__EVAL_41 = 30'h0;
  assign _EVAL_89 = _EVAL_1283;
  assign _EVAL_561 = _EVAL_404 ? 3'h2 : _EVAL_383;
  assign pma_checker_pmp__EVAL_43 = 1'h0;
  assign _EVAL_295 = _EVAL_1184 & _EVAL_1113;
  assign _EVAL_777 = _EVAL_665 == 6'h0;
  assign _EVAL_463 = _EVAL_914 ? _EVAL_731 : _EVAL_563;
  assign _EVAL_424 = |_EVAL_718;
  assign _EVAL_922 = _EVAL_952[0];
  assign _EVAL_785 = _EVAL_513 ? 3'h0 : _EVAL_414;
  assign _EVAL_575 = _EVAL_1259[3];
  assign _EVAL_352 = {1'b0,$signed(_EVAL_529)};
  assign _EVAL_1112 = _EVAL_1306[3];
  assign _EVAL_622 = 4'hd == _EVAL_733;
  assign _EVAL_314 = _EVAL_485;
  assign _EVAL_506 = &_EVAL_133;
  assign _EVAL_455 = _EVAL_938 | _EVAL_1082;
  assign _EVAL_437 = _EVAL_828 | _EVAL_877;
  assign _EVAL_579 = _EVAL_153 ? 3'h4 : _EVAL_496;
  assign _EVAL_685 = ~_EVAL_698;
  assign _EVAL_1215 = _EVAL_316 | _EVAL_300;
  assign _EVAL_546 = _EVAL_1283 == 2'h3;
  assign _EVAL_268 = _EVAL_543 | _EVAL_1340;
  assign _EVAL_431 = _EVAL_1013 & _EVAL_539;
  assign _EVAL_350 = _EVAL_369 == 3'h4;
  assign _EVAL_1357 = _EVAL_914 ? _EVAL_323 : _EVAL_148;
  assign _EVAL_102 = _EVAL_1160;
  assign _EVAL_995 = |_EVAL_945;
  assign _EVAL_860 = _EVAL_1273 - 6'h1;
  assign _EVAL_601 = _EVAL_1047[3];
  assign pma_checker_pmp__EVAL_7 = 2'h0;
  assign _EVAL_832 = _EVAL_1346 > 3'h0;
  assign _EVAL_597 = _EVAL;
  assign _EVAL_1060 = _EVAL_830 | _EVAL_358;
  assign _EVAL_398 = _EVAL_455 | _EVAL_923;
  assign _EVAL_961 = _EVAL_81;
  assign _EVAL_461 = _EVAL_177 | _EVAL_1249;
  assign _EVAL_3 = {_EVAL_1145,_EVAL_1237};
  assign _EVAL_468 = _EVAL_1284[3];
  assign _EVAL_787 = _EVAL_671 ? 1'h0 : _EVAL_989;
  assign _EVAL_1028 = _EVAL_461 | _EVAL_183;
  assign tlb_pmp__EVAL_35 = _EVAL_356;
  assign _EVAL_337 = _EVAL_763[1];
  assign _EVAL_879 = _EVAL_522 & _EVAL_771;
  assign _EVAL_331 = 4'h6 == _EVAL_733;
  assign _EVAL_629 = _EVAL_229[4];
  assign _EVAL_1254 = _EVAL_1296 - 6'h1;
  assign _EVAL_263 = {_EVAL_1305,_EVAL_1291,_EVAL_1304,_EVAL_1335};
  assign _EVAL_1181 = _EVAL_1329[1];
  assign _EVAL_412 = _EVAL_1343[13:2];
  assign _EVAL_1068 = _EVAL_651 ? _EVAL_425 : _EVAL_1329;
  assign _EVAL_964 = _EVAL_1278 == 5'h7;
  assign _EVAL_157 = $signed(_EVAL_609) & 33'sheb004000;
  assign _EVAL_383 = _EVAL_1183 ? 3'h2 : _EVAL_907;
  assign _EVAL_711 = _EVAL_1122;
  assign _EVAL_418 = _EVAL_1351 == 5'h6;
  assign _EVAL_114 = _EVAL_1331;
  assign _EVAL_264 = _EVAL_765 ? _EVAL_390 : 1'h1;
  assign _EVAL_1183 = 5'he == _EVAL_1351;
  assign _EVAL_124 = _EVAL_1351;
  assign _EVAL_886 = |_EVAL_1253;
  assign _EVAL_750 = _EVAL_1278 == 5'hb;
  assign _EVAL_1046 = _EVAL_843 ? _EVAL_602 : 14'h0;
  assign _EVAL_713 = _EVAL_921 & _EVAL_470;
  assign _EVAL_586 = |_EVAL_447;
  assign _EVAL_957 = ~_EVAL_1181;
  assign _EVAL_279 = _EVAL_626 | _EVAL_1157;
  assign _EVAL_645 = _EVAL_272 | _EVAL_1088;
  assign tlb_pmp__EVAL_40 = _EVAL_199;
  assign _EVAL_252 = _EVAL_120;
  assign _EVAL_213 = _EVAL_21;
  assign _EVAL_1207 = _EVAL_1183 ? _EVAL_1329 : _EVAL_742;
  assign pma_checker_pmp__EVAL_21 = 1'h0;
  assign tlb_pmp__EVAL_28 = _EVAL_1144;
  assign _EVAL_1246 = _EVAL_123;
  assign tlb_pmp__EVAL_37 = _EVAL_965;
  assign _EVAL_1044 = _EVAL_1037 ? _EVAL_323 : _EVAL_1151;
  assign tlb_pmp__EVAL_31 = _EVAL_213;
  assign _EVAL_562 = _EVAL_285 | _EVAL_1117;
  assign _EVAL_174 = _EVAL_87;
  assign _EVAL_628 = ~_EVAL_359;
  assign _EVAL_1156 = _EVAL_630 & _EVAL_796;
  assign _EVAL_259 = _EVAL_921 & _EVAL_427;
  assign _EVAL_1067 = _EVAL_42;
  assign _EVAL_503 = _EVAL_943 == 5'h6;
  assign _EVAL_1229 = _EVAL_1138 | _EVAL_987;
  assign _EVAL_1001 = _EVAL_156 & _EVAL_539;
  assign _EVAL_266 = _EVAL_1319 & _EVAL_605;
  assign _EVAL_422 = _EVAL_1311;
  assign _EVAL_1159 = _EVAL_1057 ? _EVAL_1329 : 32'h0;
  assign _EVAL_348 = _EVAL_422[31:12];
  assign _EVAL_1004 = {1'b0,$signed(_EVAL_405)};
  assign _EVAL_1372 = 4'h2 == _EVAL_1373;
  assign pma_checker_pmp__EVAL_2 = 1'h0;
  assign _EVAL_322 = _EVAL_104;
  assign _EVAL_1223 = _EVAL_98 == 5'hf;
  assign _EVAL_1087 = _EVAL_285 | _EVAL_1117;
  assign _EVAL_808 = _EVAL_337 & _EVAL_957;
  assign _EVAL_1232 = _EVAL_1037 ? _EVAL_1331 : _EVAL_884;
  assign _EVAL_824 = |_EVAL_438;
  assign _EVAL_930 = {_EVAL_1070,_EVAL_888};
  assign _EVAL_310 = _EVAL_419 ? 2'h3 : _EVAL_719;
  assign pma_checker_pmp__EVAL_19 = 1'h0;
  assign _EVAL_979 = _EVAL_1217 ? _EVAL_1133 : _EVAL_1330;
  assign _EVAL_475 = _EVAL_1278 == 5'hf;
  assign _EVAL_1039 = _EVAL_1251 & _EVAL_210;
  assign _EVAL_937 = {1'b0,$signed(_EVAL_1359)};
  assign _EVAL_381 = _EVAL_297 ? 2'h2 : _EVAL_639;
  assign tlb_pmp__EVAL_24 = _EVAL_317;
  assign _EVAL_83 = _EVAL_492 & _EVAL_539;
  assign _EVAL_935 = _EVAL_1384 | _EVAL_1056;
  assign _EVAL_568 = _EVAL_1053;
  assign tlb_pmp__EVAL_25 = _EVAL_249;
  assign _EVAL_700 = 4'h3 == _EVAL_733;
  assign _EVAL_364 = _EVAL_1037 ? 3'h2 : _EVAL_1236;
  assign _EVAL_696 = q__EVAL_11;
  assign _EVAL_1077 = _EVAL_39[0];
  assign _EVAL_761 = _EVAL_1077 | _EVAL_88;
  assign _EVAL_379 = _EVAL_680 | _EVAL_234;
  assign _EVAL_479 = _EVAL_242 | _EVAL_1243;
  assign _EVAL_50 = _EVAL_1267 & _EVAL_1277;
  assign tlb_pmp__EVAL_42 = _EVAL_222;
  assign _EVAL_566 = 4'h1 << _EVAL_1231;
  assign _EVAL_1376 = _EVAL_41;
  assign _EVAL_1094 = _EVAL_1234 | _EVAL_833;
  assign _EVAL_594 = _EVAL_167 ? _EVAL_1010 : 14'h0;
  assign _EVAL_288 = _EVAL_98 == 5'h11;
  assign _EVAL_683 = _EVAL_1191 | _EVAL_865;
  assign _EVAL_1155 = _EVAL_1351 == 5'h17;
  assign data__EVAL_4 = _EVAL_940;
  assign _EVAL_1015 = _EVAL_550 ? 1'h0 : _EVAL_264;
  assign _EVAL_280 = _EVAL_448;
  assign _EVAL_339 = _EVAL_1273 == 6'h1;
  assign _EVAL_1129 = _EVAL_1134;
  assign _EVAL_735 = _EVAL_679[1];
  assign q__EVAL_23 = _EVAL_153 ? 3'h0 : _EVAL_785;
  assign _EVAL_414 = _EVAL_914 ? 3'h0 : _EVAL_1085;
  assign tlb_pmp__EVAL_57 = _EVAL_1023;
  assign _EVAL_166 = _EVAL_943 == 5'h7;
  assign _EVAL_618 = 5'h8 == _EVAL_1351;
  assign _EVAL_929 = _EVAL_761 | _EVAL_1251;
  assign _EVAL_1079 = q__EVAL_13;
  assign _EVAL_1012 = _EVAL_276 & 2'h1;
  assign _EVAL_846 = _EVAL_788 | _EVAL_835;
  assign _EVAL_668 = _EVAL_831 & _EVAL_1333;
  assign _EVAL_788 = _EVAL_943 == 5'h8;
  assign _EVAL_795 = _EVAL_410 | _EVAL_407;
  assign _EVAL_1225 = _EVAL_1302 >= 2'h2;
  assign _EVAL_599 = _EVAL_121;
  assign pma_checker_pmp__EVAL_13 = 1'h0;
  assign _EVAL_840 = _EVAL_1284[1];
  assign tlb_pmp__EVAL_59 = _EVAL_129;
  assign _EVAL_411 = $signed(_EVAL_649) & -33'sh4000;
  assign data__EVAL_1 = _EVAL_497;
  assign _EVAL_72 = _EVAL_667;
  assign _EVAL_833 = _EVAL_646 | _EVAL_475;
  assign _EVAL_335 = _EVAL_1363;
  assign _EVAL_1119 = _EVAL_1278 == 5'hc;
  assign _EVAL_526 = _EVAL_1271[1];
  assign _EVAL_1389 = _EVAL_17;
  assign _EVAL_239 = data__EVAL_3;
  assign _EVAL_100 = {_EVAL_344,_EVAL_1096};
  assign _EVAL_1055 = {_EVAL_829,12'h0};
  assign _EVAL_1374 = _EVAL_811 & _EVAL_890;
  assign _EVAL_225 = ~_EVAL_244;
  assign _EVAL_738 = _EVAL_618 ? _EVAL_323 : _EVAL_1044;
  assign pma_checker_pmp__EVAL_35 = 1'h0;
  assign _EVAL_1249 = _EVAL_936 ? _EVAL_1313 : 7'h0;
  assign _EVAL_1231 = _EVAL_1263;
  assign _EVAL_578 = _EVAL_334[1];
  assign _EVAL_253 = _EVAL_342 | _EVAL_205;
  assign _EVAL_1005 = _EVAL_673 ? _EVAL_1331 : _EVAL_192;
  assign _EVAL_390 = ~_EVAL_1115;
  assign _EVAL_433 = _EVAL_567 | _EVAL_1342;
  assign _EVAL_684 = _EVAL_229[6];
  assign _EVAL_359 = {_EVAL_813,12'h0};
  assign _EVAL_557 = _EVAL_423;
  assign _EVAL_1164 = _EVAL_1333 & _EVAL_661;
  assign _EVAL_400 = _EVAL_914 ? _EVAL_1329 : _EVAL_1086;
  assign _EVAL_654 = _EVAL_1022[3:0];
  assign _EVAL_891 = _EVAL_975 | _EVAL_749;
  assign _EVAL_759 = $signed(_EVAL_826) == 33'sh0;
  assign _EVAL_498 = _EVAL_1057 ? 3'h3 : 3'h0;
  assign _EVAL_215 = _EVAL_1351 == 5'hb;
  assign _EVAL_256 = _EVAL_879 ? _EVAL_1010 : 14'h0;
  assign _EVAL_616 = _EVAL_651 & _EVAL_871;
  assign _EVAL_677 = _EVAL_32;
  assign _EVAL_254 = _EVAL_1279 > 7'h0;
  assign _EVAL_858 = _EVAL_766 ? _EVAL_731 : _EVAL_357;
  assign _EVAL_384 = _EVAL_447 ? 8'hff : 8'h0;
  assign _EVAL_1078 = {_EVAL_663,_EVAL_384,_EVAL_591,_EVAL_753};
  assign _EVAL_1166 = _EVAL_1347 | _EVAL_25;
  assign _EVAL_443 = ~_EVAL_133;
  assign _EVAL_434 = _EVAL_846 | _EVAL_176;
  assign _EVAL_509 = _EVAL_947 ? 14'h3fff : 14'h0;
  assign _EVAL_811 = ~_EVAL_812;
  assign _EVAL_955 = _EVAL_306[2:0];
  assign tlb_pmp__EVAL_10 = _EVAL_915;
  assign _EVAL_523 = _EVAL_96;
  assign _EVAL_828 = _EVAL_715 | _EVAL_191;
  assign _EVAL_281 = 1'h0;
  assign _EVAL_491 = _EVAL_812 & _EVAL_528;
  assign _EVAL_927 = _EVAL_1183 ? 3'h2 : _EVAL_160;
  assign _EVAL_404 = 5'hf == _EVAL_1351;
  assign _EVAL_1188 = _EVAL_1012 == 2'h1;
  assign _EVAL_1233 = _EVAL_44;
  assign pma_checker_pmp__EVAL_37 = _EVAL_544;
  assign _EVAL_689 = _EVAL_952[3];
  assign _EVAL_671 = 4'h6 == _EVAL_1373;
  assign _EVAL_1006 = _EVAL_91;
  assign _EVAL_284 = _EVAL_707 ? 1'h0 : _EVAL_643;
  assign _EVAL_1027 = _EVAL_866 ? _EVAL_1298 : 2'h0;
  assign _EVAL_389 = _EVAL_657 | _EVAL_1338;
  assign _EVAL_132 = _EVAL_94;
  assign _EVAL_477 = _EVAL_93;
  assign _EVAL_250 = _EVAL_163 ? 2'h3 : 2'h0;
  assign _EVAL_602 = _EVAL_644 | _EVAL_628;
  assign _EVAL_728 = 23'hff << _EVAL_362;
  assign _EVAL_697 = $signed(_EVAL_1004) & 33'sheb000000;
  assign _EVAL_1214 = _EVAL_93;
  assign _EVAL_1204 = _EVAL_604 ? 2'h3 : 2'h0;
  assign _EVAL_784 = _EVAL_1370 ? 3'h2 : _EVAL_530;
  assign _EVAL_1370 = _EVAL_443[2];
  assign _EVAL_809 = _EVAL_92;
  assign _EVAL_611 = _EVAL_1347 & _EVAL_796;
  assign _EVAL_556 = _EVAL_1333 ? _EVAL_263 : _EVAL_1331;
  assign _EVAL_1368 = ~_EVAL_45;
  assign _EVAL_244 = _EVAL_969 & _EVAL_1025;
  assign _EVAL_791 = _EVAL_1248 & _EVAL_159;
  assign _EVAL_405 = _EVAL_606 ^ 32'h2000000;
  assign _EVAL_715 = _EVAL_1364 | _EVAL_1140;
  assign _EVAL_172 = |_EVAL_892;
  assign _EVAL_1114 = {_EVAL_250,12'h0};
  assign _EVAL_674 = _EVAL_767 | _EVAL_503;
  assign _EVAL_521 = _EVAL_871 ? _EVAL_600 : _EVAL_633;
  assign _EVAL_64 = _EVAL_1345;
  assign _EVAL_690 = _EVAL_855 & _EVAL_539;
  assign _EVAL_1124 = _EVAL_141 ? _EVAL_1093 : 14'h0;
  assign pma_checker_pmp__EVAL_26 = 1'h0;
  assign tlb_pmp__EVAL_38 = {_EVAL_348,_EVAL_1125};
  assign pma_checker_pmp__EVAL_12 = 2'h0;
  assign _EVAL_1105 = _EVAL_957 & _EVAL_1132;
  assign _EVAL_450 = _EVAL_1278 == 5'ha;
  assign pma_checker_pmp__EVAL_5 = 30'h0;
  assign tlb_pmp__EVAL_22 = _EVAL_723;
  assign _EVAL_318 = _EVAL_353[13:2];
  assign _EVAL_558 = _EVAL_1037 ? _EVAL_1387 : _EVAL_289;
  assign pma_checker_pmp__EVAL_51 = 1'h0;
  assign _EVAL_721 = _EVAL_1260 | _EVAL_748;
  assign pma_checker_pmp__EVAL_36 = 1'h0;
  assign _EVAL_1024 = _EVAL_1255 | _EVAL_254;
  assign _EVAL_407 = _EVAL_156 & _EVAL_1270;
  assign _EVAL_1175 = _EVAL_1351 == 5'hd;
  assign _EVAL_754 = _EVAL_513 ? _EVAL_654 : _EVAL_463;
  assign _EVAL_996 = _EVAL_365 ? _EVAL_1275 : 2'h0;
  assign _EVAL_452 = _EVAL_818[7:0];
  assign tlb_pmp__EVAL_26 = _EVAL_1246;
  assign _EVAL_515 = |_EVAL_689;
  assign _EVAL_334 = _EVAL_603 ? _EVAL_1230 : 2'h0;
  assign tlb_pmp__EVAL_16 = _EVAL_523;
  assign q__EVAL_10 = _EVAL_1233;
  assign _EVAL_207 = _EVAL_970 & _EVAL_521;
  assign tlb_pmp__EVAL_33 = _EVAL_727;
  assign _EVAL_146 = _EVAL_1283 == 2'h2;
  assign tlb_pmp__EVAL_15 = _EVAL_1376;
  assign _EVAL_504 = _EVAL_85;
  assign _EVAL_1019 = 4'h3 == _EVAL_1373;
  assign pma_checker_pmp__EVAL_52 = 1'h0;
  assign _EVAL_309 = 4'h7 == _EVAL_1373;
  assign _EVAL_1123 = _EVAL_443[3];
  assign _EVAL_209 = _EVAL_1188 ? 2'h2 : 2'h1;
  assign _EVAL_267 = {1'b0,$signed(_EVAL_870)};
  assign _EVAL_194 = _EVAL_440 ? 3'h4 : _EVAL_204;
  assign _EVAL_319 = _EVAL_1351 == 5'ha;
  assign _EVAL_780 = _EVAL_1047[0];
  assign _EVAL_1361 = _EVAL_1170 | _EVAL_958;
  assign _EVAL_1360 = |_EVAL_623;
  assign _EVAL_1111 = _EVAL_1108[15:8];
  assign _EVAL_669 = _EVAL_98 == 5'h3;
  assign _EVAL_1173 = _EVAL_936 & _EVAL_539;
  assign _EVAL_657 = _EVAL_1319 & _EVAL_316;
  assign _EVAL_760 = _EVAL_201 ? _EVAL_1387 : _EVAL_797;
  assign _EVAL_372 = $signed(_EVAL_1004) & -33'sh10000;
  assign _EVAL_1355 = _EVAL_897 | _EVAL_197;
  assign _EVAL_152 = _EVAL_1083 | _EVAL_409;
  assign _EVAL_1354 = _EVAL_556[15:8];
  assign _EVAL_942 = ~_EVAL_295;
  assign _EVAL_188 = _EVAL_1013 & _EVAL_1299;
  assign _EVAL_1002 = _EVAL_58;
  assign _EVAL_481 = _EVAL_97;
  assign _EVAL_286 = _EVAL_606 ^ 32'h1800000;
  assign _EVAL_732 = _EVAL_1037 ? _EVAL_1329 : _EVAL_740;
  assign _EVAL_1193 = _EVAL_84;
  assign _EVAL_923 = _EVAL_1013 ? _EVAL_1312 : 32'h0;
  assign _EVAL_551 = _EVAL_149 ? _EVAL_374 : 14'h0;
  assign _EVAL_749 = _EVAL_1278 == 5'hd;
  assign _EVAL_679 = {_EVAL_678,_EVAL_446,_EVAL_158,_EVAL_886};
  assign _EVAL_889 = |_EVAL_919;
  assign _EVAL_573 = _EVAL_376 | _EVAL_1175;
  assign _EVAL_466 = _EVAL_1217 ? _EVAL_483 : _EVAL_1303;
  assign tlb_pmp__EVAL_41 = _EVAL_961;
  assign tlb_pmp__EVAL_4 = _EVAL_1383;
  assign _EVAL_453 = _EVAL_1306 & _EVAL_1016;
  assign _EVAL_938 = _EVAL_756 | _EVAL_190;
  assign _EVAL_227 = _EVAL_391 & 14'h2000;
  assign _EVAL_1222 = _EVAL_618 ? 3'h2 : _EVAL_966;
  assign _EVAL_231 = _EVAL_878 & _EVAL_856;
  assign _EVAL_164 = _EVAL_766 ? _EVAL_1387 : _EVAL_219;
  assign _EVAL_387 = _EVAL_943 == 5'h9;
  assign _EVAL_907 = _EVAL_766 ? 3'h2 : _EVAL_1106;
  assign _EVAL_1208 = _EVAL_546 | _EVAL_146;
  assign _EVAL_408 = _EVAL_1183 ? _EVAL_323 : _EVAL_1244;
  assign _EVAL_349 = _EVAL_849 | _EVAL_782;
  assign _EVAL_653 = _EVAL_281 & _EVAL_806;
  assign _EVAL_326 = _EVAL_952[2];
  assign _EVAL_1365 = _EVAL_728[7:0];
  assign _EVAL_1388 = ~_EVAL_265;
  assign _EVAL_547 = _EVAL_404 ? _EVAL_1387 : _EVAL_706;
  assign _EVAL_975 = _EVAL_581 | _EVAL_1119;
  assign tlb_pmp__EVAL_23 = _EVAL_322;
  assign _EVAL_505 = _EVAL_601 & _EVAL_539;
  assign _EVAL_529 = _EVAL_606 ^ 32'h20000000;
  assign _EVAL_1109 = _EVAL_573 | _EVAL_875;
  assign _EVAL_943 = _EVAL_1287;
  assign _EVAL_834 = _EVAL_274 & 14'h2000;
  assign _EVAL_956 = _EVAL_285 | _EVAL_1117;
  assign _EVAL_1216 = {1'b0,$signed(_EVAL_851)};
  assign _EVAL_747 = _EVAL_481 | _EVAL_132;
  assign tlb_pmp__EVAL_21 = _EVAL_621;
  assign _EVAL_1185 = _EVAL_1351 == 5'h8;
  assign _EVAL_1378 = _EVAL_691 ? _EVAL_619 : _EVAL_214;
  assign _EVAL_920 = _EVAL_714 | _EVAL_931;
  assign pma_checker_pmp__EVAL_20 = 30'h0;
  assign _EVAL_1138 = _EVAL_1225 | _EVAL_808;
  assign _EVAL_535 = _EVAL_80;
  assign _EVAL_624 = _EVAL_437 | _EVAL_211;
  assign _EVAL_415 = _EVAL_930[13:0];
  assign _EVAL_1380 = _EVAL_658 | _EVAL_1333;
  assign _EVAL_358 = _EVAL_855 ? _EVAL_1323 : 7'h0;
  assign _EVAL_347 = _EVAL_98 == 5'hd;
  assign _EVAL_1260 = _EVAL_389 & _EVAL_815;
  assign _EVAL_1252 = _EVAL_526 ? 2'h0 : _EVAL_1131;
  assign _EVAL_1251 = _EVAL_1021 | _EVAL_677;
  assign data__EVAL_2 = _EVAL_220;
  assign _EVAL_540 = 4'h1 == _EVAL_1373;
  assign _EVAL_895 = _EVAL_513 ? _EVAL_1331 : _EVAL_585;
  assign _EVAL_877 = $signed(_EVAL_1377) == 33'sh0;
  assign _EVAL_1084 = _EVAL_943 == 5'ha;
  assign _EVAL_196 = ~_EVAL_1306;
  assign _EVAL_367 = _EVAL_1026 | _EVAL_854;
  assign _EVAL_896 = _EVAL_969 | _EVAL_653;
  assign _EVAL_829 = _EVAL_442 ? 2'h3 : 2'h0;
  assign _EVAL_1248 = _EVAL_946 ? _EVAL_772 : _EVAL_1071;
  assign _EVAL_476 = _EVAL_201 ? 3'h3 : _EVAL_498;
  assign _EVAL_345 = _EVAL_65;
  assign _EVAL_1219 = _EVAL_1351 == 5'hc;
  assign _EVAL_1023 = _EVAL_75;
  assign _EVAL_427 = _EVAL_920 | _EVAL_316;
  assign _EVAL_459 = _EVAL_1224;
  assign _EVAL_1184 = ~_EVAL_981;
  assign _EVAL_467 = _EVAL_885 | _EVAL_1174;
  assign _EVAL_874 = {_EVAL_1378,_EVAL_758};
  assign _EVAL_308 = {_EVAL_862,_EVAL_836,_EVAL_228,_EVAL_480};
  assign _EVAL_580 = _EVAL_513 ? _EVAL_1387 : _EVAL_241;
  assign _EVAL_282 = |_EVAL_533;
  assign _EVAL_502 = _EVAL_1110 & _EVAL_1388;
  assign _EVAL_435 = _EVAL_844 | _EVAL_1094;
  assign _EVAL_838 = _EVAL_1259[1];
  assign _EVAL_145 = _EVAL_331 ? 2'h2 : _EVAL_310;
  assign _EVAL_1241 = {_EVAL_1199,12'h0};
  assign _EVAL_1103 = _EVAL_313[13:0];
  assign _EVAL_333 = $signed(_EVAL_302) == 33'sh0;
  assign _EVAL_726 = _EVAL_1278 == 5'he;
  assign _EVAL_9 = _EVAL_1040;
  assign _EVAL_301 = _EVAL_434 | _EVAL_693;
  assign _EVAL_1047 = _EVAL_1139[6:0];
  assign _EVAL_865 = _EVAL_1278 == 5'h6;
  assign _EVAL_448 = $signed(_EVAL_208) & 33'sh40000000;
  assign _EVAL_1066 = _EVAL_62;
  assign _EVAL_633 = |_EVAL_240;
  assign _EVAL_890 = _EVAL_1379 | _EVAL_652;
  assign _EVAL_638 = _EVAL_831 & _EVAL_924;
  assign _EVAL_625 = _EVAL_74;
  assign _EVAL_444 = _EVAL_1065[6:0];
  assign q__EVAL = _EVAL_93;
  assign _EVAL_708 = _EVAL_98 == 5'hc;
  assign _EVAL_1117 = _EVAL_610 & _EVAL_268;
  assign _EVAL_1240 = _EVAL_943 == 5'hf;
  assign _EVAL_202 = _EVAL_1351 == 5'h0;
  assign _EVAL_530 = _EVAL_1123 ? 3'h3 : _EVAL_194;
  assign _EVAL_769 = _EVAL_556[31:24];
  assign _EVAL_119 = {_EVAL_344,_EVAL_1096};
  assign _EVAL_1259 = {_EVAL_525,_EVAL_586,_EVAL_889,_EVAL_282};
  assign _EVAL_763 = _EVAL_903 | 2'h1;
  assign _EVAL_1250 = _EVAL_394 ? 2'h1 : _EVAL_974;
  assign _EVAL_1189 = _EVAL_1121;
  assign _EVAL_219 = _EVAL_673 ? _EVAL_1387 : _EVAL_1227;
  assign _EVAL_550 = _EVAL_631 & _EVAL_510;
  assign _EVAL_1375 = |_EVAL_1008;
  assign _EVAL_163 = _EVAL_878 & _EVAL_645;
  assign _EVAL_989 = _EVAL_737 ? 1'h0 : _EVAL_932;
  assign _EVAL_615 = _EVAL_874[7:0];
  assign _EVAL_392 = {1'b0,$signed(_EVAL_779)};
  assign _EVAL_1137 = _EVAL_237[2];
  assign _EVAL_804 = _EVAL_1;
  assign _EVAL_211 = $signed(_EVAL_1189) == 33'sh0;
  assign _EVAL_1221 = _EVAL_1102[3:0];
  assign amoalu__EVAL_2 = _EVAL_1331;
  assign pma_checker_pmp__EVAL_40 = 2'h0;
  assign _EVAL_1190 = _EVAL_398 | _EVAL_704;
  assign _EVAL_870 = _EVAL_606 ^ 32'h1000000;
  assign _EVAL_237 = {_EVAL_251,_EVAL_995,_EVAL_1049,_EVAL_824};
  assign _EVAL_293 = $signed(_EVAL_893) & 33'sheb000000;
  assign _EVAL_1379 = _EVAL_131 | _EVAL_789;
  assign _EVAL_489 = {{28'd0}, _EVAL_1221};
  assign _EVAL_718 = _EVAL_594 & 14'h2000;
  assign _EVAL_707 = 4'h0 == _EVAL_1373;
  assign _EVAL_821 = _EVAL_1108[23:16];
  assign _EVAL_1107 = _EVAL_368 | _EVAL_166;
  assign _EVAL_356 = _EVAL_126;
  assign _EVAL_1110 = _EVAL_713 & _EVAL_427;
  assign _EVAL_1352 = _EVAL_443[1];
  assign _EVAL_241 = _EVAL_914 ? _EVAL_1387 : _EVAL_547;
  assign _EVAL_661 = ~_EVAL_562;
  assign pma_checker_pmp__EVAL_57 = 1'h0;
  assign _EVAL_454 = $signed(_EVAL_392) & -33'sh400000;
  assign _EVAL_762 = _EVAL_1302[0];
  assign pma_checker_pmp__EVAL_47 = 2'h0;
  assign _EVAL_815 = _EVAL_484 & _EVAL_926;
  assign _EVAL_1176 = _EVAL_1237[7];
  assign pma_checker_pmp__EVAL_11 = 2'h0;
  assign _EVAL_673 = 5'hc == _EVAL_1351;
  assign _EVAL_770 = _EVAL_98 == 5'ha;
  assign _EVAL_180 = 4'h7 == _EVAL_733;
  assign _EVAL_1362 = _EVAL_765 ? 2'h1 : _EVAL_209;
  assign pma_checker_pmp__EVAL_4 = 1'h0;
  assign _EVAL_1387 = _EVAL_741 ? 3'h0 : _EVAL_518;
  assign _EVAL_141 = _EVAL_301 | _EVAL_1240;
  assign pma_checker_pmp__EVAL_46 = 32'h0;
  assign _EVAL_169 = _EVAL_871 & _EVAL_872;
  assign _EVAL_538 = _EVAL_371 & _EVAL_1186;
  assign _EVAL_1116 = _EVAL_1278 == 5'h14;
  assign _EVAL_678 = |_EVAL_822;
  assign _EVAL_820 = _EVAL_1278 == 5'h5;
  assign _EVAL_1373 = {2'h2,_EVAL_1027};
  assign _EVAL_1202 = _EVAL_579[2];
  assign _EVAL_1247 = 5'ha == _EVAL_1351;
  assign _EVAL_855 = _EVAL_1047[4];
  assign _EVAL_147 = _EVAL_983 | _EVAL_462;
  assign _EVAL_1187 = _EVAL_237[1];
  assign _EVAL_853 = q__EVAL_7;
  assign _EVAL_438 = _EVAL_1284[0];
  assign _EVAL_1140 = $signed(_EVAL_953) == 33'sh0;
  assign _EVAL_374 = ~_EVAL_1114;
  assign tlb_pmp__EVAL_50 = _EVAL_143;
  assign _EVAL_1043 = $signed(_EVAL_1369) == 33'sh0;
  assign pma_checker_pmp__EVAL_60 = 1'h0;
  assign _EVAL_827 = ~_EVAL_730;
  assign tlb_pmp__EVAL_8 = _EVAL_273;
  assign _EVAL_771 = _EVAL_1107 | _EVAL_243;
  assign _EVAL_321 = _EVAL_673 ? _EVAL_1329 : _EVAL_140;
  assign _EVAL_588 = _EVAL_805 | _EVAL_669;
  assign _EVAL_571 = ~_EVAL_956;
  assign _EVAL_177 = _EVAL_780 ? _EVAL_1325 : 7'h0;
  assign _EVAL_672 = _EVAL_601 ? _EVAL_1301 : 7'h0;
  assign _EVAL_26 = _EVAL_582;
  assign _EVAL_149 = _EVAL_943 == 5'h11;
  assign _EVAL_703 = _EVAL_389 & _EVAL_1333;
  assign _EVAL_884 = _EVAL_1247 ? _EVAL_1331 : _EVAL_847;
  assign _EVAL_730 = _EVAL_956 | _EVAL_1248;
  assign _EVAL_292 = _EVAL_1206 | _EVAL_817;
  assign _EVAL_403 = _EVAL_1062 | _EVAL_1064;
  assign _EVAL_1045 = {_EVAL_519,_EVAL_1178};
  assign _EVAL_667 = q__EVAL_12;
  assign _EVAL_205 = _EVAL_216 & _EVAL_783;
  assign pma_checker_pmp__EVAL_8 = 1'h0;
  assign _EVAL_658 = _EVAL_642 | _EVAL_1338;
  assign _EVAL_1120 = _EVAL_419 | _EVAL_283;
  assign _EVAL_981 = _EVAL_502 | _EVAL_386;
  assign q__EVAL_27 = _EVAL_1208 | _EVAL_807;
  assign _EVAL_269 = {_EVAL_1061,_EVAL_482};
  assign pma_checker_pmp__EVAL_55 = 1'h0;
  assign _EVAL_1237 = _EVAL_305 ? _EVAL_298 : _EVAL_615;
  assign _EVAL_1211 = $signed(_EVAL_557) == 33'sh0;
  assign _EVAL_706 = _EVAL_1183 ? _EVAL_1387 : _EVAL_164;
  assign _EVAL_1097 = ~_EVAL_1202;
  assign _EVAL_1096 = {_EVAL_228,_EVAL_480};
  assign _EVAL_298 = _EVAL_874[15:8];
  assign tlb_pmp__EVAL_2 = _EVAL_421;
  assign _EVAL_991 = {{30'd0}, _EVAL_537};
  assign _EVAL_242 = _EVAL_1278 == 5'h4;
  assign _EVAL_610 = _EVAL_638 | _EVAL_1333;
  assign _EVAL_798 = _EVAL_458 | _EVAL_1318;
  assign _EVAL_484 = _EVAL_531 == _EVAL_318;
  assign _EVAL_323 = {{2'd0}, _EVAL_1302};
  assign _EVAL_1049 = |_EVAL_840;
  assign _EVAL_1113 = _EVAL_1160;
  assign _EVAL_1102 = _EVAL_566 - 4'h1;
  assign _EVAL_488 = _EVAL_51;
  assign _EVAL_1070 = _EVAL_1286[31:14];
  assign _EVAL_1196 = _EVAL_651 ? _EVAL_1341 : _EVAL_1268;
  assign tlb_pmp__EVAL_7 = _EVAL_1098;
  assign _EVAL_447 = _EVAL_1306[2];
  assign _EVAL_1131 = {_EVAL_417,_EVAL_230};
  assign _EVAL_779 = _EVAL_606 ^ 32'hc000000;
  assign _EVAL_151 = q__EVAL_21;
  assign _EVAL_430 = _EVAL_1271[11:0];
  assign _EVAL_70 = _EVAL_946 ? _EVAL_699 : _EVAL_439;
  assign _EVAL_510 = ~_EVAL_571;
  assign _EVAL_410 = _EVAL_694 | _EVAL_1030;
  assign _EVAL_1042 = _EVAL_1103;
  assign _EVAL_257 = _EVAL_1248 ? _EVAL_1042 : _EVAL_984;
  assign pma_checker_pmp__EVAL_44 = 1'h0;
  assign _EVAL_183 = _EVAL_156 ? _EVAL_1314 : 7'h0;
  assign _EVAL_841 = _EVAL_618 ? _EVAL_731 : _EVAL_801;
  assign tlb_pmp__EVAL_61 = _EVAL_393;
  assign _EVAL_620 = _EVAL_549 | _EVAL_1009;
  assign _EVAL_880 = {1'b0,$signed(_EVAL_178)};
  assign _EVAL_563 = _EVAL_404 ? _EVAL_731 : _EVAL_139;
  assign _EVAL_753 = _EVAL_533 ? 8'hff : 8'h0;
  assign _EVAL_182 = _EVAL_1317 >= 2'h1;
  assign _EVAL_953 = _EVAL_411;
  assign _EVAL_756 = _EVAL_379 | _EVAL_441;
  assign _EVAL_1157 = _EVAL_855 & _EVAL_1289;
  assign _EVAL_758 = _EVAL_1181 ? _EVAL_214 : _EVAL_262;
  assign _EVAL_1085 = _EVAL_404 ? 3'h3 : _EVAL_927;
  assign _EVAL_1126 = ~_EVAL_470;
  assign _EVAL_544 = gated_clock_dcache_clock_gate_out;
  assign _EVAL_1011 = _EVAL_1296 == 6'h0;
  assign _EVAL_480 = _EVAL_1308[7:0];
  assign _EVAL_483 = _EVAL_1198 | _EVAL_1303;
  assign _EVAL_704 = _EVAL_365 ? _EVAL_1269 : 32'h0;
  assign _EVAL_1056 = _EVAL_1351 == 5'h9;
  assign _EVAL_802 = _EVAL_914 ? 3'h0 : _EVAL_561;
  assign _EVAL_1142 = $signed(_EVAL_459) == 33'sh0;
  assign _EVAL_519 = |_EVAL_949;
  assign tlb_pmp__EVAL_55 = _EVAL_909;
  assign _EVAL_1100 = {_EVAL_1061,_EVAL_415};
  assign _EVAL_130 = _EVAL_1217 ? _EVAL_798 : _EVAL_1318;
  assign _EVAL_313 = _EVAL_1333 ? _EVAL_1343 : _EVAL_1295;
  assign _EVAL_596 = _EVAL_67;
  assign _EVAL_1150 = _EVAL_180 | _EVAL_925;
  assign tlb_pmp__EVAL_52 = _EVAL_702;
  assign _EVAL_1385 = ~_EVAL_481;
  assign _EVAL_273 = _EVAL_40;
  assign _EVAL_191 = $signed(_EVAL_346) == 33'sh0;
  assign _EVAL_329 = ~_EVAL_25;
  assign _EVAL_951 = q__EVAL_16;
  assign pma_checker_pmp__EVAL_16 = 2'h0;
  assign _EVAL_959 = _EVAL_238 ? _EVAL_239 : 32'h0;
  assign _EVAL_659 = _EVAL_556[7:0];
  assign _EVAL_1174 = _EVAL_365 ? _EVAL_1321 : 7'h0;
  assign _EVAL_1228 = _EVAL_30;
  assign _EVAL_1200 = $signed(_EVAL_1216) & 33'sheb002000;
  assign _EVAL_893 = {1'b0,$signed(_EVAL_426)};
  assign tlb_pmp__EVAL_34 = _EVAL_1002;
  assign _EVAL_973 = _EVAL_1138 | _EVAL_752;
  assign _EVAL_393 = _EVAL_47;
  assign _EVAL_1108 = _EVAL_636 | _EVAL_976;
  assign _EVAL_1016 = {_EVAL_147,_EVAL_1252};
  assign _EVAL_783 = _EVAL_1181 & _EVAL_305;
  assign _EVAL_1003 = _EVAL_1109 | _EVAL_332;
  assign _EVAL_354 = _EVAL_464[7:2];
  assign _EVAL_342 = _EVAL_1225 | _EVAL_1165;
  assign _EVAL_966 = _EVAL_1037 ? 3'h3 : _EVAL_850;
  assign _EVAL_208 = {1'b0,$signed(_EVAL_606)};
  assign _EVAL_522 = |_EVAL_495;
  assign _EVAL_545 = _EVAL_1046 | _EVAL_551;
  assign _EVAL_1366 = q__EVAL_6;
  assign _EVAL_574 = _EVAL_545 | _EVAL_524;
  assign _EVAL_525 = |_EVAL_1112;
  assign _EVAL_634 = _EVAL_425 < 32'h80004000;
  assign _EVAL_861 = _EVAL_1347 & _EVAL_258;
  assign _EVAL_1238 = _EVAL_1057 ? _EVAL_1331 : 32'h0;
  assign _EVAL_361 = _EVAL_513 ? _EVAL_1329 : _EVAL_400;
  assign _EVAL_531 = _EVAL_1295[13:2];
  assign _EVAL_799 = _EVAL_1017 == 6'h0;
  assign tlb_pmp__EVAL_18 = _EVAL_1193;
  assign _EVAL_1206 = $signed(_EVAL_711) == 33'sh0;
  assign _EVAL_954 = _EVAL_679[3];
  assign _EVAL_324 = _EVAL_820 & _EVAL_395;
  assign tlb_pmp__EVAL_6 = _EVAL_1066;
  assign pma_checker_pmp__EVAL_58 = 1'h0;
  assign _EVAL_552 = _EVAL_59;
  assign _EVAL_377 = _EVAL_1279 > 7'h3;
  assign _EVAL_1198 = _EVAL_229[3];
  assign pma_checker_pmp__EVAL_3 = 1'h0;
  assign _EVAL_316 = _EVAL_1355 | _EVAL_931;
  assign _EVAL_1057 = 5'h4 == _EVAL_1351;
  assign _EVAL_501 = _EVAL_1149 ? 2'h1 : 2'h0;
  assign _EVAL_1255 = _EVAL_1380 | _EVAL_782;
  assign _EVAL_402 = _EVAL_502 | _EVAL_386;
  assign _EVAL_737 = 4'h5 == _EVAL_1373;
  assign _EVAL_357 = _EVAL_673 ? _EVAL_731 : _EVAL_841;
  assign _EVAL_1227 = _EVAL_618 ? _EVAL_1387 : _EVAL_558;
  assign _EVAL_167 = _EVAL_522 & _EVAL_1226;
  assign _EVAL_497 = _EVAL_956 ? _EVAL_1103 : _EVAL_257;
  assign _EVAL_919 = _EVAL_1306[1];
  assign _EVAL_1121 = $signed(_EVAL_880) & -33'sh1000;
  assign _EVAL_694 = _EVAL_780 & _EVAL_1348;
  assign tlb_pmp__EVAL_44 = _EVAL_986;
  assign _EVAL_985 = _EVAL_473 <= 3'h3;
  assign _EVAL_53 = _EVAL_1161;
  assign _EVAL_238 = _EVAL_334[0];
  assign _EVAL_905 = _EVAL_16;
  assign _EVAL_555 = _EVAL_1265 & _EVAL_873;
  assign _EVAL_1220 = _EVAL_848 | _EVAL_486;
  assign _EVAL_380 = _EVAL_201 ? 3'h0 : _EVAL_498;
  assign _EVAL_426 = _EVAL_606 ^ 32'h8000000;
  assign _EVAL_494 = {_EVAL_1081,_EVAL_248};
  assign pma_checker_pmp__EVAL_33 = 30'h0;
  assign _EVAL_1356 = _EVAL_16[5:0];
  assign _EVAL_294 = _EVAL_574 | _EVAL_1124;
  assign _EVAL_814 = _EVAL_1265 & _EVAL_1176;
  assign _EVAL_903 = 2'h1 << _EVAL_762;
  assign tlb_pmp__EVAL_0 = _EVAL_1051;
  assign _EVAL_1169 = $signed(_EVAL_208) & 33'she9000000;
  assign _EVAL_1212 = _EVAL_370 | _EVAL_1367;
  assign _EVAL_220 = _EVAL_956 ? _EVAL_494 : _EVAL_590;
  assign lfsr_prng__EVAL_14 = _EVAL_93;
  assign _EVAL_369 = {{1'd0}, _EVAL_276};
  assign _EVAL_258 = _EVAL_435 & _EVAL_721;
  assign _EVAL_185 = _EVAL_679[0];
  assign _EVAL_24 = _EVAL_1268;
  assign _EVAL_976 = _EVAL_308 & _EVAL_134;
  assign _EVAL_736 = _EVAL_8;
  assign _EVAL_236 = _EVAL_386 ? _EVAL_1100 : _EVAL_905;
  assign _EVAL_741 = _EVAL_443[0];
  assign _EVAL_899 = |_EVAL_1371;
  assign _EVAL_600 = |_EVAL_675;
  assign _EVAL_106 = _EVAL_687;
  assign _EVAL_234 = _EVAL_936 ? _EVAL_1322 : 32'h0;
  assign _EVAL_1359 = _EVAL_606 ^ 32'h3000;
  assign _EVAL_13 = _EVAL_853;
  assign _EVAL_1009 = _EVAL_365 & _EVAL_1337;
  assign _EVAL_165 = _EVAL_1172 ? 2'h0 : _EVAL_381;
  assign _EVAL_371 = _EVAL_1347 & _EVAL_1368;
  assign _EVAL_1178 = |_EVAL_922;
  assign amoalu__EVAL_1 = _EVAL_1292;
  assign _EVAL_1210 = _EVAL_365 & _EVAL_539;
  assign _EVAL_631 = _EVAL_369 == 3'h5;
  assign _EVAL_1242 = _EVAL_1235 | _EVAL_1223;
  assign q__EVAL_2 = _EVAL_153 ? 3'h4 : _EVAL_496;
  assign _EVAL_1098 = _EVAL_14;
  assign _EVAL_136 = ~_EVAL_800;
  assign _EVAL_1017 = _EVAL_1097 ? _EVAL_354 : 6'h0;
  assign _EVAL_216 = _EVAL_763[0];
  assign tlb_pmp__EVAL_60 = _EVAL_810;
  assign _EVAL_918 = _EVAL_539 & _EVAL_776;
  assign q__EVAL_1 = _EVAL_153 ? _EVAL_323 : _EVAL_650;
  assign _EVAL_1053 = _EVAL_946 ? 1'h0 : _EVAL_1015;
  assign pma_checker_pmp__EVAL_56 = 1'h0;
  assign _EVAL_803 = |_EVAL_227;
  assign tlb_pmp__EVAL_3 = _EVAL_804;
  assign _EVAL_612 = _EVAL_1247 ? _EVAL_731 : _EVAL_577;
  assign _EVAL_723 = _EVAL_43;
  assign _EVAL_1245 = _EVAL_372;
  assign _EVAL_681 = _EVAL_1057 ? _EVAL_323 : 4'h0;
  assign _EVAL_144 = _EVAL_622 ? 2'h2 : _EVAL_501;
  assign _EVAL_275 = _EVAL_1013 ? _EVAL_1326 : 2'h0;
  assign _EVAL_251 = |_EVAL_468;
  assign _EVAL_1236 = _EVAL_1247 ? 3'h1 : _EVAL_380;
  assign _EVAL_1050 = _EVAL_492 ? 1'h0 : _EVAL_1087;
  assign _EVAL_245 = _EVAL_98 == 5'h0;
  assign _EVAL_56 = _EVAL_568;
  assign _EVAL_179 = _EVAL_1154 | _EVAL_991;
  assign _EVAL_1022 = {{15'd0}, _EVAL_1306};
  assign tlb_pmp__EVAL_5 = _EVAL_270;
  assign _EVAL_457 = _EVAL_700 ? 2'h3 : _EVAL_401;
  assign _EVAL_156 = _EVAL_1047[2];
  assign _EVAL_428 = _EVAL_635 | _EVAL_872;
  assign _EVAL_792 = _EVAL_832 ? _EVAL_955 : _EVAL_1346;
  assign _EVAL_714 = _EVAL_311 | _EVAL_197;
  assign _EVAL_142 = _EVAL_805 | _EVAL_288;
  assign _EVAL_520 = _EVAL_142 | _EVAL_789;
  assign _EVAL_512 = _EVAL_1217 ? _EVAL_1032 : _EVAL_1272;
  assign pma_checker_pmp__EVAL_14 = 1'h0;
  assign _EVAL_590 = _EVAL_1248 ? _EVAL_485 : _EVAL_314;
  assign _EVAL_362 = _EVAL_153 ? _EVAL_323 : _EVAL_650;
  assign _EVAL_1367 = _EVAL_32 & _EVAL_338;
  assign _EVAL_826 = _EVAL_697;
  assign _EVAL_686 = _EVAL_320 | _EVAL_1332;
  assign _EVAL_1224 = $signed(_EVAL_1216) & -33'sh2000;
  assign _EVAL_1218 = ~_EVAL_452;
  assign _EVAL_513 = _EVAL_1351 == 5'h11;
  assign _EVAL_773 = _EVAL_98 == 5'he;
  assign _EVAL_195 = _EVAL_1110 & _EVAL_1388;
  assign _EVAL_297 = 4'h5 == _EVAL_733;
  assign _EVAL_439 = _EVAL_942 ? 1'h0 : _EVAL_312;
  assign _EVAL_564 = _EVAL_425[31:2];
  assign _EVAL_878 = _EVAL_624 | _EVAL_1142;
  assign _EVAL_1034 = _EVAL_156 ? _EVAL_1290 : 2'h0;
  assign _EVAL_140 = _EVAL_618 ? _EVAL_1329 : _EVAL_732;
  assign _EVAL_998 = _EVAL_425 >= 32'h80000000;
  assign _EVAL_1235 = _EVAL_793 | _EVAL_773;
  assign _EVAL_972 = _EVAL_647[31:6];
  assign _EVAL_365 = _EVAL_1047[6];
  assign _EVAL_752 = _EVAL_216 & _EVAL_1075;
  assign _EVAL_850 = _EVAL_1247 ? 3'h3 : _EVAL_476;
  assign _EVAL_471 = _EVAL_1016[2];
  assign _EVAL_636 = amoalu__EVAL & _EVAL_1078;
  assign pma_checker_pmp__EVAL_22 = 1'h0;
  assign _EVAL_805 = _EVAL_98 == 5'h1;
  assign _EVAL_417 = _EVAL_278 | _EVAL_182;
  assign tlb_pmp__EVAL_29 = _EVAL_688;
  assign _EVAL_419 = 4'hf == _EVAL_733;
  assign _EVAL_274 = _EVAL_843 ? 14'h1fff : 14'h0;
  assign _EVAL_549 = _EVAL_279 | _EVAL_188;
  assign _EVAL_440 = _EVAL_443[4];
  assign _EVAL_539 = _EVAL_339 | _EVAL_777;
  assign _EVAL_486 = _EVAL_601 ? _EVAL_1281 : 2'h0;
  assign tlb_pmp__EVAL_13 = _EVAL_535;
  assign _EVAL_338 = ~_EVAL_588;
  assign _EVAL_592 = _EVAL_1108[7:0];
  assign q__EVAL_17 = _EVAL_153 ? _EVAL_1387 : _EVAL_580;
  assign _EVAL_1048 = _EVAL_90;
  assign _EVAL_199 = _EVAL_55;
  assign _EVAL_745 = _EVAL_1259[0];
  assign pma_checker_pmp__EVAL_34 = 32'h0;
  assign _EVAL_739 = _EVAL_292 | _EVAL_960;
  assign _EVAL_1143 = q__EVAL_8;
  assign _EVAL_849 = _EVAL_611 | _EVAL_968;
  assign _EVAL_396 = _EVAL_435 | _EVAL_871;
  assign _EVAL_1253 = _EVAL_1016[0];
  assign _EVAL_1081 = {_EVAL_769,_EVAL_1386};
  assign _EVAL_868 = _EVAL_874[31:8];
  assign _EVAL_569 = _EVAL_679[2];
  assign _EVAL_800 = {_EVAL_1204,12'h0};
  assign _EVAL_201 = 5'h9 == _EVAL_1351;
  assign _EVAL_470 = _EVAL_700 | _EVAL_982;
  assign pma_checker_pmp__EVAL_39 = 32'h0;
  assign _EVAL_719 = _EVAL_283 ? 2'h3 : _EVAL_165;
  assign _EVAL_693 = _EVAL_943 == 5'he;
  assign pma_checker_pmp__EVAL_49 = 1'h0;
  assign _EVAL_1130 = _EVAL_913 | _EVAL_387;
  assign _EVAL_1217 = _EVAL_1025 & _EVAL_896;
  assign _EVAL_960 = $signed(_EVAL_1245) == 33'sh0;
  assign pma_checker_pmp__EVAL_50 = 1'h0;
  assign _EVAL_291 = _EVAL_985 & _EVAL_1147;
  assign _EVAL_635 = _EVAL_1278 == 5'h1;
  assign _EVAL_246 = $signed(_EVAL_335) == 33'sh0;
  assign tlb_pmp__EVAL_46 = _EVAL_1048;
  assign _EVAL_54 = _EVAL_1328 ? _EVAL_1274 : _EVAL_1329;
  assign _EVAL_733 = {_EVAL_316,_EVAL_341,_EVAL_1298};
  assign _EVAL_306 = _EVAL_1346 - 3'h1;
  assign _EVAL_965 = gated_clock_dcache_clock_gate_out;
  assign _EVAL_79 = _EVAL_863;
  assign _EVAL_603 = _EVAL_329 ? _EVAL_1280 : 1'h1;
  assign _EVAL_320 = _EVAL_1347 & _EVAL_871;
  assign _EVAL_442 = _EVAL_878 & _EVAL_212;
  assign _EVAL_496 = _EVAL_513 ? 3'h1 : _EVAL_802;
  assign _EVAL_967 = _EVAL_601 & _EVAL_1266;
  assign _EVAL_980 = _EVAL_674 | _EVAL_166;
  assign _EVAL_1030 = _EVAL_936 & _EVAL_1294;
  assign _EVAL_336 = _EVAL_259 & _EVAL_1126;
  assign pma_checker_pmp__EVAL_23 = 1'h0;
  assign _EVAL_1125 = _EVAL_422[11:0];
  assign pma_checker_pmp__EVAL_17 = 1'h0;
  assign _EVAL_1167 = _EVAL_831 & _EVAL_933;
  assign _EVAL_869 = 1'h0;
  assign _EVAL_793 = _EVAL_1201 | _EVAL_347;
  assign pma_checker_pmp__EVAL_27 = 32'h0;
  assign _EVAL_25 = _EVAL_776 & _EVAL_1188;
  assign _EVAL_862 = _EVAL_1308[31:24];
  assign _EVAL_924 = ~_EVAL_1332;
  assign _EVAL_909 = _EVAL_0;
  assign _EVAL_27 = _EVAL_1267 & _EVAL_1324;
  assign _EVAL_548 = _EVAL_765 & _EVAL_539;
  assign _EVAL_287 = _EVAL_929 | _EVAL_1347;
  assign _EVAL_1088 = $signed(_EVAL_1163) == 33'sh0;
  assign _EVAL_378 = {_EVAL_954,_EVAL_569,_EVAL_735,_EVAL_185};
  assign _EVAL_1115 = _EVAL_1273 == 6'h0;
  assign _EVAL_190 = _EVAL_601 ? _EVAL_1316 : 32'h0;
  assign _EVAL_931 = _EVAL_187 | _EVAL_1003;
  assign _EVAL_445 = ~_EVAL_852;
  assign _EVAL_656 = _EVAL_237[3];
  assign _EVAL_327 = _EVAL_1057 ? _EVAL_731 : 4'h0;
  assign _EVAL_993 = ~_EVAL_506;
  assign _EVAL_644 = _EVAL_1197 | _EVAL_509;
  assign _EVAL_740 = _EVAL_1247 ? _EVAL_1329 : _EVAL_304;
  assign _EVAL_370 = ~_EVAL_827;
  assign _EVAL_1154 = {_EVAL_564, 2'h0};
  assign _EVAL_842 = _EVAL_578 ? _EVAL_1090 : 32'h0;
  assign _EVAL_343 = _EVAL_1218[7:2];
  assign _EVAL_1133 = _EVAL_664 | _EVAL_1330;
  assign _EVAL_709 = _EVAL_2 | _EVAL_195;
  assign _EVAL_1383 = _EVAL_110;
  assign _EVAL_1051 = _EVAL_57;
  assign _EVAL_830 = _EVAL_1028 | _EVAL_672;
  assign _EVAL_712 = _EVAL_673 ? _EVAL_323 : _EVAL_738;
  assign _EVAL_688 = _EVAL_125;
  assign tlb_pmp__EVAL_48 = _EVAL_597;
  assign _EVAL_373 = _EVAL_644 | _EVAL_136;
  assign pma_checker_pmp__EVAL_15 = 1'h0;
  assign _EVAL_818 = 23'hff << _EVAL_174;
  assign _EVAL_158 = |_EVAL_138;
  assign _EVAL_139 = _EVAL_1183 ? _EVAL_731 : _EVAL_858;
  assign _EVAL_1062 = _EVAL_98 == 5'h4;
  assign _EVAL_312 = _EVAL_1374 ? 1'h0 : _EVAL_685;
  assign _EVAL_34 = _EVAL_1267 & _EVAL_1282;
  assign _EVAL_958 = _EVAL_936 ? _EVAL_1344 : 2'h0;
  assign _EVAL_844 = _EVAL_683 | _EVAL_964;
  assign _EVAL_1377 = _EVAL_1029;
  assign _EVAL_363 = |_EVAL_834;
  assign _EVAL_458 = _EVAL_229[1];
  assign _EVAL_831 = _EVAL_725 | _EVAL_1338;
  assign pma_checker_pmp__EVAL_29 = 32'h0;
  assign pma_checker_pmp__EVAL_42 = 30'h0;
  assign _EVAL_950 = _EVAL_1108[31:24];
  assign _EVAL_822 = _EVAL_1016[3];
  assign tlb_pmp__EVAL_12 = _EVAL_682;
  assign pma_checker_pmp__EVAL_25 = 1'h0;
  assign pma_checker_pmp__EVAL_48 = 1'h0;
  assign _EVAL_605 = ~_EVAL_1360;
  assign _EVAL_305 = _EVAL_1329[0];
  assign _EVAL_1226 = _EVAL_980 | _EVAL_243;
  assign _EVAL_987 = _EVAL_216 & _EVAL_1105;
  assign _EVAL_984 = _EVAL_269[13:0];
  assign _EVAL_300 = _EVAL_1351 == 5'h3;
  assign _EVAL_171 = _EVAL_766 ? _EVAL_1331 : _EVAL_1005;
  assign _EVAL_817 = $signed(_EVAL_1059) == 33'sh0;
  assign _EVAL_249 = _EVAL_109;
  assign _EVAL_1082 = _EVAL_855 ? _EVAL_1276 : 32'h0;
  assign _EVAL_499 = _EVAL_943 == 5'hb;
  assign _EVAL_5 = _EVAL_776 & _EVAL_747;
  assign _EVAL_626 = _EVAL_795 | _EVAL_967;
  assign _EVAL_875 = _EVAL_1351 == 5'he;
  assign _EVAL_340 = $signed(_EVAL_609) & -33'sh4000;
  assign _EVAL_1382 = _EVAL_1351 == 5'h1;
  assign _EVAL_1032 = _EVAL_629 | _EVAL_1272;
  assign _EVAL_888 = _EVAL_1329[13:0];
  assign _EVAL_28 = _EVAL_714 | _EVAL_931;
  assign _EVAL_344 = {_EVAL_862,_EVAL_836};
  assign _EVAL_101 = 1'h0;
  assign _EVAL_528 = _EVAL_32 & _EVAL_429;
  assign _EVAL_429 = _EVAL_890 | _EVAL_576;
  assign _EVAL_716 = {_EVAL_1182,_EVAL_1125};
  assign _EVAL_775 = _EVAL_921 & _EVAL_377;
  assign _EVAL_1127 = _EVAL_342 | _EVAL_1020;
  assign _EVAL_1104 = _EVAL_46;
  assign _EVAL_154 = _EVAL_201 ? _EVAL_323 : _EVAL_681;
  assign _EVAL_687 = q__EVAL_15;
  assign _EVAL_1161 = q__EVAL_22;
  assign _EVAL_224 = _EVAL_73;
  assign _EVAL_4 = _EVAL_670;
  assign pma_checker_pmp__EVAL_45 = 30'h0;
  assign _EVAL_1013 = _EVAL_1047[5];
  assign _EVAL_643 = _EVAL_309 | _EVAL_787;
  assign _EVAL_789 = _EVAL_98 == 5'h7;
  assign _EVAL_641 = _EVAL_1226 ? _EVAL_373 : 14'h0;
  always @(posedge _EVAL_112) begin
    _EVAL_1160 <= _EVAL_1024 | _EVAL_832;
  end
  always @(posedge gated_clock_dcache_clock_gate_out) begin
    if (_EVAL_1039) begin
      _EVAL_1263 <= _EVAL_111;
    end
    if (_EVAL_651) begin
      _EVAL_1264 <= _EVAL_363;
    end
    if (_EVAL_776) begin
      if (_EVAL_765) begin
        _EVAL_1265 <= _EVAL_1089;
      end else if (_EVAL_1188) begin
        _EVAL_1265 <= _EVAL_620;
      end else begin
        _EVAL_1265 <= _EVAL_1089;
      end
    end else begin
      _EVAL_1265 <= _EVAL_1089;
    end
    if (_EVAL_1217) begin
      if (_EVAL_1198) begin
        _EVAL_1266 <= _EVAL_1265;
      end
    end
    _EVAL_1267 <= _EVAL_1156 & _EVAL_685;
    if (_EVAL_776) begin
      if (_EVAL_765) begin
        _EVAL_1268 <= _EVAL_1196;
      end else if (_EVAL_1188) begin
        _EVAL_1268 <= _EVAL_467;
      end else begin
        _EVAL_1268 <= _EVAL_1196;
      end
    end else begin
      _EVAL_1268 <= _EVAL_1196;
    end
    if (_EVAL_1217) begin
      if (_EVAL_684) begin
        _EVAL_1269 <= _EVAL_1329;
      end
    end
    if (_EVAL_1217) begin
      if (_EVAL_567) begin
        _EVAL_1270 <= _EVAL_1265;
      end
    end
    if (_EVAL_1039) begin
      _EVAL_1271 <= _EVAL_1092;
    end
    if (_EVAL_93) begin
      _EVAL_1272 <= 1'h0;
    end else if (_EVAL_776) begin
      if (_EVAL_765) begin
        _EVAL_1272 <= _EVAL_512;
      end else if (_EVAL_690) begin
        _EVAL_1272 <= 1'h0;
      end else begin
        _EVAL_1272 <= _EVAL_512;
      end
    end else begin
      _EVAL_1272 <= _EVAL_512;
    end
    if (_EVAL_93) begin
      _EVAL_1273 <= 6'h0;
    end else if (_EVAL_776) begin
      if (_EVAL_1115) begin
        if (_EVAL_743) begin
          _EVAL_1273 <= _EVAL_343;
        end else begin
          _EVAL_1273 <= 6'h0;
        end
      end else begin
        _EVAL_1273 <= _EVAL_451;
      end
    end
    if (_EVAL_776) begin
      if (!(_EVAL_765)) begin
        if (_EVAL_1188) begin
          _EVAL_1274 <= _EVAL_1190;
        end
      end
    end
    if (_EVAL_1217) begin
      if (_EVAL_684) begin
        _EVAL_1275 <= _EVAL_1302;
      end
    end
    if (_EVAL_1217) begin
      if (_EVAL_629) begin
        _EVAL_1276 <= _EVAL_1329;
      end
    end
    if (_EVAL_651) begin
      _EVAL_1277 <= _EVAL_803;
    end
    if (_EVAL_1039) begin
      _EVAL_1278 <= _EVAL_98;
    end
    if (_EVAL_93) begin
      _EVAL_1279 <= 7'h0;
    end else if (_EVAL_775) begin
      _EVAL_1279 <= 7'h3;
    end else if (_EVAL_254) begin
      _EVAL_1279 <= _EVAL_444;
    end else if (_EVAL_281) begin
      _EVAL_1279 <= _EVAL_1171;
    end
    if (_EVAL_1039) begin
      _EVAL_1280 <= _EVAL_491;
    end
    if (_EVAL_1217) begin
      if (_EVAL_1198) begin
        _EVAL_1281 <= _EVAL_1302;
      end
    end
    if (_EVAL_651) begin
      _EVAL_1282 <= _EVAL_420;
    end
    if (_EVAL_651) begin
      _EVAL_1283 <= _EVAL_1315;
    end
    if (_EVAL_1167) begin
      _EVAL_1284 <= _EVAL_328;
    end
    if (_EVAL_946) begin
      if (_EVAL_492) begin
        _EVAL_1285 <= _EVAL_510;
      end else begin
        _EVAL_1285 <= _EVAL_1212;
      end
    end else begin
      _EVAL_1285 <= _EVAL_1212;
    end
    if (_EVAL_651) begin
      _EVAL_1286 <= _EVAL_353;
    end
    if (_EVAL_1039) begin
      _EVAL_1287 <= _EVAL_98;
    end
    if (_EVAL_1217) begin
      if (_EVAL_487) begin
        _EVAL_1288 <= _EVAL_1302;
      end
    end
    if (_EVAL_1217) begin
      if (_EVAL_629) begin
        _EVAL_1289 <= _EVAL_1265;
      end
    end
    if (_EVAL_1217) begin
      if (_EVAL_567) begin
        _EVAL_1290 <= _EVAL_1302;
      end
    end
    if (_EVAL_1167) begin
      _EVAL_1291 <= _EVAL_821;
    end
    if (_EVAL_616) begin
      _EVAL_1292 <= _EVAL_1278;
    end
    _EVAL_1293 <= ~_EVAL_698;
    if (_EVAL_1217) begin
      if (_EVAL_458) begin
        _EVAL_1294 <= _EVAL_1265;
      end
    end
    if (_EVAL_616) begin
      _EVAL_1295 <= _EVAL_353;
    end
    if (_EVAL_93) begin
      _EVAL_1296 <= 6'h0;
    end else if (_EVAL_1217) begin
      if (_EVAL_1011) begin
        if (_EVAL_1097) begin
          _EVAL_1296 <= _EVAL_354;
        end else begin
          _EVAL_1296 <= 6'h0;
        end
      end else begin
        _EVAL_1296 <= _EVAL_155;
      end
    end
    if (_EVAL_1217) begin
      if (_EVAL_487) begin
        _EVAL_1297 <= _EVAL_1329;
      end
    end
    if (_EVAL_651) begin
      if (_EVAL_416) begin
        _EVAL_1298 <= 2'h3;
      end else begin
        _EVAL_1298 <= 2'h0;
      end
    end
    if (_EVAL_1217) begin
      if (_EVAL_664) begin
        _EVAL_1299 <= _EVAL_1265;
      end
    end
    if (_EVAL_1039) begin
      _EVAL_1300 <= _EVAL_36;
    end
    if (_EVAL_1217) begin
      if (_EVAL_1198) begin
        _EVAL_1301 <= _EVAL_1268;
      end
    end
    if (_EVAL_776) begin
      if (_EVAL_765) begin
        _EVAL_1302 <= _EVAL_1261;
      end else if (_EVAL_1188) begin
        _EVAL_1302 <= _EVAL_406;
      end else begin
        _EVAL_1302 <= _EVAL_1261;
      end
    end else begin
      _EVAL_1302 <= _EVAL_1261;
    end
    if (_EVAL_93) begin
      _EVAL_1303 <= 1'h0;
    end else if (_EVAL_776) begin
      if (_EVAL_765) begin
        _EVAL_1303 <= _EVAL_466;
      end else if (_EVAL_505) begin
        _EVAL_1303 <= 1'h0;
      end else begin
        _EVAL_1303 <= _EVAL_466;
      end
    end else begin
      _EVAL_1303 <= _EVAL_466;
    end
    if (_EVAL_1167) begin
      _EVAL_1304 <= _EVAL_1111;
    end
    if (_EVAL_1167) begin
      _EVAL_1305 <= _EVAL_950;
    end
    if (_EVAL_616) begin
      if (_EVAL_872) begin
        _EVAL_1306 <= _EVAL_6;
      end else begin
        _EVAL_1306 <= _EVAL_1016;
      end
    end
    if (_EVAL_93) begin
      _EVAL_1307 <= 1'h0;
    end else if (_EVAL_776) begin
      if (_EVAL_765) begin
        _EVAL_1307 <= _EVAL_757;
      end else if (_EVAL_593) begin
        _EVAL_1307 <= 1'h0;
      end else begin
        _EVAL_1307 <= _EVAL_757;
      end
    end else begin
      _EVAL_1307 <= _EVAL_757;
    end
    if (_EVAL_1166) begin
      _EVAL_1308 <= _EVAL_617;
    end
    if (_EVAL_1217) begin
      if (_EVAL_664) begin
        _EVAL_1309 <= _EVAL_1268;
      end
    end
    if (_EVAL_1217) begin
      if (_EVAL_629) begin
        _EVAL_1310 <= _EVAL_1302;
      end
    end
    if (_EVAL_1039) begin
      _EVAL_1311 <= _EVAL_1092;
    end
    if (_EVAL_1217) begin
      if (_EVAL_664) begin
        _EVAL_1312 <= _EVAL_1329;
      end
    end
    if (_EVAL_1217) begin
      if (_EVAL_458) begin
        _EVAL_1313 <= _EVAL_1268;
      end
    end
    if (_EVAL_1217) begin
      if (_EVAL_567) begin
        _EVAL_1314 <= _EVAL_1268;
      end
    end
    if (_EVAL_1039) begin
      _EVAL_1315 <= _EVAL_122;
    end
    if (_EVAL_1217) begin
      if (_EVAL_1198) begin
        _EVAL_1316 <= _EVAL_1329;
      end
    end
    if (_EVAL_1039) begin
      _EVAL_1317 <= _EVAL_111;
    end
    if (_EVAL_93) begin
      _EVAL_1318 <= 1'h0;
    end else if (_EVAL_776) begin
      if (_EVAL_765) begin
        _EVAL_1318 <= _EVAL_130;
      end else if (_EVAL_1173) begin
        _EVAL_1318 <= 1'h0;
      end else begin
        _EVAL_1318 <= _EVAL_130;
      end
    end else begin
      _EVAL_1318 <= _EVAL_130;
    end
    if (_EVAL_93) begin
      _EVAL_1319 <= 1'h0;
    end else begin
      _EVAL_1319 <= _EVAL_538;
    end
    if (_EVAL_1039) begin
      _EVAL_1320 <= _EVAL_15;
    end
    if (_EVAL_1217) begin
      if (_EVAL_684) begin
        _EVAL_1321 <= _EVAL_1268;
      end
    end
    if (_EVAL_1217) begin
      if (_EVAL_458) begin
        _EVAL_1322 <= _EVAL_1329;
      end
    end
    if (_EVAL_1217) begin
      if (_EVAL_629) begin
        _EVAL_1323 <= _EVAL_1268;
      end
    end
    if (_EVAL_651) begin
      _EVAL_1324 <= _EVAL_424;
    end
    if (_EVAL_1217) begin
      if (_EVAL_487) begin
        _EVAL_1325 <= _EVAL_1268;
      end
    end
    if (_EVAL_1217) begin
      if (_EVAL_664) begin
        _EVAL_1326 <= _EVAL_1302;
      end
    end
    if (_EVAL_651) begin
      _EVAL_1327 <= _EVAL_172;
    end
    _EVAL_1328 <= _EVAL_25;
    if (_EVAL_776) begin
      if (_EVAL_765) begin
        _EVAL_1329 <= _EVAL_1068;
      end else if (_EVAL_1188) begin
        _EVAL_1329 <= _EVAL_179;
      end else begin
        _EVAL_1329 <= _EVAL_1068;
      end
    end else begin
      _EVAL_1329 <= _EVAL_1068;
    end
    if (_EVAL_93) begin
      _EVAL_1330 <= 1'h0;
    end else if (_EVAL_776) begin
      if (_EVAL_765) begin
        _EVAL_1330 <= _EVAL_979;
      end else if (_EVAL_431) begin
        _EVAL_1330 <= 1'h0;
      end else begin
        _EVAL_1330 <= _EVAL_979;
      end
    end else begin
      _EVAL_1330 <= _EVAL_979;
    end
    if (_EVAL_616) begin
      _EVAL_1331 <= _EVAL_52;
    end
    if (_EVAL_616) begin
      _EVAL_1332 <= _EVAL_570;
    end
    if (_EVAL_93) begin
      _EVAL_1333 <= 1'h0;
    end else begin
      _EVAL_1333 <= _EVAL_203;
    end
    if (_EVAL_651) begin
      _EVAL_1334 <= _EVAL_899;
    end
    if (_EVAL_1167) begin
      _EVAL_1335 <= _EVAL_592;
    end
    if (_EVAL_1039) begin
      _EVAL_1336 <= _EVAL_115;
    end
    if (_EVAL_1217) begin
      if (_EVAL_684) begin
        _EVAL_1337 <= _EVAL_1265;
      end
    end
    if (_EVAL_93) begin
      _EVAL_1338 <= 1'h0;
    end else begin
      _EVAL_1338 <= _EVAL_221;
    end
    if (_EVAL_651) begin
      _EVAL_1339 <= _EVAL_1320;
    end
    _EVAL_1340 <= _EVAL_2;
    if (_EVAL_1039) begin
      _EVAL_1341 <= _EVAL_77;
    end
    if (_EVAL_93) begin
      _EVAL_1342 <= 1'h0;
    end else if (_EVAL_776) begin
      if (_EVAL_765) begin
        _EVAL_1342 <= _EVAL_906;
      end else if (_EVAL_1001) begin
        _EVAL_1342 <= 1'h0;
      end else begin
        _EVAL_1342 <= _EVAL_906;
      end
    end else begin
      _EVAL_1342 <= _EVAL_906;
    end
    if (_EVAL_1167) begin
      _EVAL_1343 <= _EVAL_1295;
    end
    if (_EVAL_1217) begin
      if (_EVAL_458) begin
        _EVAL_1344 <= _EVAL_1302;
      end
    end
    if (_EVAL_651) begin
      _EVAL_1345 <= _EVAL_1336;
    end
    if (_EVAL_93) begin
      _EVAL_1346 <= 3'h0;
    end else if (_EVAL_776) begin
      if (_EVAL_765) begin
        if (_EVAL_539) begin
          _EVAL_1346 <= 3'h7;
        end else begin
          _EVAL_1346 <= _EVAL_792;
        end
      end else begin
        _EVAL_1346 <= _EVAL_792;
      end
    end else begin
      _EVAL_1346 <= _EVAL_792;
    end
    if (_EVAL_93) begin
      _EVAL_1347 <= 1'h0;
    end else begin
      _EVAL_1347 <= _EVAL_198;
    end
    if (_EVAL_1217) begin
      if (_EVAL_487) begin
        _EVAL_1348 <= _EVAL_1265;
      end
    end
    if (_EVAL_1217) begin
      if (_EVAL_567) begin
        _EVAL_1349 <= _EVAL_1329;
      end
    end
    if (_EVAL_93) begin
      _EVAL_1350 <= 1'h0;
    end else if (_EVAL_776) begin
      if (_EVAL_765) begin
        _EVAL_1350 <= _EVAL_511;
      end else if (_EVAL_1210) begin
        _EVAL_1350 <= 1'h0;
      end else begin
        _EVAL_1350 <= _EVAL_511;
      end
    end else begin
      _EVAL_1350 <= _EVAL_511;
    end
    if (_EVAL_776) begin
      if (_EVAL_765) begin
        _EVAL_1351 <= _EVAL_729;
      end else if (_EVAL_1188) begin
        _EVAL_1351 <= 5'h0;
      end else begin
        _EVAL_1351 <= _EVAL_729;
      end
    end else begin
      _EVAL_1351 <= _EVAL_729;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_1160 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_1263 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_1264 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_1265 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_1266 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_1267 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_1268 = _RAND_6[6:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_1269 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_1270 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_1271 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_1272 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_1273 = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_1274 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_1275 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_1276 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_1277 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_1278 = _RAND_16[4:0];
  _RAND_17 = {1{`RANDOM}};
  _EVAL_1279 = _RAND_17[6:0];
  _RAND_18 = {1{`RANDOM}};
  _EVAL_1280 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  _EVAL_1281 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  _EVAL_1282 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _EVAL_1283 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  _EVAL_1284 = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  _EVAL_1285 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  _EVAL_1286 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  _EVAL_1287 = _RAND_25[4:0];
  _RAND_26 = {1{`RANDOM}};
  _EVAL_1288 = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  _EVAL_1289 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  _EVAL_1290 = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  _EVAL_1291 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  _EVAL_1292 = _RAND_30[4:0];
  _RAND_31 = {1{`RANDOM}};
  _EVAL_1293 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  _EVAL_1294 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  _EVAL_1295 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  _EVAL_1296 = _RAND_34[5:0];
  _RAND_35 = {1{`RANDOM}};
  _EVAL_1297 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  _EVAL_1298 = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  _EVAL_1299 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  _EVAL_1300 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  _EVAL_1301 = _RAND_39[6:0];
  _RAND_40 = {1{`RANDOM}};
  _EVAL_1302 = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  _EVAL_1303 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  _EVAL_1304 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  _EVAL_1305 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  _EVAL_1306 = _RAND_44[3:0];
  _RAND_45 = {1{`RANDOM}};
  _EVAL_1307 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  _EVAL_1308 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  _EVAL_1309 = _RAND_47[6:0];
  _RAND_48 = {1{`RANDOM}};
  _EVAL_1310 = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  _EVAL_1311 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  _EVAL_1312 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  _EVAL_1313 = _RAND_51[6:0];
  _RAND_52 = {1{`RANDOM}};
  _EVAL_1314 = _RAND_52[6:0];
  _RAND_53 = {1{`RANDOM}};
  _EVAL_1315 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  _EVAL_1316 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  _EVAL_1317 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  _EVAL_1318 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  _EVAL_1319 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  _EVAL_1320 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  _EVAL_1321 = _RAND_59[6:0];
  _RAND_60 = {1{`RANDOM}};
  _EVAL_1322 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  _EVAL_1323 = _RAND_61[6:0];
  _RAND_62 = {1{`RANDOM}};
  _EVAL_1324 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  _EVAL_1325 = _RAND_63[6:0];
  _RAND_64 = {1{`RANDOM}};
  _EVAL_1326 = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  _EVAL_1327 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  _EVAL_1328 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  _EVAL_1329 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  _EVAL_1330 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  _EVAL_1331 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  _EVAL_1332 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  _EVAL_1333 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  _EVAL_1334 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  _EVAL_1335 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  _EVAL_1336 = _RAND_74[3:0];
  _RAND_75 = {1{`RANDOM}};
  _EVAL_1337 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  _EVAL_1338 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  _EVAL_1339 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  _EVAL_1340 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  _EVAL_1341 = _RAND_79[6:0];
  _RAND_80 = {1{`RANDOM}};
  _EVAL_1342 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  _EVAL_1343 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  _EVAL_1344 = _RAND_82[1:0];
  _RAND_83 = {1{`RANDOM}};
  _EVAL_1345 = _RAND_83[3:0];
  _RAND_84 = {1{`RANDOM}};
  _EVAL_1346 = _RAND_84[2:0];
  _RAND_85 = {1{`RANDOM}};
  _EVAL_1347 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  _EVAL_1348 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  _EVAL_1349 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  _EVAL_1350 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  _EVAL_1351 = _RAND_89[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
