//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_20(
  input         _EVAL,
  output [1:0]  _EVAL_0,
  output        _EVAL_1,
  output        _EVAL_2,
  input  [3:0]  _EVAL_3,
  output [31:0] _EVAL_4,
  output        _EVAL_5,
  input  [31:0] _EVAL_6,
  output        _EVAL_7,
  input         _EVAL_8,
  input  [2:0]  _EVAL_9,
  input         _EVAL_10,
  output [2:0]  _EVAL_11,
  output [2:0]  _EVAL_12,
  input  [2:0]  _EVAL_13,
  input         _EVAL_14,
  output [1:0]  _EVAL_15,
  output [4:0]  _EVAL_16,
  output [2:0]  _EVAL_17,
  input         _EVAL_18,
  input  [2:0]  _EVAL_19,
  input         _EVAL_20,
  input         _EVAL_21,
  output        _EVAL_22,
  input         _EVAL_23,
  output        _EVAL_24,
  output [3:0]  _EVAL_25,
  input         _EVAL_26,
  output [2:0]  _EVAL_27,
  input  [4:0]  _EVAL_28,
  input  [31:0] _EVAL_29,
  input  [30:0] _EVAL_30,
  input         _EVAL_31,
  input         _EVAL_32,
  output [30:0] _EVAL_33,
  output [31:0] _EVAL_34
);
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire [3:0] _EVAL_37;
  wire [2:0] _EVAL_38;
  wire [2:0] _EVAL_39;
  wire [31:0] _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire [4:0] buffer__EVAL;
  wire [30:0] buffer__EVAL_0;
  wire [2:0] buffer__EVAL_1;
  wire [2:0] buffer__EVAL_2;
  wire [31:0] buffer__EVAL_3;
  wire [31:0] buffer__EVAL_4;
  wire  buffer__EVAL_5;
  wire [2:0] buffer__EVAL_6;
  wire  buffer__EVAL_7;
  wire [30:0] buffer__EVAL_8;
  wire [2:0] buffer__EVAL_9;
  wire  buffer__EVAL_10;
  wire  buffer__EVAL_11;
  wire [2:0] buffer__EVAL_12;
  wire [4:0] buffer__EVAL_13;
  wire [31:0] buffer__EVAL_14;
  wire [2:0] buffer__EVAL_15;
  wire [2:0] buffer__EVAL_16;
  wire  buffer__EVAL_17;
  wire  buffer__EVAL_18;
  wire [4:0] buffer__EVAL_19;
  wire  buffer__EVAL_20;
  wire  buffer__EVAL_21;
  wire  buffer__EVAL_22;
  wire  buffer__EVAL_23;
  wire  buffer__EVAL_24;
  wire [3:0] buffer__EVAL_25;
  wire  buffer__EVAL_26;
  wire  buffer__EVAL_27;
  wire [1:0] buffer__EVAL_28;
  wire  buffer__EVAL_29;
  wire  buffer__EVAL_30;
  wire [2:0] buffer__EVAL_31;
  wire  buffer__EVAL_32;
  wire  buffer__EVAL_33;
  wire  buffer__EVAL_34;
  wire  buffer__EVAL_35;
  wire  buffer__EVAL_36;
  wire [4:0] buffer__EVAL_37;
  wire  buffer__EVAL_38;
  wire  buffer__EVAL_39;
  wire [1:0] buffer__EVAL_40;
  wire [2:0] buffer__EVAL_41;
  wire [2:0] buffer__EVAL_42;
  wire [31:0] buffer__EVAL_43;
  wire [3:0] buffer__EVAL_44;
  wire  buffer__EVAL_45;
  wire  buffer__EVAL_46;
  wire  buffer__EVAL_47;
  wire  buffer__EVAL_48;
  wire [4:0] _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire [3:0] _EVAL_47;
  wire [3:0] _EVAL_48;
  wire [2:0] _EVAL_49;
  wire  _EVAL_50;
  wire [1:0] _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire [2:0] _EVAL_55;
  wire  _EVAL_56;
  wire [2:0] _EVAL_57;
  wire  _EVAL_58;
  wire [2:0] _EVAL_59;
  wire  _EVAL_60;
  wire [2:0] _EVAL_61;
  wire [1:0] _EVAL_62;
  wire [2:0] _EVAL_63;
  wire [2:0] _EVAL_64;
  wire  _EVAL_65;
  wire [4:0] _EVAL_66;
  wire [30:0] _EVAL_67;
  wire [30:0] _EVAL_68;
  wire [2:0] _EVAL_69;
  wire [30:0] _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire [4:0] _EVAL_73;
  wire  _EVAL_74;
  wire [31:0] _EVAL_75;
  wire [2:0] _EVAL_76;
  wire [2:0] _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire [31:0] _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire [2:0] _EVAL_84;
  wire [31:0] _EVAL_85;
  wire [2:0] _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire [31:0] _EVAL_89;
  wire  _EVAL_90;
  wire [2:0] _EVAL_91;
  wire [31:0] _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire [2:0] _EVAL_95;
  wire  _EVAL_96;
  wire [2:0] _EVAL_97;
  wire [4:0] _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire [31:0] _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire [30:0] _EVAL_108;
  wire  _EVAL_109;
  wire [2:0] _EVAL_110;
  wire  tl2ahb__EVAL;
  wire  tl2ahb__EVAL_0;
  wire [30:0] tl2ahb__EVAL_1;
  wire  tl2ahb__EVAL_2;
  wire  tl2ahb__EVAL_3;
  wire [2:0] tl2ahb__EVAL_4;
  wire  tl2ahb__EVAL_5;
  wire [1:0] tl2ahb__EVAL_6;
  wire [3:0] tl2ahb__EVAL_7;
  wire  tl2ahb__EVAL_8;
  wire [31:0] tl2ahb__EVAL_9;
  wire  tl2ahb__EVAL_10;
  wire [31:0] tl2ahb__EVAL_11;
  wire  tl2ahb__EVAL_12;
  wire  tl2ahb__EVAL_13;
  wire [2:0] tl2ahb__EVAL_14;
  wire [2:0] tl2ahb__EVAL_15;
  wire  tl2ahb__EVAL_16;
  wire [3:0] tl2ahb__EVAL_17;
  wire [2:0] tl2ahb__EVAL_18;
  wire  tl2ahb__EVAL_19;
  wire [2:0] tl2ahb__EVAL_20;
  wire [2:0] tl2ahb__EVAL_21;
  wire [31:0] tl2ahb__EVAL_22;
  wire [4:0] tl2ahb__EVAL_23;
  wire  tl2ahb__EVAL_24;
  wire [30:0] tl2ahb__EVAL_25;
  wire  tl2ahb__EVAL_26;
  wire  tl2ahb__EVAL_27;
  wire  tl2ahb__EVAL_28;
  wire  tl2ahb__EVAL_29;
  wire [31:0] tl2ahb__EVAL_30;
  wire [1:0] tl2ahb__EVAL_31;
  wire  tl2ahb__EVAL_32;
  wire [2:0] tl2ahb__EVAL_33;
  wire [4:0] tl2ahb__EVAL_34;
  wire  _EVAL_111;
  wire [31:0] _EVAL_112;
  wire [2:0] _EVAL_113;
  wire  _EVAL_114;
  wire [1:0] _EVAL_115;
  wire [2:0] _EVAL_116;
  wire [3:0] _EVAL_117;
  wire  _EVAL_118;
  wire [4:0] _EVAL_119;
  wire  _EVAL_120;
  wire [2:0] _EVAL_121;
  wire [2:0] _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire [30:0] _EVAL_127;
  wire [31:0] _EVAL_128;
  wire [4:0] _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire [2:0] _EVAL_132;
  wire [1:0] _EVAL_133;
  wire [3:0] _EVAL_134;
  wire [1:0] _EVAL_135;
  wire [31:0] _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire [2:0] _EVAL_139;
  wire  _EVAL_140;
  wire [4:0] _EVAL_141;
  wire [4:0] _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire [4:0] _EVAL_145;
  wire [2:0] _EVAL_146;
  wire [4:0] _EVAL_147;
  wire  _EVAL_148;
  wire [2:0] _EVAL_149;
  wire [2:0] _EVAL_150;
  wire  _EVAL_151;
  wire [2:0] _EVAL_152;
  wire  _EVAL_153;
  wire [4:0] _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire [4:0] _EVAL_157;
  wire [31:0] _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire [1:0] _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire [2:0] _EVAL_166;
  wire [3:0] _EVAL_167;
  wire [2:0] _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire [31:0] _EVAL_177;
  wire [30:0] _EVAL_178;
  _EVAL_19 buffer (
    ._EVAL(buffer__EVAL),
    ._EVAL_0(buffer__EVAL_0),
    ._EVAL_1(buffer__EVAL_1),
    ._EVAL_2(buffer__EVAL_2),
    ._EVAL_3(buffer__EVAL_3),
    ._EVAL_4(buffer__EVAL_4),
    ._EVAL_5(buffer__EVAL_5),
    ._EVAL_6(buffer__EVAL_6),
    ._EVAL_7(buffer__EVAL_7),
    ._EVAL_8(buffer__EVAL_8),
    ._EVAL_9(buffer__EVAL_9),
    ._EVAL_10(buffer__EVAL_10),
    ._EVAL_11(buffer__EVAL_11),
    ._EVAL_12(buffer__EVAL_12),
    ._EVAL_13(buffer__EVAL_13),
    ._EVAL_14(buffer__EVAL_14),
    ._EVAL_15(buffer__EVAL_15),
    ._EVAL_16(buffer__EVAL_16),
    ._EVAL_17(buffer__EVAL_17),
    ._EVAL_18(buffer__EVAL_18),
    ._EVAL_19(buffer__EVAL_19),
    ._EVAL_20(buffer__EVAL_20),
    ._EVAL_21(buffer__EVAL_21),
    ._EVAL_22(buffer__EVAL_22),
    ._EVAL_23(buffer__EVAL_23),
    ._EVAL_24(buffer__EVAL_24),
    ._EVAL_25(buffer__EVAL_25),
    ._EVAL_26(buffer__EVAL_26),
    ._EVAL_27(buffer__EVAL_27),
    ._EVAL_28(buffer__EVAL_28),
    ._EVAL_29(buffer__EVAL_29),
    ._EVAL_30(buffer__EVAL_30),
    ._EVAL_31(buffer__EVAL_31),
    ._EVAL_32(buffer__EVAL_32),
    ._EVAL_33(buffer__EVAL_33),
    ._EVAL_34(buffer__EVAL_34),
    ._EVAL_35(buffer__EVAL_35),
    ._EVAL_36(buffer__EVAL_36),
    ._EVAL_37(buffer__EVAL_37),
    ._EVAL_38(buffer__EVAL_38),
    ._EVAL_39(buffer__EVAL_39),
    ._EVAL_40(buffer__EVAL_40),
    ._EVAL_41(buffer__EVAL_41),
    ._EVAL_42(buffer__EVAL_42),
    ._EVAL_43(buffer__EVAL_43),
    ._EVAL_44(buffer__EVAL_44),
    ._EVAL_45(buffer__EVAL_45),
    ._EVAL_46(buffer__EVAL_46),
    ._EVAL_47(buffer__EVAL_47),
    ._EVAL_48(buffer__EVAL_48)
  );
  _EVAL_15 tl2ahb (
    ._EVAL(tl2ahb__EVAL),
    ._EVAL_0(tl2ahb__EVAL_0),
    ._EVAL_1(tl2ahb__EVAL_1),
    ._EVAL_2(tl2ahb__EVAL_2),
    ._EVAL_3(tl2ahb__EVAL_3),
    ._EVAL_4(tl2ahb__EVAL_4),
    ._EVAL_5(tl2ahb__EVAL_5),
    ._EVAL_6(tl2ahb__EVAL_6),
    ._EVAL_7(tl2ahb__EVAL_7),
    ._EVAL_8(tl2ahb__EVAL_8),
    ._EVAL_9(tl2ahb__EVAL_9),
    ._EVAL_10(tl2ahb__EVAL_10),
    ._EVAL_11(tl2ahb__EVAL_11),
    ._EVAL_12(tl2ahb__EVAL_12),
    ._EVAL_13(tl2ahb__EVAL_13),
    ._EVAL_14(tl2ahb__EVAL_14),
    ._EVAL_15(tl2ahb__EVAL_15),
    ._EVAL_16(tl2ahb__EVAL_16),
    ._EVAL_17(tl2ahb__EVAL_17),
    ._EVAL_18(tl2ahb__EVAL_18),
    ._EVAL_19(tl2ahb__EVAL_19),
    ._EVAL_20(tl2ahb__EVAL_20),
    ._EVAL_21(tl2ahb__EVAL_21),
    ._EVAL_22(tl2ahb__EVAL_22),
    ._EVAL_23(tl2ahb__EVAL_23),
    ._EVAL_24(tl2ahb__EVAL_24),
    ._EVAL_25(tl2ahb__EVAL_25),
    ._EVAL_26(tl2ahb__EVAL_26),
    ._EVAL_27(tl2ahb__EVAL_27),
    ._EVAL_28(tl2ahb__EVAL_28),
    ._EVAL_29(tl2ahb__EVAL_29),
    ._EVAL_30(tl2ahb__EVAL_30),
    ._EVAL_31(tl2ahb__EVAL_31),
    ._EVAL_32(tl2ahb__EVAL_32),
    ._EVAL_33(tl2ahb__EVAL_33),
    ._EVAL_34(tl2ahb__EVAL_34)
  );
  assign buffer__EVAL_14 = tl2ahb__EVAL_22;
  assign _EVAL_48 = _EVAL_167;
  assign _EVAL_7 = tl2ahb__EVAL_5;
  assign _EVAL_62 = _EVAL_162;
  assign _EVAL_154 = _EVAL_129;
  assign _EVAL_46 = _EVAL_100;
  assign _EVAL_160 = _EVAL_118;
  assign _EVAL_67 = _EVAL_178;
  assign _EVAL_36 = _EVAL_155;
  assign _EVAL_40 = _EVAL_112;
  assign _EVAL_128 = buffer__EVAL_43;
  assign _EVAL_86 = _EVAL_76;
  assign buffer__EVAL_11 = _EVAL_105;
  assign buffer__EVAL_21 = _EVAL_65;
  assign _EVAL_125 = _EVAL_130;
  assign _EVAL_119 = _EVAL_145;
  assign buffer__EVAL_39 = _EVAL_148;
  assign buffer__EVAL_45 = _EVAL_170;
  assign buffer__EVAL_26 = _EVAL_44;
  assign _EVAL_136 = _EVAL_102;
  assign _EVAL_27 = tl2ahb__EVAL_18;
  assign _EVAL_135 = buffer__EVAL_28;
  assign _EVAL_170 = _EVAL_144;
  assign _EVAL_150 = _EVAL_77;
  assign _EVAL_123 = _EVAL_23;
  assign _EVAL_131 = _EVAL_54;
  assign _EVAL_49 = _EVAL_132;
  assign _EVAL_11 = tl2ahb__EVAL_33;
  assign _EVAL_142 = buffer__EVAL;
  assign _EVAL_178 = _EVAL_30;
  assign _EVAL_144 = _EVAL_171;
  assign _EVAL_33 = tl2ahb__EVAL_25;
  assign _EVAL_45 = _EVAL_72;
  assign _EVAL_58 = _EVAL_41;
  assign _EVAL_109 = _EVAL_90;
  assign _EVAL_0 = tl2ahb__EVAL_6;
  assign _EVAL_41 = buffer__EVAL_7;
  assign _EVAL_153 = _EVAL_120;
  assign _EVAL_105 = _EVAL_35;
  assign _EVAL_130 = _EVAL_159;
  assign buffer__EVAL_22 = _EVAL_14;
  assign _EVAL_162 = _EVAL_115;
  assign _EVAL_75 = _EVAL_85;
  assign _EVAL_82 = _EVAL_137;
  assign _EVAL_72 = _EVAL_36;
  assign _EVAL_53 = _EVAL;
  assign _EVAL_145 = _EVAL_157;
  assign _EVAL_122 = _EVAL_86;
  assign _EVAL_89 = _EVAL_128;
  assign _EVAL_121 = _EVAL_146;
  assign _EVAL_146 = _EVAL_97;
  assign _EVAL_124 = _EVAL_123;
  assign _EVAL_159 = _EVAL_131;
  assign _EVAL_103 = _EVAL_176;
  assign _EVAL_117 = _EVAL_3;
  assign _EVAL_24 = _EVAL_52;
  assign _EVAL_152 = buffer__EVAL_6;
  assign buffer__EVAL_46 = _EVAL_32;
  assign tl2ahb__EVAL_3 = buffer__EVAL_35;
  assign _EVAL_143 = _EVAL_78;
  assign tl2ahb__EVAL_32 = buffer__EVAL_5;
  assign _EVAL_52 = _EVAL_153;
  assign tl2ahb__EVAL_29 = buffer__EVAL_18;
  assign _EVAL_17 = _EVAL_39;
  assign _EVAL_101 = _EVAL_53;
  assign _EVAL_84 = _EVAL_168;
  assign _EVAL_63 = _EVAL_13;
  assign buffer__EVAL_3 = _EVAL_75;
  assign tl2ahb__EVAL_28 = _EVAL_32;
  assign _EVAL_175 = _EVAL_163;
  assign _EVAL_127 = _EVAL_108;
  assign _EVAL_167 = _EVAL_37;
  assign _EVAL_151 = _EVAL_88;
  assign tl2ahb__EVAL_30 = buffer__EVAL_4;
  assign _EVAL_111 = _EVAL_160;
  assign _EVAL_22 = _EVAL_93;
  assign tl2ahb__EVAL_20 = buffer__EVAL_42;
  assign tl2ahb__EVAL_27 = _EVAL_10;
  assign _EVAL_94 = _EVAL_101;
  assign _EVAL_133 = _EVAL_62;
  assign _EVAL_50 = _EVAL_106;
  assign _EVAL_1 = _EVAL_109;
  assign _EVAL_80 = _EVAL_124;
  assign buffer__EVAL_0 = _EVAL_70;
  assign tl2ahb__EVAL_9 = _EVAL_29;
  assign _EVAL_155 = buffer__EVAL_24;
  assign buffer__EVAL_34 = tl2ahb__EVAL_0;
  assign buffer__EVAL_1 = _EVAL_55;
  assign _EVAL_138 = _EVAL_172;
  assign _EVAL_134 = _EVAL_48;
  assign _EVAL_37 = _EVAL_47;
  assign _EVAL_76 = _EVAL_113;
  assign _EVAL_129 = _EVAL_28;
  assign _EVAL_42 = _EVAL_18;
  assign _EVAL_174 = _EVAL_80;
  assign _EVAL_66 = _EVAL_98;
  assign _EVAL_35 = _EVAL_156;
  assign buffer__EVAL_12 = tl2ahb__EVAL_4;
  assign _EVAL_140 = _EVAL_82;
  assign _EVAL_81 = _EVAL_92;
  assign _EVAL_115 = _EVAL_135;
  assign buffer__EVAL_17 = tl2ahb__EVAL_24;
  assign _EVAL_5 = _EVAL_96;
  assign _EVAL_44 = _EVAL_99;
  assign _EVAL_176 = _EVAL_143;
  assign _EVAL_97 = _EVAL_149;
  assign _EVAL_79 = _EVAL_45;
  assign _EVAL_4 = tl2ahb__EVAL_11;
  assign _EVAL_87 = _EVAL_26;
  assign buffer__EVAL_10 = tl2ahb__EVAL_19;
  assign buffer__EVAL_40 = tl2ahb__EVAL_31;
  assign _EVAL_99 = _EVAL_174;
  assign tl2ahb__EVAL_10 = _EVAL_14;
  assign tl2ahb__EVAL_17 = buffer__EVAL_44;
  assign tl2ahb__EVAL_13 = buffer__EVAL_29;
  assign buffer__EVAL_25 = _EVAL_134;
  assign buffer__EVAL_13 = tl2ahb__EVAL_34;
  assign _EVAL_148 = _EVAL_125;
  assign buffer__EVAL_32 = _EVAL_83;
  assign tl2ahb__EVAL = buffer__EVAL_48;
  assign _EVAL_68 = _EVAL_67;
  assign _EVAL_164 = _EVAL_60;
  assign _EVAL_165 = _EVAL_74;
  assign _EVAL_60 = buffer__EVAL_47;
  assign _EVAL_158 = _EVAL_89;
  assign _EVAL_69 = _EVAL_63;
  assign buffer__EVAL_19 = _EVAL_43;
  assign _EVAL_106 = _EVAL_175;
  assign _EVAL_65 = _EVAL_126;
  assign _EVAL_78 = _EVAL_31;
  assign _EVAL_92 = _EVAL_40;
  assign tl2ahb__EVAL_2 = buffer__EVAL_38;
  assign _EVAL_61 = _EVAL_64;
  assign _EVAL_43 = _EVAL_119;
  assign tl2ahb__EVAL_16 = _EVAL_8;
  assign _EVAL_59 = _EVAL_121;
  assign _EVAL_77 = _EVAL_139;
  assign buffer__EVAL_23 = _EVAL_114;
  assign _EVAL_114 = _EVAL_56;
  assign _EVAL_112 = _EVAL_6;
  assign _EVAL_116 = _EVAL_110;
  assign _EVAL_139 = _EVAL_116;
  assign _EVAL_73 = _EVAL_142;
  assign _EVAL_132 = _EVAL_84;
  assign _EVAL_57 = _EVAL_38;
  assign buffer__EVAL_30 = tl2ahb__EVAL_26;
  assign _EVAL_15 = _EVAL_51;
  assign _EVAL_85 = _EVAL_81;
  assign tl2ahb__EVAL_21 = buffer__EVAL_16;
  assign _EVAL_16 = _EVAL_66;
  assign _EVAL_2 = _EVAL_138;
  assign _EVAL_177 = _EVAL_136;
  assign _EVAL_55 = _EVAL_59;
  assign tl2ahb__EVAL_23 = buffer__EVAL_37;
  assign _EVAL_102 = _EVAL_158;
  assign _EVAL_88 = _EVAL_42;
  assign _EVAL_173 = _EVAL_20;
  assign _EVAL_107 = _EVAL_140;
  assign _EVAL_161 = _EVAL_164;
  assign _EVAL_64 = _EVAL_57;
  assign tl2ahb__EVAL_8 = buffer__EVAL_20;
  assign _EVAL_104 = _EVAL_173;
  assign _EVAL_38 = _EVAL_69;
  assign _EVAL_149 = _EVAL_19;
  assign _EVAL_71 = _EVAL_104;
  assign _EVAL_83 = _EVAL_46;
  assign _EVAL_95 = _EVAL_122;
  assign _EVAL_108 = _EVAL_68;
  assign tl2ahb__EVAL_1 = buffer__EVAL_8;
  assign _EVAL_98 = _EVAL_147;
  assign _EVAL_90 = _EVAL_107;
  assign _EVAL_163 = buffer__EVAL_36;
  assign _EVAL_166 = _EVAL_95;
  assign _EVAL_168 = _EVAL_152;
  assign _EVAL_93 = _EVAL_79;
  assign _EVAL_56 = _EVAL_169;
  assign _EVAL_172 = _EVAL_50;
  assign _EVAL_12 = _EVAL_91;
  assign _EVAL_141 = _EVAL_73;
  assign _EVAL_47 = _EVAL_117;
  assign buffer__EVAL_2 = _EVAL_166;
  assign _EVAL_51 = _EVAL_133;
  assign _EVAL_74 = _EVAL_87;
  assign buffer__EVAL_33 = tl2ahb__EVAL_12;
  assign _EVAL_120 = _EVAL_161;
  assign _EVAL_96 = _EVAL_111;
  assign _EVAL_118 = _EVAL_58;
  assign buffer__EVAL_31 = tl2ahb__EVAL_14;
  assign _EVAL_156 = _EVAL_94;
  assign tl2ahb__EVAL_15 = buffer__EVAL_15;
  assign _EVAL_100 = _EVAL_71;
  assign _EVAL_147 = _EVAL_141;
  assign buffer__EVAL_41 = _EVAL_61;
  assign _EVAL_171 = _EVAL_151;
  assign _EVAL_54 = _EVAL_21;
  assign _EVAL_34 = _EVAL_177;
  assign _EVAL_169 = _EVAL_165;
  assign _EVAL_137 = buffer__EVAL_27;
  assign _EVAL_70 = _EVAL_127;
  assign _EVAL_39 = _EVAL_49;
  assign _EVAL_25 = tl2ahb__EVAL_7;
  assign _EVAL_91 = _EVAL_150;
  assign _EVAL_110 = buffer__EVAL_9;
  assign _EVAL_157 = _EVAL_154;
  assign _EVAL_113 = _EVAL_9;
  assign _EVAL_126 = _EVAL_103;
endmodule
