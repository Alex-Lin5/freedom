//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_21(
  output        _EVAL,
  input  [4:0]  _EVAL_0,
  input  [31:0] _EVAL_1,
  input         _EVAL_2,
  output [30:0] _EVAL_3,
  output [2:0]  _EVAL_4,
  input  [2:0]  _EVAL_5,
  input  [31:0] _EVAL_6,
  output        _EVAL_7,
  output        _EVAL_8,
  output        _EVAL_9,
  input  [30:0] _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input  [2:0]  _EVAL_15,
  input         _EVAL_16,
  output [4:0]  _EVAL_17,
  output [1:0]  _EVAL_18,
  input         _EVAL_19,
  output [2:0]  _EVAL_20,
  input         _EVAL_21,
  input  [3:0]  _EVAL_22,
  output [1:0]  _EVAL_23,
  input         _EVAL_24,
  input         _EVAL_25,
  output [3:0]  _EVAL_26,
  output [31:0] _EVAL_27,
  output [2:0]  _EVAL_28,
  output        _EVAL_29,
  output [2:0]  _EVAL_30,
  output        _EVAL_31,
  input         _EVAL_32,
  output [31:0] _EVAL_33,
  input         _EVAL_34
);
  wire  bridge_for_ahb_sys_port__EVAL;
  wire [1:0] bridge_for_ahb_sys_port__EVAL_0;
  wire  bridge_for_ahb_sys_port__EVAL_1;
  wire  bridge_for_ahb_sys_port__EVAL_2;
  wire [3:0] bridge_for_ahb_sys_port__EVAL_3;
  wire [31:0] bridge_for_ahb_sys_port__EVAL_4;
  wire  bridge_for_ahb_sys_port__EVAL_5;
  wire [31:0] bridge_for_ahb_sys_port__EVAL_6;
  wire  bridge_for_ahb_sys_port__EVAL_7;
  wire  bridge_for_ahb_sys_port__EVAL_8;
  wire [2:0] bridge_for_ahb_sys_port__EVAL_9;
  wire  bridge_for_ahb_sys_port__EVAL_10;
  wire [2:0] bridge_for_ahb_sys_port__EVAL_11;
  wire [2:0] bridge_for_ahb_sys_port__EVAL_12;
  wire [2:0] bridge_for_ahb_sys_port__EVAL_13;
  wire  bridge_for_ahb_sys_port__EVAL_14;
  wire [1:0] bridge_for_ahb_sys_port__EVAL_15;
  wire [4:0] bridge_for_ahb_sys_port__EVAL_16;
  wire [2:0] bridge_for_ahb_sys_port__EVAL_17;
  wire  bridge_for_ahb_sys_port__EVAL_18;
  wire [2:0] bridge_for_ahb_sys_port__EVAL_19;
  wire  bridge_for_ahb_sys_port__EVAL_20;
  wire  bridge_for_ahb_sys_port__EVAL_21;
  wire  bridge_for_ahb_sys_port__EVAL_22;
  wire  bridge_for_ahb_sys_port__EVAL_23;
  wire  bridge_for_ahb_sys_port__EVAL_24;
  wire [3:0] bridge_for_ahb_sys_port__EVAL_25;
  wire  bridge_for_ahb_sys_port__EVAL_26;
  wire [2:0] bridge_for_ahb_sys_port__EVAL_27;
  wire [4:0] bridge_for_ahb_sys_port__EVAL_28;
  wire [31:0] bridge_for_ahb_sys_port__EVAL_29;
  wire [30:0] bridge_for_ahb_sys_port__EVAL_30;
  wire  bridge_for_ahb_sys_port__EVAL_31;
  wire  bridge_for_ahb_sys_port__EVAL_32;
  wire [30:0] bridge_for_ahb_sys_port__EVAL_33;
  wire [31:0] bridge_for_ahb_sys_port__EVAL_34;
  _EVAL_20 bridge_for_ahb_sys_port (
    ._EVAL(bridge_for_ahb_sys_port__EVAL),
    ._EVAL_0(bridge_for_ahb_sys_port__EVAL_0),
    ._EVAL_1(bridge_for_ahb_sys_port__EVAL_1),
    ._EVAL_2(bridge_for_ahb_sys_port__EVAL_2),
    ._EVAL_3(bridge_for_ahb_sys_port__EVAL_3),
    ._EVAL_4(bridge_for_ahb_sys_port__EVAL_4),
    ._EVAL_5(bridge_for_ahb_sys_port__EVAL_5),
    ._EVAL_6(bridge_for_ahb_sys_port__EVAL_6),
    ._EVAL_7(bridge_for_ahb_sys_port__EVAL_7),
    ._EVAL_8(bridge_for_ahb_sys_port__EVAL_8),
    ._EVAL_9(bridge_for_ahb_sys_port__EVAL_9),
    ._EVAL_10(bridge_for_ahb_sys_port__EVAL_10),
    ._EVAL_11(bridge_for_ahb_sys_port__EVAL_11),
    ._EVAL_12(bridge_for_ahb_sys_port__EVAL_12),
    ._EVAL_13(bridge_for_ahb_sys_port__EVAL_13),
    ._EVAL_14(bridge_for_ahb_sys_port__EVAL_14),
    ._EVAL_15(bridge_for_ahb_sys_port__EVAL_15),
    ._EVAL_16(bridge_for_ahb_sys_port__EVAL_16),
    ._EVAL_17(bridge_for_ahb_sys_port__EVAL_17),
    ._EVAL_18(bridge_for_ahb_sys_port__EVAL_18),
    ._EVAL_19(bridge_for_ahb_sys_port__EVAL_19),
    ._EVAL_20(bridge_for_ahb_sys_port__EVAL_20),
    ._EVAL_21(bridge_for_ahb_sys_port__EVAL_21),
    ._EVAL_22(bridge_for_ahb_sys_port__EVAL_22),
    ._EVAL_23(bridge_for_ahb_sys_port__EVAL_23),
    ._EVAL_24(bridge_for_ahb_sys_port__EVAL_24),
    ._EVAL_25(bridge_for_ahb_sys_port__EVAL_25),
    ._EVAL_26(bridge_for_ahb_sys_port__EVAL_26),
    ._EVAL_27(bridge_for_ahb_sys_port__EVAL_27),
    ._EVAL_28(bridge_for_ahb_sys_port__EVAL_28),
    ._EVAL_29(bridge_for_ahb_sys_port__EVAL_29),
    ._EVAL_30(bridge_for_ahb_sys_port__EVAL_30),
    ._EVAL_31(bridge_for_ahb_sys_port__EVAL_31),
    ._EVAL_32(bridge_for_ahb_sys_port__EVAL_32),
    ._EVAL_33(bridge_for_ahb_sys_port__EVAL_33),
    ._EVAL_34(bridge_for_ahb_sys_port__EVAL_34)
  );
  assign bridge_for_ahb_sys_port__EVAL_26 = _EVAL_21;
  assign bridge_for_ahb_sys_port__EVAL_30 = _EVAL_10;
  assign _EVAL_8 = bridge_for_ahb_sys_port__EVAL_2;
  assign bridge_for_ahb_sys_port__EVAL_6 = _EVAL_6;
  assign _EVAL_9 = bridge_for_ahb_sys_port__EVAL_24;
  assign _EVAL_29 = bridge_for_ahb_sys_port__EVAL_22;
  assign _EVAL_23 = bridge_for_ahb_sys_port__EVAL_0;
  assign _EVAL_28 = bridge_for_ahb_sys_port__EVAL_17;
  assign _EVAL_17 = bridge_for_ahb_sys_port__EVAL_16;
  assign _EVAL_7 = bridge_for_ahb_sys_port__EVAL_5;
  assign _EVAL = bridge_for_ahb_sys_port__EVAL_7;
  assign bridge_for_ahb_sys_port__EVAL_29 = _EVAL_1;
  assign bridge_for_ahb_sys_port__EVAL = _EVAL_13;
  assign bridge_for_ahb_sys_port__EVAL_32 = _EVAL_32;
  assign _EVAL_26 = bridge_for_ahb_sys_port__EVAL_25;
  assign _EVAL_18 = bridge_for_ahb_sys_port__EVAL_15;
  assign bridge_for_ahb_sys_port__EVAL_20 = _EVAL_24;
  assign bridge_for_ahb_sys_port__EVAL_23 = _EVAL_14;
  assign bridge_for_ahb_sys_port__EVAL_19 = _EVAL_12;
  assign _EVAL_27 = bridge_for_ahb_sys_port__EVAL_34;
  assign bridge_for_ahb_sys_port__EVAL_18 = _EVAL_2;
  assign bridge_for_ahb_sys_port__EVAL_14 = _EVAL_11;
  assign bridge_for_ahb_sys_port__EVAL_9 = _EVAL_15;
  assign bridge_for_ahb_sys_port__EVAL_13 = _EVAL_5;
  assign _EVAL_3 = bridge_for_ahb_sys_port__EVAL_33;
  assign _EVAL_20 = bridge_for_ahb_sys_port__EVAL_11;
  assign bridge_for_ahb_sys_port__EVAL_28 = _EVAL_0;
  assign bridge_for_ahb_sys_port__EVAL_8 = _EVAL_34;
  assign bridge_for_ahb_sys_port__EVAL_21 = _EVAL_25;
  assign bridge_for_ahb_sys_port__EVAL_10 = _EVAL_19;
  assign bridge_for_ahb_sys_port__EVAL_31 = _EVAL_16;
  assign _EVAL_30 = bridge_for_ahb_sys_port__EVAL_27;
  assign bridge_for_ahb_sys_port__EVAL_3 = _EVAL_22;
  assign _EVAL_31 = bridge_for_ahb_sys_port__EVAL_1;
  assign _EVAL_33 = bridge_for_ahb_sys_port__EVAL_4;
  assign _EVAL_4 = bridge_for_ahb_sys_port__EVAL_12;
endmodule
