//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_2_assert(
  input  [31:0] _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input  [2:0]  _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input  [3:0]  _EVAL_6,
  input  [3:0]  _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input  [3:0]  _EVAL_10,
  input  [1:0]  _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input  [3:0]  _EVAL_14,
  input  [3:0]  _EVAL_15,
  input  [2:0]  _EVAL_16,
  input         _EVAL_17,
  input  [2:0]  _EVAL_18
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_19;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire [32:0] _EVAL_25;
  wire  _EVAL_26;
  wire [5:0] _EVAL_27;
  wire  _EVAL_28;
  wire [31:0] _EVAL_29;
  wire [31:0] _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire [32:0] _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_36;
  wire [2:0] _EVAL_37;
  wire [32:0] _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire [3:0] _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire [32:0] _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire [8:0] _EVAL_66;
  wire [5:0] _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire [31:0] _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire [8:0] _EVAL_77;
  wire  _EVAL_78;
  wire [1:0] _EVAL_79;
  wire  _EVAL_80;
  wire [7:0] _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire [6:0] _EVAL_84;
  wire [32:0] _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire [7:0] _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire [22:0] _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire [32:0] _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  reg [3:0] _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire [32:0] _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  reg [5:0] _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire [32:0] _EVAL_118;
  wire [32:0] _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire [7:0] _EVAL_122;
  reg [3:0] _EVAL_123;
  wire [32:0] _EVAL_124;
  wire  _EVAL_125;
  wire [15:0] _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire [3:0] _EVAL_129;
  reg [5:0] _EVAL_130;
  wire [1:0] _EVAL_131;
  wire  _EVAL_132;
  wire [31:0] _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire [32:0] _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire [5:0] _EVAL_149;
  wire [5:0] _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire [32:0] _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire [31:0] _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  reg [2:0] _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire [3:0] _EVAL_179;
  wire [32:0] _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire [31:0] _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire [32:0] _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire [32:0] _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire [32:0] _EVAL_210;
  reg [2:0] _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  reg [8:0] _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire [15:0] _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire [32:0] _EVAL_238;
  wire [32:0] _EVAL_239;
  reg [5:0] _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  reg [1:0] _EVAL_243;
  wire  _EVAL_244;
  wire [31:0] _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  reg  _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire [15:0] _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire [8:0] _EVAL_263;
  wire [31:0] _EVAL_264;
  reg [5:0] _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire [5:0] _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire [8:0] _EVAL_278;
  wire  _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  reg [3:0] _EVAL_283;
  wire  _EVAL_284;
  wire [31:0] _EVAL_285;
  wire [8:0] _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire [6:0] _EVAL_291;
  wire  _EVAL_292;
  wire [22:0] _EVAL_293;
  wire  _EVAL_294;
  wire  _EVAL_295;
  reg  _EVAL_296;
  wire [32:0] _EVAL_297;
  reg [3:0] _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire [32:0] _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_307;
  wire  _EVAL_308;
  wire  _EVAL_309;
  wire [32:0] _EVAL_310;
  wire  _EVAL_311;
  wire [6:0] _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_314;
  reg [31:0] _EVAL_315;
  wire [6:0] _EVAL_316;
  wire  _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_320;
  wire [2:0] _EVAL_321;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_322;
  wire  _EVAL_323;
  reg [2:0] _EVAL_324;
  wire  _EVAL_326;
  wire [32:0] _EVAL_327;
  wire  _EVAL_328;
  wire  _EVAL_329;
  wire  _EVAL_330;
  wire [32:0] _EVAL_331;
  wire [3:0] _EVAL_332;
  wire  _EVAL_333;
  wire  _EVAL_334;
  wire  _EVAL_335;
  wire  _EVAL_336;
  wire [7:0] _EVAL_337;
  wire  _EVAL_338;
  wire [32:0] _EVAL_339;
  wire  _EVAL_340;
  wire  _EVAL_341;
  wire  _EVAL_342;
  wire [31:0] _EVAL_343;
  wire [32:0] _EVAL_344;
  wire  _EVAL_345;
  reg [31:0] _EVAL_346;
  wire  _EVAL_347;
  wire [15:0] _EVAL_349;
  wire  _EVAL_350;
  wire [8:0] _EVAL_351;
  wire  _EVAL_352;
  wire [8:0] _EVAL_353;
  wire [8:0] _EVAL_354;
  wire  _EVAL_355;
  wire  _EVAL_356;
  wire  _EVAL_358;
  wire  _EVAL_359;
  wire  _EVAL_360;
  wire  _EVAL_361;
  wire  _EVAL_362;
  wire [5:0] _EVAL_363;
  wire  _EVAL_364;
  wire  _EVAL_365;
  wire  _EVAL_366;
  wire  _EVAL_367;
  wire  _EVAL_368;
  wire  _EVAL_369;
  wire  _EVAL_370;
  wire  _EVAL_371;
  wire  _EVAL_372;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_173 = _EVAL_168 & _EVAL_71;
  assign _EVAL_187 = _EVAL_2 & _EVAL_13;
  assign _EVAL_206 = $signed(_EVAL_210) & -33'sh1000;
  assign _EVAL_195 = ~_EVAL_31;
  assign _EVAL_138 = $signed(_EVAL_57) & -33'sh5000;
  assign _EVAL_219 = _EVAL_45 & _EVAL_74;
  assign _EVAL_152 = _EVAL_1 & _EVAL_365;
  assign _EVAL_233 = ~_EVAL_248;
  assign _EVAL_288 = _EVAL_371 | _EVAL_202;
  assign _EVAL_139 = _EVAL_45 & _EVAL_359;
  assign _EVAL_316 = _EVAL_240 - 6'h1;
  assign _EVAL_210 = {1'b0,$signed(_EVAL_161)};
  assign _EVAL_77 = _EVAL_349[8:0];
  assign _EVAL_147 = _EVAL_3[0];
  assign _EVAL_311 = _EVAL_98 | _EVAL_12;
  assign _EVAL_279 = ~_EVAL_54;
  assign _EVAL_212 = _EVAL_1 & _EVAL_216;
  assign _EVAL_168 = 4'h2 == _EVAL_10;
  assign _EVAL_340 = ~_EVAL_257;
  assign _EVAL_102 = _EVAL[0];
  assign _EVAL_208 = _EVAL_32 | _EVAL_12;
  assign _EVAL_96 = ~_EVAL_311;
  assign _EVAL_46 = plusarg_reader_out == 32'h0;
  assign _EVAL_282 = _EVAL_144 | _EVAL_12;
  assign _EVAL_215 = _EVAL_13 & _EVAL_125;
  assign _EVAL_310 = _EVAL_206;
  assign _EVAL_238 = $signed(_EVAL_85) & -33'sh400000;
  assign _EVAL_22 = _EVAL_130 == 6'h0;
  assign _EVAL_235 = _EVAL_164 | _EVAL_12;
  assign _EVAL_104 = _EVAL_18 <= 3'h4;
  assign _EVAL_178 = _EVAL_163 | _EVAL_12;
  assign _EVAL_79 = _EVAL_131 | 2'h1;
  assign _EVAL_231 = ~_EVAL_242;
  assign _EVAL_360 = _EVAL_179 == 4'h0;
  assign _EVAL_284 = _EVAL_11 != 2'h2;
  assign _EVAL_226 = 16'h1 << _EVAL_7;
  assign _EVAL_266 = _EVAL_342 & _EVAL_250;
  assign _EVAL_323 = _EVAL_320 | _EVAL_0;
  assign _EVAL_141 = _EVAL_49 | _EVAL_372;
  assign _EVAL_53 = _EVAL_6 & _EVAL_129;
  assign _EVAL_304 = _EVAL_10 == _EVAL_103;
  assign _EVAL_137 = _EVAL_182 | _EVAL_299;
  assign _EVAL_89 = _EVAL_186 & _EVAL_221;
  assign _EVAL_118 = $signed(_EVAL_33) & -33'sh4000;
  assign _EVAL_368 = _EVAL_7 == _EVAL_123;
  assign _EVAL_267 = _EVAL_16 == 3'h3;
  assign _EVAL_135 = _EVAL_110 == 6'h0;
  assign _EVAL_263 = _EVAL_278 >> _EVAL_7;
  assign _EVAL_309 = _EVAL_71 | _EVAL_116;
  assign _EVAL_327 = _EVAL_297;
  assign _EVAL_370 = _EVAL_87 | _EVAL_12;
  assign _EVAL_314 = _EVAL_7[3];
  assign _EVAL_156 = _EVAL_227 | _EVAL_36;
  assign _EVAL_329 = _EVAL_13 & _EVAL_64;
  assign _EVAL_225 = ~_EVAL_183;
  assign _EVAL_34 = _EVAL_18 <= 3'h2;
  assign _EVAL_58 = _EVAL_13 & _EVAL_356;
  assign _EVAL_38 = {1'b0,$signed(_EVAL_343)};
  assign _EVAL_244 = _EVAL_29 == 32'h0;
  assign _EVAL_82 = _EVAL_70 | _EVAL_139;
  assign _EVAL_88 = _EVAL_94[7:0];
  assign _EVAL_334 = ~_EVAL_160;
  assign _EVAL_190 = ~_EVAL_314;
  assign _EVAL_191 = ~_EVAL_167;
  assign _EVAL_230 = _EVAL_1 & _EVAL_19;
  assign _EVAL_192 = _EVAL_16[2];
  assign _EVAL_144 = _EVAL_70 | _EVAL_219;
  assign _EVAL_253 = _EVAL_220 | _EVAL_247;
  assign _EVAL_237 = _EVAL_347 | _EVAL_12;
  assign _EVAL_76 = ~_EVAL_52;
  assign _EVAL_47 = _EVAL_13 & _EVAL_267;
  assign _EVAL_91 = _EVAL_18 <= 3'h1;
  assign _EVAL_171 = ~_EVAL_235;
  assign _EVAL_161 = _EVAL ^ 32'h3000;
  assign _EVAL_259 = _EVAL_78 | _EVAL_12;
  assign _EVAL_185 = ~_EVAL_23;
  assign _EVAL_229 = _EVAL_173 & _EVAL_90;
  assign _EVAL_294 = ~_EVAL_102;
  assign _EVAL_242 = |_EVAL_217;
  assign _EVAL_75 = ~_EVAL_303;
  assign _EVAL_196 = ~_EVAL_43;
  assign _EVAL_216 = ~_EVAL_135;
  assign _EVAL_83 = _EVAL_145 | _EVAL_12;
  assign _EVAL_303 = _EVAL_15[3];
  assign _EVAL_280 = ~_EVAL_62;
  assign _EVAL_158 = ~_EVAL_313;
  assign _EVAL_121 = _EVAL_1 & _EVAL_140;
  assign _EVAL_98 = _EVAL_18 == _EVAL_176;
  assign _EVAL_307 = _EVAL_268 & _EVAL_102;
  assign _EVAL_163 = _EVAL_165 | _EVAL_301;
  assign _EVAL_318 = _EVAL_5 & _EVAL_1;
  assign _EVAL_19 = _EVAL_3 == 3'h0;
  assign _EVAL_299 = _EVAL_346 < plusarg_reader_out;
  assign _EVAL_74 = _EVAL_367 | _EVAL_202;
  assign _EVAL_363 = _EVAL_291[5:0];
  assign _EVAL_291 = _EVAL_130 - 6'h1;
  assign _EVAL_112 = _EVAL_18 != 3'h0;
  assign _EVAL_300 = $signed(_EVAL_119) == 33'sh0;
  assign _EVAL_349 = _EVAL_289 ? _EVAL_226 : 16'h0;
  assign _EVAL_172 = _EVAL_229 | _EVAL_12;
  assign _EVAL_107 = _EVAL_238;
  assign _EVAL_68 = ~_EVAL_50;
  assign _EVAL_111 = _EVAL_112 | _EVAL_12;
  assign _EVAL_287 = _EVAL_16 == 3'h1;
  assign _EVAL_199 = _EVAL_244 | _EVAL_12;
  assign _EVAL_223 = _EVAL_37 <= 3'h6;
  assign _EVAL_108 = _EVAL_177 | _EVAL_12;
  assign _EVAL_193 = _EVAL_366 | _EVAL_12;
  assign _EVAL_148 = _EVAL_56 | _EVAL_12;
  assign _EVAL_371 = _EVAL_141 | _EVAL_120;
  assign _EVAL_164 = _EVAL_3 == _EVAL_324;
  assign _EVAL_331 = {1'b0,$signed(_EVAL_188)};
  assign _EVAL_249 = ~_EVAL_236;
  assign _EVAL_87 = ~_EVAL_0;
  assign _EVAL_356 = _EVAL_16 == 3'h4;
  assign _EVAL_330 = _EVAL_11 <= 2'h2;
  assign _EVAL_33 = {1'b0,$signed(_EVAL_72)};
  assign _EVAL_245 = _EVAL ^ 32'h2000000;
  assign _EVAL_115 = _EVAL_187 | _EVAL_318;
  assign _EVAL_258 = _EVAL_318 & _EVAL_135;
  assign _EVAL_165 = _EVAL_190 & _EVAL_26;
  assign _EVAL_69 = _EVAL_10 >= 4'h2;
  assign _EVAL_281 = _EVAL_322 | _EVAL_12;
  assign _EVAL_166 = ~_EVAL_370;
  assign _EVAL_116 = _EVAL_15 == 4'h8;
  assign _EVAL_213 = ~_EVAL_41;
  assign _EVAL_326 = ~_EVAL_83;
  assign _EVAL_127 = _EVAL_1 & _EVAL_336;
  assign _EVAL_109 = ~_EVAL_172;
  assign _EVAL_218 = ~_EVAL_51;
  assign _EVAL_257 = _EVAL_162 | _EVAL_12;
  assign _EVAL_301 = _EVAL_7 == 4'h8;
  assign _EVAL_305 = ~_EVAL_207;
  assign _EVAL_42 = _EVAL_11 == _EVAL_243;
  assign _EVAL_342 = _EVAL_79[0];
  assign _EVAL_202 = $signed(_EVAL_180) == 33'sh0;
  assign _EVAL_61 = ~_EVAL_358;
  assign _EVAL_322 = _EVAL_18 <= 3'h3;
  assign _EVAL_271 = _EVAL_81[7:2];
  assign _EVAL_162 = _EVAL_16 == _EVAL_211;
  assign _EVAL_286 = _EVAL_260[8:0];
  assign _EVAL_197 = _EVAL_186 & _EVAL_268;
  assign _EVAL_224 = _EVAL_13 & _EVAL_195;
  assign _EVAL_358 = _EVAL_320 | _EVAL_12;
  assign _EVAL_50 = _EVAL_328 | _EVAL_12;
  assign _EVAL_337 = ~_EVAL_88;
  assign _EVAL_222 = ~_EVAL_39;
  assign _EVAL_319 = _EVAL_14 >= 4'h2;
  assign _EVAL_131 = 2'h1 << _EVAL_157;
  assign _EVAL_99 = _EVAL_290 | _EVAL_12;
  assign _EVAL_44 = ~_EVAL_198;
  assign _EVAL_339 = _EVAL_25;
  assign _EVAL_201 = _EVAL_3 == 3'h1;
  assign _EVAL_134 = _EVAL_203[31:0];
  assign _EVAL_106 = _EVAL_3 <= 3'h6;
  assign _EVAL_355 = _EVAL_367 | _EVAL_120;
  assign _EVAL_200 = $signed(_EVAL_339) == 33'sh0;
  assign _EVAL_122 = _EVAL_293[7:0];
  assign _EVAL_55 = ~_EVAL_199;
  assign _EVAL_234 = ~_EVAL_86;
  assign _EVAL_81 = ~_EVAL_122;
  assign _EVAL_228 = _EVAL_1 & _EVAL_335;
  assign _EVAL_295 = _EVAL_82 | _EVAL_12;
  assign _EVAL_151 = ~_EVAL_99;
  assign _EVAL_113 = _EVAL_265 == 6'h0;
  assign _EVAL_270 = _EVAL_10 <= 4'h8;
  assign _EVAL_313 = _EVAL_69 | _EVAL_12;
  assign _EVAL_100 = _EVAL_138;
  assign _EVAL_272 = _EVAL_16 == 3'h5;
  assign _EVAL_92 = _EVAL_69 | _EVAL_89;
  assign _EVAL_30 = {{24'd0}, _EVAL_337};
  assign _EVAL_247 = $signed(_EVAL_310) == 33'sh0;
  assign _EVAL_335 = _EVAL_3 == 3'h4;
  assign _EVAL_150 = _EVAL_312[5:0];
  assign _EVAL_169 = _EVAL_45 & _EVAL_255;
  assign _EVAL_188 = _EVAL ^ 32'h1800000;
  assign _EVAL_209 = ~_EVAL_232;
  assign _EVAL_362 = ~_EVAL_17;
  assign _EVAL_26 = _EVAL_321 <= 3'h6;
  assign _EVAL_24 = _EVAL_16 == 3'h6;
  assign _EVAL_145 = _EVAL_15 == _EVAL_283;
  assign _EVAL_155 = _EVAL_104 | _EVAL_12;
  assign _EVAL_182 = _EVAL_231 | _EVAL_46;
  assign _EVAL_154 = _EVAL_268 & _EVAL_294;
  assign _EVAL_367 = _EVAL_308 | _EVAL_372;
  assign _EVAL_23 = _EVAL_254 | _EVAL_12;
  assign _EVAL_278 = _EVAL_286 | _EVAL_217;
  assign _EVAL_174 = ~_EVAL_365;
  assign _EVAL_353 = _EVAL_351 & _EVAL_66;
  assign _EVAL_32 = _EVAL_273 | _EVAL_218;
  assign _EVAL_347 = _EVAL_263[0];
  assign _EVAL_241 = _EVAL_42 | _EVAL_12;
  assign _EVAL_142 = _EVAL_187 & _EVAL_22;
  assign _EVAL_52 = _EVAL_368 | _EVAL_12;
  assign _EVAL_264 = _EVAL ^ 32'hc000000;
  assign _EVAL_251 = ~_EVAL_259;
  assign _EVAL_344 = _EVAL_124;
  assign _EVAL_157 = _EVAL_10[0];
  assign _EVAL_128 = ~_EVAL_97;
  assign _EVAL_129 = ~_EVAL_332;
  assign _EVAL_239 = $signed(_EVAL_331) & -33'sh4000;
  assign _EVAL_269 = _EVAL_187 & _EVAL_31;
  assign _EVAL_204 = ~_EVAL_93;
  assign _EVAL_359 = _EVAL_120 | _EVAL_146;
  assign _EVAL_86 = _EVAL_341 | _EVAL_12;
  assign _EVAL_85 = {1'b0,$signed(_EVAL_264)};
  assign _EVAL_170 = ~_EVAL_237;
  assign _EVAL_54 = _EVAL_330 | _EVAL_12;
  assign _EVAL_183 = _EVAL_252 | _EVAL_12;
  assign _EVAL_214 = _EVAL_16 == 3'h0;
  assign _EVAL_306 = _EVAL_91 | _EVAL_12;
  assign _EVAL_252 = _EVAL_14 == _EVAL_298;
  assign _EVAL_184 = _EVAL_13 & _EVAL_272;
  assign _EVAL_203 = _EVAL_346 + 32'h1;
  assign _EVAL_198 = _EVAL_95 | _EVAL_12;
  assign _EVAL_73 = _EVAL_318 & _EVAL_113;
  assign _EVAL_153 = {1'b0,$signed(_EVAL_285)};
  assign _EVAL_94 = 23'hff << _EVAL_10;
  assign _EVAL_27 = _EVAL_84[5:0];
  assign _EVAL_293 = 23'hff << _EVAL_14;
  assign _EVAL_37 = _EVAL_15[2:0];
  assign _EVAL_194 = ~_EVAL_192;
  assign _EVAL_49 = _EVAL_159 | _EVAL_200;
  assign _EVAL_101 = ~_EVAL_208;
  assign _EVAL_132 = 4'h6 == _EVAL_10;
  assign _EVAL_40 = ~_EVAL_281;
  assign _EVAL_124 = $signed(_EVAL_153) & -33'sh2000;
  assign _EVAL_343 = _EVAL ^ 32'h40000000;
  assign _EVAL_70 = _EVAL_270 & _EVAL_247;
  assign _EVAL_268 = ~_EVAL_221;
  assign _EVAL_338 = _EVAL_355 | _EVAL_146;
  assign _EVAL_180 = _EVAL_118;
  assign _EVAL_146 = $signed(_EVAL_327) == 33'sh0;
  assign _EVAL_60 = _EVAL_132 & _EVAL_116;
  assign _EVAL_39 = _EVAL_106 | _EVAL_12;
  assign _EVAL_186 = _EVAL_79[1];
  assign _EVAL_250 = _EVAL_221 & _EVAL_294;
  assign _EVAL_341 = _EVAL_11 == 2'h0;
  assign _EVAL_125 = _EVAL_16 == 3'h7;
  assign _EVAL_289 = _EVAL_73 & _EVAL_174;
  assign _EVAL_43 = _EVAL_323 | _EVAL_12;
  assign _EVAL_321 = _EVAL_7[2:0];
  assign _EVAL_336 = _EVAL_3 == 3'h5;
  assign _EVAL_273 = _EVAL_286 != _EVAL_77;
  assign _EVAL_105 = ~_EVAL_178;
  assign _EVAL_352 = _EVAL_92 | _EVAL_266;
  assign _EVAL_207 = _EVAL_319 | _EVAL_12;
  assign _EVAL_246 = ~_EVAL_295;
  assign _EVAL_140 = _EVAL_3 == 3'h2;
  assign _EVAL_312 = _EVAL_265 - 6'h1;
  assign _EVAL_262 = _EVAL_13 & _EVAL_287;
  assign _EVAL_189 = ~_EVAL_148;
  assign _EVAL_63 = ~_EVAL_108;
  assign _EVAL_345 = _EVAL_342 & _EVAL_277;
  assign _EVAL_290 = _EVAL == _EVAL_315;
  assign _EVAL_350 = _EVAL_13 & _EVAL_214;
  assign _EVAL_365 = _EVAL_3 == 3'h6;
  assign _EVAL_21 = ~_EVAL_241;
  assign _EVAL_72 = _EVAL ^ 32'h80000000;
  assign _EVAL_332 = {_EVAL_364,_EVAL_352,_EVAL_156,_EVAL_80};
  assign _EVAL_64 = _EVAL_16 == 3'h2;
  assign _EVAL_160 = _EVAL_249 | _EVAL_12;
  assign _EVAL_84 = _EVAL_110 - 6'h1;
  assign _EVAL_51 = |_EVAL_286;
  assign _EVAL_254 = _EVAL_53 == 4'h0;
  assign _EVAL_361 = _EVAL_13 & _EVAL_24;
  assign _EVAL_227 = _EVAL_69 | _EVAL_197;
  assign _EVAL_36 = _EVAL_342 & _EVAL_307;
  assign _EVAL_372 = $signed(_EVAL_107) == 33'sh0;
  assign _EVAL_45 = _EVAL_10 <= 4'h6;
  assign _EVAL_57 = {1'b0,$signed(_EVAL)};
  assign _EVAL_28 = ~_EVAL_306;
  assign _EVAL_159 = _EVAL_253 | _EVAL_300;
  assign _EVAL_181 = ~_EVAL_12;
  assign _EVAL_232 = _EVAL_360 | _EVAL_12;
  assign _EVAL_120 = $signed(_EVAL_344) == 33'sh0;
  assign _EVAL_308 = _EVAL_117 | _EVAL_200;
  assign _EVAL_62 = _EVAL_309 | _EVAL_12;
  assign _EVAL_167 = _EVAL_362 | _EVAL_12;
  assign _EVAL_119 = _EVAL_239;
  assign _EVAL_261 = ~_EVAL_155;
  assign _EVAL_369 = _EVAL_10 <= 4'h2;
  assign _EVAL_177 = _EVAL_18 == 3'h0;
  assign _EVAL_90 = _EVAL_369 & _EVAL_288;
  assign _EVAL_260 = _EVAL_142 ? _EVAL_126 : 16'h0;
  assign _EVAL_56 = _EVAL_6 == _EVAL_332;
  assign _EVAL_277 = _EVAL_221 & _EVAL_102;
  assign _EVAL_364 = _EVAL_92 | _EVAL_345;
  assign _EVAL_67 = _EVAL_316[5:0];
  assign _EVAL_328 = _EVAL_70 | _EVAL_169;
  assign _EVAL_276 = _EVAL_205 | _EVAL_60;
  assign _EVAL_221 = _EVAL[1];
  assign _EVAL_297 = $signed(_EVAL_38) & -33'sh2000;
  assign _EVAL_95 = _EVAL_8 == _EVAL_296;
  assign _EVAL_143 = ~_EVAL_59;
  assign _EVAL_136 = ~_EVAL_282;
  assign _EVAL_93 = _EVAL_34 | _EVAL_12;
  assign _EVAL_351 = _EVAL_217 | _EVAL_286;
  assign _EVAL_149 = _EVAL_337[7:2];
  assign _EVAL_333 = _EVAL_1 & _EVAL_201;
  assign _EVAL_285 = _EVAL ^ 32'h20000000;
  assign _EVAL_117 = _EVAL_220 | _EVAL_300;
  assign _EVAL_80 = _EVAL_227 | _EVAL_275;
  assign _EVAL_41 = _EVAL_137 | _EVAL_12;
  assign _EVAL_59 = _EVAL_304 | _EVAL_12;
  assign _EVAL_78 = _EVAL_4 == _EVAL_256;
  assign _EVAL_25 = $signed(_EVAL_302) & -33'sh10000;
  assign _EVAL_248 = _EVAL_284 | _EVAL_12;
  assign _EVAL_302 = {1'b0,$signed(_EVAL_245)};
  assign _EVAL_366 = _EVAL_205 & _EVAL_328;
  assign _EVAL_275 = _EVAL_342 & _EVAL_154;
  assign _EVAL_179 = ~_EVAL_6;
  assign _EVAL_320 = ~_EVAL_4;
  assign _EVAL_205 = _EVAL_369 & _EVAL_71;
  assign _EVAL_236 = _EVAL_354[0];
  assign _EVAL_66 = ~_EVAL_77;
  assign _EVAL_126 = 16'h1 << _EVAL_15;
  assign _EVAL_29 = _EVAL & _EVAL_30;
  assign _EVAL_31 = _EVAL_240 == 6'h0;
  assign _EVAL_71 = _EVAL_75 & _EVAL_223;
  assign _EVAL_354 = _EVAL_217 >> _EVAL_15;
  assign _EVAL_255 = _EVAL_338 | _EVAL_202;
  assign _EVAL_97 = _EVAL_276 | _EVAL_12;
  assign _EVAL_292 = ~_EVAL_111;
  assign _EVAL_220 = $signed(_EVAL_100) == 33'sh0;
  assign _EVAL_175 = ~_EVAL_193;
  always @(posedge _EVAL_9) begin
    if (_EVAL_269) begin
      _EVAL_103 <= _EVAL_10;
    end
    if (_EVAL_12) begin
      _EVAL_110 <= 6'h0;
    end else if (_EVAL_318) begin
      if (_EVAL_135) begin
        if (_EVAL_147) begin
          _EVAL_110 <= _EVAL_271;
        end else begin
          _EVAL_110 <= 6'h0;
        end
      end else begin
        _EVAL_110 <= _EVAL_27;
      end
    end
    if (_EVAL_258) begin
      _EVAL_123 <= _EVAL_7;
    end
    if (_EVAL_12) begin
      _EVAL_130 <= 6'h0;
    end else if (_EVAL_187) begin
      if (_EVAL_22) begin
        if (_EVAL_194) begin
          _EVAL_130 <= _EVAL_149;
        end else begin
          _EVAL_130 <= 6'h0;
        end
      end else begin
        _EVAL_130 <= _EVAL_363;
      end
    end
    if (_EVAL_269) begin
      _EVAL_176 <= _EVAL_18;
    end
    if (_EVAL_269) begin
      _EVAL_211 <= _EVAL_16;
    end
    if (_EVAL_12) begin
      _EVAL_217 <= 9'h0;
    end else begin
      _EVAL_217 <= _EVAL_353;
    end
    if (_EVAL_12) begin
      _EVAL_240 <= 6'h0;
    end else if (_EVAL_187) begin
      if (_EVAL_31) begin
        if (_EVAL_194) begin
          _EVAL_240 <= _EVAL_149;
        end else begin
          _EVAL_240 <= 6'h0;
        end
      end else begin
        _EVAL_240 <= _EVAL_67;
      end
    end
    if (_EVAL_258) begin
      _EVAL_243 <= _EVAL_11;
    end
    if (_EVAL_258) begin
      _EVAL_256 <= _EVAL_4;
    end
    if (_EVAL_12) begin
      _EVAL_265 <= 6'h0;
    end else if (_EVAL_318) begin
      if (_EVAL_113) begin
        if (_EVAL_147) begin
          _EVAL_265 <= _EVAL_271;
        end else begin
          _EVAL_265 <= 6'h0;
        end
      end else begin
        _EVAL_265 <= _EVAL_150;
      end
    end
    if (_EVAL_269) begin
      _EVAL_283 <= _EVAL_15;
    end
    if (_EVAL_258) begin
      _EVAL_296 <= _EVAL_8;
    end
    if (_EVAL_258) begin
      _EVAL_298 <= _EVAL_14;
    end
    if (_EVAL_269) begin
      _EVAL_315 <= _EVAL;
    end
    if (_EVAL_258) begin
      _EVAL_324 <= _EVAL_3;
    end
    if (_EVAL_12) begin
      _EVAL_346 <= 32'h0;
    end else if (_EVAL_115) begin
      _EVAL_346 <= 32'h0;
    end else begin
      _EVAL_346 <= _EVAL_134;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd32edb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_334) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc5df332)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_305) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_96) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_329 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50dbcb66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf18667)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_329 & _EVAL_261) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e911f3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_350 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba0c689a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7aa4e25a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bd69cdd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a520eb5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78dccd4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cc4c8ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf40a209)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(673025e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_350 & _EVAL_175) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b425311f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_151) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_128) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4cd65140)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_305) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4965884b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5098eeb9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2944ab2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_329 & _EVAL_261) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_329 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c823235)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f27aa2a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b6ed1a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2604591a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74d7a379)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(866d1427)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc92f8fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4c43ff4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3fe0f66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_305) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_350 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b33fb96d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8960701a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_340) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1716f46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e09c0a1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_326) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26005506)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_333 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3c3832c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(428a8031)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_305) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69c3f14e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_350 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(372680bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5afe4a02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_329 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_329 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c83bc2bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cdc8723)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4355f22a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_151) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0c5e0ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_333 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_350 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d82cfb5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_334) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_233) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_171) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_333 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_21) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8567bdd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c693ccd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_350 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(239265bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9dab4af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b89ee5e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_21) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_28) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_329 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_329 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c83d618)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba9d95a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1760bfe4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d68e1cff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_350 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(487ed2a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_189) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16e2c774)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bac9332)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(673025e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(270ee79b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(704a3c6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12e82b18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_292) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(668c1373)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_329 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_28) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(925a94f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a74b8f6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_63) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b61e7c11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca9c913c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db284749)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20b10ecf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_128) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_333 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af98b544)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_222) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_105) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd1d627b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1 & _EVAL_222) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc9e5fc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(380484fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_233) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ea753dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_305) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a228683e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41f888d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d488a9b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_171) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4b8a785)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1515931c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_305) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb74aef3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8450a04a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_350 & _EVAL_175) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77084b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_333 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86fe575a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a59fcd76)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_333 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5b3da55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b7b7742)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_340) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bf91190)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_215 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(196cbe9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d9a5927)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_350 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ebcfdb69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_96) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b52ab7e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f68e7df8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_361 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5d7f0dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_105) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_127 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db72bd6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_329 & _EVAL_189) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f31f87f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_58 & _EVAL_63) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2f46065)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_224 & _EVAL_326) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_350 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_152 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c52c166)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(126d057a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_103 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_110 = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_123 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_130 = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_176 = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_211 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_217 = _RAND_6[8:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_240 = _RAND_7[5:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_243 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_256 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_265 = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_283 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_296 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_298 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_315 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_324 = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_346 = _RAND_16[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
