//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_102_assert(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [1:0]  _EVAL_2,
  input         _EVAL_3,
  input  [2:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input  [31:0] _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input  [3:0]  _EVAL_11
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] _EVAL_12;
  wire  _EVAL_13;
  wire  _EVAL_14;
  wire [32:0] _EVAL_15;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire [6:0] _EVAL_19;
  wire [32:0] _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire [22:0] _EVAL_27;
  wire  _EVAL_28;
  wire [31:0] _EVAL_29;
  wire  _EVAL_30;
  wire [32:0] _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire [32:0] _EVAL_34;
  wire [32:0] _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  reg [2:0] _EVAL_39;
  wire  _EVAL_40;
  wire [31:0] _EVAL_41;
  wire  _EVAL_42;
  reg [31:0] _EVAL_43;
  wire [7:0] _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire [5:0] _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire [32:0] _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire [31:0] _EVAL_54;
  wire  _EVAL_56;
  wire  _EVAL_58;
  wire [31:0] _EVAL_59;
  wire [7:0] _EVAL_60;
  wire [5:0] _EVAL_61;
  wire [31:0] _EVAL_62;
  wire  _EVAL_63;
  wire [32:0] _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire [32:0] _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_75;
  wire [32:0] _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire [6:0] _EVAL_84;
  wire [32:0] _EVAL_85;
  reg [5:0] _EVAL_86;
  wire  _EVAL_87;
  wire [32:0] _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire [32:0] _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  reg [5:0] _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire [32:0] _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  reg [3:0] _EVAL_114;
  wire  _EVAL_115;
  wire [32:0] _EVAL_116;
  wire  _EVAL_117;
  reg  _EVAL_118;
  wire  _EVAL_119;
  wire [32:0] _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire [32:0] _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire [32:0] _EVAL_128;
  wire  _EVAL_129;
  reg [5:0] _EVAL_130;
  wire [32:0] _EVAL_131;
  wire  _EVAL_132;
  wire [32:0] _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_139;
  wire [32:0] _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire [32:0] _EVAL_147;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire [6:0] _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire [32:0] _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire [5:0] _EVAL_165;
  wire  _EVAL_166;
  wire [5:0] _EVAL_167;
  wire [32:0] _EVAL_169;
  wire  _EVAL_170;
  wire [31:0] plusarg_reader_out;
  reg  _EVAL_171;
  wire  _EVAL_172;
  wire [31:0] _EVAL_173;
  reg [1:0] _EVAL_174;
  wire  _EVAL_175;
  wire [32:0] _EVAL_176;
  wire [31:0] _EVAL_177;
  reg [5:0] _EVAL_178;
  wire  _EVAL_179;
  wire [31:0] _EVAL_180;
  wire  _EVAL_181;
  wire [6:0] _EVAL_182;
  wire  _EVAL_183;
  wire [32:0] _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire [31:0] _EVAL_189;
  wire [1:0] _EVAL_190;
  wire [5:0] _EVAL_191;
  wire  _EVAL_193;
  reg  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire [1:0] _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_83 = _EVAL_90 | _EVAL_6;
  assign _EVAL_188 = _EVAL_91 & _EVAL_66;
  assign _EVAL_14 = _EVAL_23 | _EVAL_94;
  assign _EVAL_123 = _EVAL_86 == 6'h0;
  assign _EVAL_63 = _EVAL_22 | _EVAL_6;
  assign _EVAL_173 = _EVAL_128[31:0];
  assign _EVAL_93 = _EVAL_169;
  assign _EVAL_33 = ~_EVAL_13;
  assign _EVAL_102 = _EVAL_0 & _EVAL_24;
  assign _EVAL_197 = _EVAL_159 ? 2'h1 : 2'h0;
  assign _EVAL_51 = $signed(_EVAL_76) & -33'sh1000;
  assign _EVAL_142 = _EVAL_11 >= 4'h2;
  assign _EVAL_34 = _EVAL_184;
  assign _EVAL_84 = _EVAL_178 - 6'h1;
  assign _EVAL_41 = _EVAL_8 ^ 32'h1800000;
  assign _EVAL_76 = {1'b0,$signed(_EVAL_180)};
  assign _EVAL_129 = $signed(_EVAL_15) == 33'sh0;
  assign _EVAL_71 = {1'b0,$signed(_EVAL_29)};
  assign _EVAL_131 = _EVAL_121;
  assign _EVAL_156 = _EVAL_196 | _EVAL_154;
  assign _EVAL_80 = ~_EVAL_149;
  assign _EVAL_161 = _EVAL_110 | _EVAL_6;
  assign _EVAL_104 = _EVAL_46 | _EVAL_179;
  assign _EVAL_144 = _EVAL_163 & _EVAL_150;
  assign _EVAL_163 = _EVAL_9 & _EVAL;
  assign _EVAL_78 = _EVAL_8 == _EVAL_12;
  assign _EVAL_146 = _EVAL_4 == 3'h1;
  assign _EVAL_19 = _EVAL_96 - 6'h1;
  assign _EVAL_44 = _EVAL_27[7:0];
  assign _EVAL_189 = _EVAL_8 ^ 32'hc000000;
  assign _EVAL_121 = $signed(_EVAL_88) & -33'sh5000;
  assign _EVAL_37 = ~_EVAL_47;
  assign _EVAL_151 = _EVAL_130 - 6'h1;
  assign _EVAL_85 = $signed(_EVAL_176) & -33'sh400000;
  assign _EVAL_65 = ~_EVAL_68;
  assign _EVAL_139 = _EVAL_4 <= 3'h6;
  assign _EVAL_195 = ~_EVAL_150;
  assign _EVAL_116 = {1'b0,$signed(_EVAL_62)};
  assign _EVAL_97 = _EVAL_45 | _EVAL_3;
  assign _EVAL_82 = _EVAL_0 & _EVAL_100;
  assign _EVAL_159 = _EVAL_163 & _EVAL_53;
  assign _EVAL_162 = ~_EVAL_72;
  assign _EVAL_196 = ~_EVAL_112;
  assign _EVAL_108 = ~_EVAL_25;
  assign _EVAL_183 = _EVAL_4 == 3'h4;
  assign _EVAL_110 = _EVAL_4 == _EVAL_39;
  assign _EVAL_53 = _EVAL_96 == 6'h0;
  assign _EVAL_64 = $signed(_EVAL_71) & -33'sh2000;
  assign _EVAL_155 = _EVAL_2 <= 2'h2;
  assign _EVAL_191 = _EVAL_151[5:0];
  assign _EVAL_15 = _EVAL_147;
  assign _EVAL_42 = ~_EVAL_6;
  assign _EVAL_35 = {1'b0,$signed(_EVAL_54)};
  assign _EVAL_49 = _EVAL_50 & _EVAL_124;
  assign _EVAL_141 = _EVAL_11 == _EVAL_114;
  assign _EVAL_198 = _EVAL_0 & _EVAL_137;
  assign _EVAL_54 = _EVAL_8 ^ 32'h20000000;
  assign _EVAL_169 = $signed(_EVAL_125) & -33'sh10000;
  assign _EVAL_153 = $signed(_EVAL_140) == 33'sh0;
  assign _EVAL_176 = {1'b0,$signed(_EVAL_189)};
  assign _EVAL_164 = _EVAL_1 & _EVAL_0;
  assign _EVAL_73 = _EVAL_177 == 32'h0;
  assign _EVAL_56 = ~_EVAL_193;
  assign _EVAL_45 = ~_EVAL_10;
  assign _EVAL_17 = _EVAL_190[0];
  assign _EVAL_165 = _EVAL_19[5:0];
  assign _EVAL_133 = $signed(_EVAL_31) & -33'sh4000;
  assign _EVAL_50 = _EVAL_164 & _EVAL_170;
  assign _EVAL_147 = $signed(_EVAL_116) & -33'sh4000;
  assign _EVAL_60 = ~_EVAL_44;
  assign _EVAL_132 = _EVAL_77 | _EVAL_6;
  assign _EVAL_88 = {1'b0,$signed(_EVAL_8)};
  assign _EVAL_87 = ~_EVAL_21;
  assign _EVAL_22 = _EVAL_187 | _EVAL_194;
  assign _EVAL_149 = _EVAL_78 | _EVAL_6;
  assign _EVAL_23 = _EVAL_52 | _EVAL_153;
  assign _EVAL_150 = _EVAL_130 == 6'h0;
  assign _EVAL_193 = _EVAL_199 | _EVAL_6;
  assign _EVAL_100 = _EVAL_4 == 3'h0;
  assign _EVAL_47 = _EVAL_181 | _EVAL_6;
  assign _EVAL_58 = _EVAL_119 | _EVAL_6;
  assign _EVAL_124 = ~_EVAL_98;
  assign _EVAL_13 = _EVAL_139 | _EVAL_6;
  assign _EVAL_24 = ~_EVAL_123;
  assign _EVAL_126 = _EVAL_164 & _EVAL_123;
  assign _EVAL_177 = _EVAL_8 & 32'h3f;
  assign _EVAL_32 = _EVAL_187 != _EVAL_17;
  assign _EVAL_98 = _EVAL_4 == 3'h6;
  assign _EVAL_59 = _EVAL_8 ^ 32'h2000000;
  assign _EVAL_128 = _EVAL_43 + 32'h1;
  assign _EVAL_109 = _EVAL_4 == 3'h2;
  assign _EVAL_20 = _EVAL_51;
  assign _EVAL_111 = ~_EVAL_38;
  assign _EVAL_122 = _EVAL_0 & _EVAL_98;
  assign _EVAL_119 = _EVAL_2 == _EVAL_174;
  assign _EVAL_175 = _EVAL_0 & _EVAL_109;
  assign _EVAL_66 = ~_EVAL_17;
  assign _EVAL_172 = _EVAL_0 & _EVAL_183;
  assign _EVAL_18 = _EVAL_2 == 2'h0;
  assign _EVAL_127 = _EVAL_101 | _EVAL_6;
  assign _EVAL_81 = _EVAL_97 | _EVAL_6;
  assign _EVAL_77 = ~_EVAL_3;
  assign _EVAL_103 = _EVAL_0 & _EVAL_146;
  assign _EVAL_31 = {1'b0,$signed(_EVAL_41)};
  assign _EVAL_62 = _EVAL_8 ^ 32'h80000000;
  assign _EVAL_184 = $signed(_EVAL_35) & -33'sh2000;
  assign _EVAL_46 = _EVAL_70 | _EVAL_69;
  assign _EVAL_158 = ~_EVAL_127;
  assign _EVAL_187 = _EVAL_197[0];
  assign _EVAL_89 = _EVAL_10 == _EVAL_118;
  assign _EVAL_16 = _EVAL_73 | _EVAL_6;
  assign _EVAL_186 = $signed(_EVAL_20) == 33'sh0;
  assign _EVAL_70 = _EVAL_14 | _EVAL_26;
  assign _EVAL_30 = _EVAL_5 == _EVAL_171;
  assign _EVAL_38 = _EVAL_135 | _EVAL_6;
  assign _EVAL_113 = ~_EVAL_58;
  assign _EVAL_105 = _EVAL_85;
  assign _EVAL_95 = ~_EVAL_92;
  assign _EVAL_61 = _EVAL_182[5:0];
  assign _EVAL_75 = ~_EVAL_81;
  assign _EVAL_152 = _EVAL_163 | _EVAL_164;
  assign _EVAL_117 = ~_EVAL_106;
  assign _EVAL_170 = _EVAL_178 == 6'h0;
  assign _EVAL_112 = |_EVAL_194;
  assign _EVAL_94 = $signed(_EVAL_93) == 33'sh0;
  assign _EVAL_134 = ~_EVAL_161;
  assign _EVAL_99 = _EVAL_104 | _EVAL_129;
  assign _EVAL_180 = _EVAL_8 ^ 32'h3000;
  assign _EVAL_140 = _EVAL_133;
  assign _EVAL_79 = _EVAL_89 | _EVAL_6;
  assign _EVAL_166 = ~_EVAL_28;
  assign _EVAL_106 = _EVAL_45 | _EVAL_6;
  assign _EVAL_26 = $signed(_EVAL_105) == 33'sh0;
  assign _EVAL_52 = $signed(_EVAL_131) == 33'sh0;
  assign _EVAL_154 = plusarg_reader_out == 32'h0;
  assign _EVAL_125 = {1'b0,$signed(_EVAL_59)};
  assign _EVAL_28 = _EVAL_30 | _EVAL_6;
  assign _EVAL_136 = ~_EVAL_16;
  assign _EVAL_181 = _EVAL_2 != 2'h2;
  assign _EVAL_92 = _EVAL_155 | _EVAL_6;
  assign _EVAL_199 = _EVAL_186 | _EVAL_99;
  assign _EVAL_68 = _EVAL_18 | _EVAL_6;
  assign _EVAL_115 = ~_EVAL_63;
  assign _EVAL_190 = _EVAL_49 ? 2'h1 : 2'h0;
  assign _EVAL_25 = _EVAL_142 | _EVAL_6;
  assign _EVAL_90 = _EVAL_156 | _EVAL_36;
  assign _EVAL_69 = $signed(_EVAL_34) == 33'sh0;
  assign _EVAL_91 = _EVAL_194 | _EVAL_187;
  assign _EVAL_137 = _EVAL_4 == 3'h5;
  assign _EVAL_179 = $signed(_EVAL_157) == 33'sh0;
  assign _EVAL_167 = _EVAL_84[5:0];
  assign _EVAL_72 = _EVAL_141 | _EVAL_6;
  assign _EVAL_157 = _EVAL_64;
  assign _EVAL_101 = ~_EVAL_194;
  assign _EVAL_40 = ~_EVAL_83;
  assign _EVAL_48 = _EVAL_60[7:2];
  assign _EVAL_27 = 23'hff << _EVAL_11;
  assign _EVAL_107 = _EVAL_4[0];
  assign _EVAL_29 = _EVAL_8 ^ 32'h40000000;
  assign _EVAL_36 = _EVAL_43 < plusarg_reader_out;
  assign _EVAL_21 = |_EVAL_187;
  assign _EVAL_145 = _EVAL & _EVAL_195;
  assign _EVAL_143 = ~_EVAL_132;
  assign _EVAL_185 = ~_EVAL_79;
  assign _EVAL_135 = _EVAL_32 | _EVAL_87;
  assign _EVAL_182 = _EVAL_86 - 6'h1;
  always @(posedge _EVAL_7) begin
    if (_EVAL_144) begin
      _EVAL_12 <= _EVAL_8;
    end
    if (_EVAL_126) begin
      _EVAL_39 <= _EVAL_4;
    end
    if (_EVAL_6) begin
      _EVAL_43 <= 32'h0;
    end else if (_EVAL_152) begin
      _EVAL_43 <= 32'h0;
    end else begin
      _EVAL_43 <= _EVAL_173;
    end
    if (_EVAL_6) begin
      _EVAL_86 <= 6'h0;
    end else if (_EVAL_164) begin
      if (_EVAL_123) begin
        if (_EVAL_107) begin
          _EVAL_86 <= _EVAL_48;
        end else begin
          _EVAL_86 <= 6'h0;
        end
      end else begin
        _EVAL_86 <= _EVAL_61;
      end
    end
    if (_EVAL_6) begin
      _EVAL_96 <= 6'h0;
    end else if (_EVAL_163) begin
      if (_EVAL_53) begin
        _EVAL_96 <= 6'h0;
      end else begin
        _EVAL_96 <= _EVAL_165;
      end
    end
    if (_EVAL_126) begin
      _EVAL_114 <= _EVAL_11;
    end
    if (_EVAL_126) begin
      _EVAL_118 <= _EVAL_10;
    end
    if (_EVAL_6) begin
      _EVAL_130 <= 6'h0;
    end else if (_EVAL_163) begin
      if (_EVAL_150) begin
        _EVAL_130 <= 6'h0;
      end else begin
        _EVAL_130 <= _EVAL_191;
      end
    end
    if (_EVAL_126) begin
      _EVAL_171 <= _EVAL_5;
    end
    if (_EVAL_126) begin
      _EVAL_174 <= _EVAL_2;
    end
    if (_EVAL_6) begin
      _EVAL_178 <= 6'h0;
    end else if (_EVAL_164) begin
      if (_EVAL_170) begin
        if (_EVAL_107) begin
          _EVAL_178 <= _EVAL_48;
        end else begin
          _EVAL_178 <= 6'h0;
        end
      end else begin
        _EVAL_178 <= _EVAL_167;
      end
    end
    if (_EVAL_6) begin
      _EVAL_194 <= 1'h0;
    end else begin
      _EVAL_194 <= _EVAL_188;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd4938f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6710e30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(832b957d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8a33a7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72966b06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_158) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85976b6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(566f3ff9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_0 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1f4cedf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4068dadb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea39d966)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_37) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_162) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98df4d4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fda4cb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_117) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e567447)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e74e6b14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf41452a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56c71061)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b711732)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6417bae5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_42) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3cf02463)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bdde700)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_158) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf8bcccc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_117) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7ac52c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5f7baec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_108) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4daa66ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69b0e161)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(baa0e81f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_143) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ae04dd3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3fded718)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0a8363d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_108) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68853594)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_37) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d44c5d12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_102 & _EVAL_162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_172 & _EVAL_42) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_103 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_82 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_143) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc60fc8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9166c134)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_122 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_12 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_39 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_43 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_86 = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_96 = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_114 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_118 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_130 = _RAND_7[5:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_171 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_174 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_178 = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_194 = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
