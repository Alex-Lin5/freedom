//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_13_assert(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  input  [30:0] _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input  [4:0]  _EVAL_4,
  input  [4:0]  _EVAL_5,
  input  [2:0]  _EVAL_6,
  input         _EVAL_7,
  input  [2:0]  _EVAL_8,
  input         _EVAL_9,
  input  [1:0]  _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input  [2:0]  _EVAL_14,
  input         _EVAL_15,
  input  [3:0]  _EVAL_16,
  input         _EVAL_17,
  input  [2:0]  _EVAL_18
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire [17:0] _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire [12:0] _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  reg [4:0] _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire [17:0] _EVAL_38;
  wire [3:0] _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  reg [2:0] _EVAL_48;
  reg [3:0] _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire [3:0] _EVAL_54;
  wire  _EVAL_55;
  wire [4:0] _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire [5:0] _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_69;
  wire  _EVAL_70;
  reg [4:0] _EVAL_71;
  wire  _EVAL_72;
  wire [31:0] _EVAL_73;
  reg [1:0] _EVAL_74;
  wire  _EVAL_75;
  wire [31:0] _EVAL_76;
  wire  _EVAL_77;
  wire [3:0] _EVAL_78;
  wire  _EVAL_79;
  reg [2:0] _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire [31:0] _EVAL_84;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  reg [2:0] _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire [3:0] _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire [17:0] _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  reg [3:0] _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire [5:0] _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire [4:0] _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire [17:0] _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire [3:0] _EVAL_130;
  wire  _EVAL_131;
  wire [5:0] _EVAL_132;
  wire [2:0] _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire [17:0] _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_146;
  wire  _EVAL_147;
  reg [31:0] _EVAL_148;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire [3:0] _EVAL_152;
  wire [5:0] _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_156;
  wire [12:0] _EVAL_157;
  wire [30:0] _EVAL_158;
  wire  _EVAL_159;
  wire [31:0] _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire [32:0] _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire [17:0] _EVAL_173;
  wire  _EVAL_174;
  wire [4:0] _EVAL_175;
  wire [2:0] _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire [31:0] _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  reg [3:0] _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  reg [3:0] _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire [3:0] _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire [30:0] _EVAL_220;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  reg [30:0] _EVAL_227;
  wire [31:0] _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire [1:0] _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire [1:0] _EVAL_236;
  wire [30:0] _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire [17:0] _EVAL_243;
  reg [17:0] _EVAL_244;
  wire  _EVAL_245;
  wire [3:0] _EVAL_246;
  reg [2:0] _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  reg  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire [31:0] _EVAL_265;
  wire  _EVAL_266;
  wire [31:0] _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  reg [2:0] _EVAL_272;
  wire  _EVAL_273;
  reg  _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire [1:0] _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire [17:0] _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire [4:0] _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_294;
  wire [3:0] _EVAL_295;
  wire  _EVAL_296;
  wire  _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_307;
  wire  _EVAL_308;
  wire  _EVAL_309;
  wire [3:0] _EVAL_310;
  wire  _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire [1:0] _EVAL_317;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_117 = ~_EVAL_62;
  assign _EVAL_23 = ~_EVAL_21;
  assign _EVAL_240 = _EVAL_13 == _EVAL_274;
  assign _EVAL_307 = _EVAL_9 & _EVAL_290;
  assign _EVAL_51 = _EVAL_150 & _EVAL_40;
  assign _EVAL_245 = _EVAL_317 == 2'h0;
  assign _EVAL_225 = ~_EVAL_110;
  assign _EVAL_224 = _EVAL_6 == 3'h1;
  assign _EVAL_165 = _EVAL_3 & _EVAL_151;
  assign _EVAL_111 = _EVAL_200 | _EVAL_101;
  assign _EVAL_138 = _EVAL_0 == _EVAL_272;
  assign _EVAL_276 = ~_EVAL_11;
  assign _EVAL_122 = _EVAL_27 | _EVAL_184;
  assign _EVAL_64 = _EVAL_10 == 2'h0;
  assign _EVAL_69 = _EVAL_28 | _EVAL_11;
  assign _EVAL_124 = _EVAL_243 & _EVAL_103;
  assign _EVAL_304 = _EVAL_9 & _EVAL_275;
  assign _EVAL_103 = ~_EVAL_38;
  assign _EVAL_192 = _EVAL_281 & _EVAL_241;
  assign _EVAL_232 = _EVAL_6 == 3'h0;
  assign _EVAL_231 = _EVAL_229 | _EVAL_11;
  assign _EVAL_228 = _EVAL_63 ? _EVAL_187 : 32'h0;
  assign _EVAL_44 = _EVAL_77 & _EVAL_219;
  assign _EVAL_87 = _EVAL_90 | _EVAL_96;
  assign _EVAL_115 = _EVAL_0 <= 3'h2;
  assign _EVAL_55 = _EVAL_18 == 3'h0;
  assign _EVAL_213 = _EVAL_147 & _EVAL_293;
  assign _EVAL_116 = _EVAL_55 | _EVAL_11;
  assign _EVAL_161 = _EVAL_3 & _EVAL_218;
  assign _EVAL_56 = _EVAL_107 - 4'h1;
  assign _EVAL_295 = _EVAL_16 & _EVAL_130;
  assign _EVAL_282 = _EVAL_193 | _EVAL_11;
  assign _EVAL_252 = _EVAL_300 | _EVAL_11;
  assign _EVAL_46 = _EVAL_259 | _EVAL_11;
  assign _EVAL_177 = ~_EVAL_262;
  assign _EVAL_255 = _EVAL_226 | _EVAL_11;
  assign _EVAL_136 = ~_EVAL_289;
  assign _EVAL_226 = _EVAL_34 & _EVAL_143;
  assign _EVAL_246 = _EVAL_56[3:0];
  assign _EVAL_125 = _EVAL_183 & _EVAL_119;
  assign _EVAL_222 = _EVAL_3 & _EVAL_266;
  assign _EVAL_263 = _EVAL_300 | _EVAL_51;
  assign _EVAL_204 = _EVAL_281 & _EVAL_202;
  assign _EVAL_273 = ~_EVAL_17;
  assign _EVAL_100 = |_EVAL_244;
  assign _EVAL_158 = _EVAL_1 & _EVAL_237;
  assign _EVAL_218 = _EVAL_14 == 3'h0;
  assign _EVAL_34 = _EVAL_0 <= 3'h6;
  assign _EVAL_75 = _EVAL_14[0];
  assign _EVAL_313 = ~_EVAL_69;
  assign _EVAL_206 = _EVAL_5 == 5'h10;
  assign _EVAL_258 = ~_EVAL_46;
  assign _EVAL_254 = _EVAL_250 | _EVAL_314;
  assign _EVAL_310 = _EVAL_132[5:2];
  assign _EVAL_188 = _EVAL_270 | _EVAL_11;
  assign _EVAL_76 = _EVAL_166[31:0];
  assign _EVAL_108 = _EVAL_107 == 4'h0;
  assign _EVAL_73 = {1'b0,$signed(_EVAL_220)};
  assign _EVAL_131 = _EVAL_6 == 3'h4;
  assign _EVAL_211 = _EVAL_182 | _EVAL_11;
  assign _EVAL_269 = _EVAL_14 <= 3'h6;
  assign _EVAL_283 = _EVAL_5 == _EVAL_35;
  assign _EVAL_140 = _EVAL_9 & _EVAL_224;
  assign _EVAL_82 = ~_EVAL_164;
  assign _EVAL_185 = _EVAL_14 == 3'h1;
  assign _EVAL_65 = _EVAL_273 | _EVAL_11;
  assign _EVAL_212 = ~_EVAL_306;
  assign _EVAL_233 = 2'h1 << _EVAL_32;
  assign _EVAL_236 = _EVAL_5[4:3];
  assign _EVAL_291 = ~_EVAL_203;
  assign _EVAL_146 = ~_EVAL_114;
  assign _EVAL_114 = _EVAL_64 | _EVAL_11;
  assign _EVAL_142 = _EVAL_109 | _EVAL_11;
  assign _EVAL_297 = ~_EVAL_271;
  assign _EVAL_174 = _EVAL_111 & _EVAL_226;
  assign _EVAL_279 = _EVAL_233 | 2'h1;
  assign _EVAL_219 = ~_EVAL_195;
  assign _EVAL_156 = ~_EVAL_102;
  assign _EVAL_40 = ~_EVAL_77;
  assign _EVAL_109 = _EVAL_4 == _EVAL_71;
  assign _EVAL_118 = _EVAL_14 == 3'h5;
  assign _EVAL_98 = _EVAL_315 | _EVAL_11;
  assign _EVAL_81 = _EVAL_158 == 31'h0;
  assign _EVAL_25 = _EVAL_5 == 5'h11;
  assign _EVAL_284 = ~_EVAL_261;
  assign _EVAL_202 = _EVAL_77 & _EVAL_195;
  assign _EVAL_311 = _EVAL_242 | _EVAL_11;
  assign _EVAL_198 = 3'h6 == _EVAL_0;
  assign _EVAL_33 = _EVAL_87 | _EVAL_11;
  assign _EVAL_50 = ~_EVAL_100;
  assign _EVAL_182 = _EVAL_16 == _EVAL_214;
  assign _EVAL_120 = _EVAL_194 - 4'h1;
  assign _EVAL_86 = ~_EVAL_301;
  assign _EVAL_31 = _EVAL_40 & _EVAL_195;
  assign _EVAL_137 = plusarg_reader_out == 32'h0;
  assign _EVAL_173 = _EVAL_244 >> _EVAL_4;
  assign _EVAL_267 = _EVAL_125 ? _EVAL_160 : 32'h0;
  assign _EVAL_22 = ~_EVAL_129;
  assign _EVAL_238 = _EVAL_250 | _EVAL_101;
  assign _EVAL_216 = ~_EVAL_141;
  assign _EVAL_19 = _EVAL_288 | _EVAL_244;
  assign _EVAL_70 = ~_EVAL_24;
  assign _EVAL_93 = _EVAL_277 | _EVAL_11;
  assign _EVAL_110 = _EVAL_81 | _EVAL_11;
  assign _EVAL_59 = ~_EVAL_299;
  assign _EVAL_170 = _EVAL_173[0];
  assign _EVAL_92 = _EVAL_300 | _EVAL_309;
  assign _EVAL_196 = _EVAL_6 == 3'h6;
  assign _EVAL_24 = _EVAL_248 | _EVAL_11;
  assign _EVAL_97 = ~_EVAL_231;
  assign _EVAL_301 = _EVAL_26 | _EVAL_11;
  assign _EVAL_96 = _EVAL_5 == 5'h8;
  assign _EVAL_205 = _EVAL_194 == 4'h0;
  assign _EVAL_287 = _EVAL_236 == 2'h0;
  assign _EVAL_63 = _EVAL_147 & _EVAL_205;
  assign _EVAL_250 = _EVAL_4 == 5'h11;
  assign _EVAL_259 = _EVAL_8 == _EVAL_80;
  assign _EVAL_256 = _EVAL_1 == _EVAL_227;
  assign _EVAL_178 = _EVAL_263 | _EVAL_30;
  assign _EVAL_39 = _EVAL_120[3:0];
  assign _EVAL_163 = ~_EVAL_154;
  assign _EVAL_239 = _EVAL_238 | _EVAL_314;
  assign _EVAL_241 = _EVAL_40 & _EVAL_219;
  assign _EVAL_278 = ~_EVAL_93;
  assign _EVAL_234 = _EVAL_295 == 4'h0;
  assign _EVAL_294 = _EVAL_6 == 3'h5;
  assign _EVAL_306 = _EVAL_283 | _EVAL_11;
  assign _EVAL_298 = _EVAL_8 >= 3'h2;
  assign _EVAL_121 = ~_EVAL_88;
  assign _EVAL_223 = ~_EVAL_65;
  assign _EVAL_45 = _EVAL_9 & _EVAL_232;
  assign _EVAL_203 = _EVAL_138 | _EVAL_11;
  assign _EVAL_54 = _EVAL_292[3:0];
  assign _EVAL_264 = ~_EVAL_257;
  assign _EVAL_183 = _EVAL_217 & _EVAL_108;
  assign _EVAL_312 = ~_EVAL_235;
  assign _EVAL_184 = _EVAL_148 < plusarg_reader_out;
  assign _EVAL_21 = _EVAL_234 | _EVAL_11;
  assign _EVAL_235 = _EVAL_240 | _EVAL_11;
  assign _EVAL_166 = _EVAL_148 + 32'h1;
  assign _EVAL_102 = |_EVAL_288;
  assign _EVAL_58 = _EVAL_92 | _EVAL_41;
  assign _EVAL_126 = _EVAL_18 != 3'h0;
  assign _EVAL_315 = _EVAL_12 == _EVAL_253;
  assign _EVAL_101 = _EVAL_4 == 5'h10;
  assign _EVAL_141 = _EVAL_126 | _EVAL_11;
  assign _EVAL_160 = 32'h1 << _EVAL_5;
  assign _EVAL_20 = _EVAL_9 & _EVAL_294;
  assign _EVAL_36 = _EVAL_9 & _EVAL_196;
  assign _EVAL_132 = ~_EVAL_153;
  assign _EVAL_171 = _EVAL_9 & _EVAL_131;
  assign _EVAL_127 = ~_EVAL_255;
  assign _EVAL_41 = _EVAL_281 & _EVAL_44;
  assign _EVAL_90 = _EVAL_230 | _EVAL_249;
  assign _EVAL_190 = _EVAL_18 <= 3'h2;
  assign _EVAL_43 = ~_EVAL_13;
  assign _EVAL_248 = _EVAL_18 <= 3'h3;
  assign _EVAL_270 = _EVAL_18 <= 3'h4;
  assign _EVAL_186 = ~_EVAL_179;
  assign _EVAL_242 = _EVAL_111 | _EVAL_61;
  assign _EVAL_249 = _EVAL_287 & _EVAL_99;
  assign _EVAL_26 = ~_EVAL_170;
  assign _EVAL_66 = _EVAL_133 <= 3'h6;
  assign _EVAL_266 = ~_EVAL_189;
  assign _EVAL_83 = _EVAL_4 == 5'h8;
  assign _EVAL_37 = _EVAL_3 & _EVAL_215;
  assign _EVAL_72 = ~_EVAL_144;
  assign _EVAL_305 = ~_EVAL_188;
  assign _EVAL_285 = _EVAL_14 == _EVAL_89;
  assign _EVAL_277 = _EVAL_10 != 2'h2;
  assign _EVAL_135 = ~_EVAL_142;
  assign _EVAL_230 = _EVAL_25 | _EVAL_206;
  assign _EVAL_208 = _EVAL_263 | _EVAL_192;
  assign _EVAL_95 = ~_EVAL_280;
  assign _EVAL_129 = _EVAL_79 | _EVAL_11;
  assign _EVAL_27 = _EVAL_50 | _EVAL_137;
  assign _EVAL_299 = _EVAL_112 | _EVAL_11;
  assign _EVAL_112 = _EVAL_152 == 4'h0;
  assign _EVAL_220 = _EVAL_1 ^ 31'h40000000;
  assign _EVAL_197 = _EVAL_43 | _EVAL_17;
  assign _EVAL_147 = _EVAL_7 & _EVAL_9;
  assign _EVAL_189 = _EVAL_209 == 4'h0;
  assign _EVAL_84 = $signed(_EVAL_73) & -32'sh2000;
  assign _EVAL_143 = $signed(_EVAL_265) == 32'sh0;
  assign _EVAL_79 = _EVAL_139[0];
  assign _EVAL_257 = _EVAL_169 | _EVAL_11;
  assign _EVAL_57 = _EVAL_174 | _EVAL_11;
  assign _EVAL_187 = 32'h1 << _EVAL_4;
  assign _EVAL_78 = _EVAL_175[3:0];
  assign _EVAL_159 = _EVAL_6 == 3'h2;
  assign _EVAL_113 = ~_EVAL_251;
  assign _EVAL_290 = _EVAL_6 == 3'h3;
  assign _EVAL_309 = _EVAL_150 & _EVAL_77;
  assign _EVAL_292 = _EVAL_209 - 4'h1;
  assign _EVAL_217 = _EVAL_2 & _EVAL_3;
  assign _EVAL_288 = _EVAL_228[17:0];
  assign _EVAL_167 = _EVAL_67 | _EVAL_156;
  assign _EVAL_271 = _EVAL_285 | _EVAL_11;
  assign _EVAL_317 = _EVAL_4[4:3];
  assign _EVAL_172 = _EVAL_10 == _EVAL_74;
  assign _EVAL_175 = _EVAL_49 - 4'h1;
  assign _EVAL_286 = _EVAL_217 & _EVAL_189;
  assign _EVAL_275 = ~_EVAL_293;
  assign _EVAL_195 = _EVAL_1[0];
  assign _EVAL_215 = _EVAL_14 == 3'h4;
  assign _EVAL_28 = _EVAL_18 == _EVAL_48;
  assign _EVAL_52 = ~_EVAL_98;
  assign _EVAL_94 = _EVAL_117[5:2];
  assign _EVAL_61 = _EVAL_198 & _EVAL_83;
  assign _EVAL_214 = {_EVAL_104,_EVAL_58,_EVAL_178,_EVAL_208};
  assign _EVAL_207 = _EVAL_3 & _EVAL_316;
  assign _EVAL_210 = _EVAL_3 & _EVAL_118;
  assign _EVAL_201 = ~_EVAL_211;
  assign _EVAL_193 = _EVAL_10 <= 2'h2;
  assign _EVAL_133 = _EVAL_4[2:0];
  assign _EVAL_262 = _EVAL_105 | _EVAL_11;
  assign _EVAL_106 = ~_EVAL_252;
  assign _EVAL_42 = _EVAL_3 & _EVAL_185;
  assign _EVAL_303 = _EVAL_9 & _EVAL_47;
  assign _EVAL_168 = _EVAL_9 & _EVAL_159;
  assign _EVAL_77 = _EVAL_1[1];
  assign _EVAL_60 = ~_EVAL_116;
  assign _EVAL_157 = 13'h3f << _EVAL_8;
  assign _EVAL_300 = _EVAL_0 >= 3'h2;
  assign _EVAL_151 = _EVAL_14 == 3'h2;
  assign _EVAL_314 = _EVAL_245 & _EVAL_66;
  assign _EVAL_280 = _EVAL_256 | _EVAL_11;
  assign _EVAL_268 = _EVAL_147 | _EVAL_217;
  assign _EVAL_302 = ~_EVAL_308;
  assign _EVAL_62 = _EVAL_29[5:0];
  assign _EVAL_144 = _EVAL_122 | _EVAL_11;
  assign _EVAL_164 = _EVAL_190 | _EVAL_11;
  assign _EVAL_134 = _EVAL_6 == _EVAL_247;
  assign _EVAL_152 = ~_EVAL_16;
  assign _EVAL_32 = _EVAL_0[0];
  assign _EVAL_176 = _EVAL_5[2:0];
  assign _EVAL_293 = _EVAL_49 == 4'h0;
  assign _EVAL_153 = _EVAL_157[5:0];
  assign _EVAL_130 = ~_EVAL_214;
  assign _EVAL_91 = ~_EVAL_128;
  assign _EVAL_67 = _EVAL_288 != _EVAL_38;
  assign _EVAL_154 = _EVAL_134 | _EVAL_11;
  assign _EVAL_38 = _EVAL_267[17:0];
  assign _EVAL_105 = ~_EVAL;
  assign _EVAL_123 = ~_EVAL_57;
  assign _EVAL_128 = _EVAL_167 | _EVAL_11;
  assign _EVAL_104 = _EVAL_92 | _EVAL_204;
  assign _EVAL_289 = _EVAL_43 | _EVAL_11;
  assign _EVAL_191 = ~_EVAL_33;
  assign _EVAL_200 = _EVAL_115 & _EVAL_254;
  assign _EVAL_181 = ~_EVAL_311;
  assign _EVAL_47 = _EVAL_6 == 3'h7;
  assign _EVAL_150 = _EVAL_279[1];
  assign _EVAL_261 = _EVAL_269 | _EVAL_11;
  assign _EVAL_265 = _EVAL_84;
  assign _EVAL_243 = _EVAL_244 | _EVAL_288;
  assign _EVAL_308 = _EVAL_172 | _EVAL_11;
  assign _EVAL_99 = _EVAL_176 <= 3'h6;
  assign _EVAL_229 = _EVAL_239 | _EVAL_83;
  assign _EVAL_88 = _EVAL_298 | _EVAL_11;
  assign _EVAL_29 = 13'h3f << _EVAL_0;
  assign _EVAL_237 = {{25'd0}, _EVAL_117};
  assign _EVAL_139 = _EVAL_19 >> _EVAL_5;
  assign _EVAL_296 = ~_EVAL_282;
  assign _EVAL_30 = _EVAL_281 & _EVAL_31;
  assign _EVAL_119 = ~_EVAL_316;
  assign _EVAL_281 = _EVAL_279[0];
  assign _EVAL_179 = _EVAL_6[2];
  assign _EVAL_169 = _EVAL_18 <= 3'h1;
  assign _EVAL_316 = _EVAL_14 == 3'h6;
  assign _EVAL_251 = _EVAL_197 | _EVAL_11;
  always @(posedge _EVAL_15) begin
    if (_EVAL_286) begin
      _EVAL_35 <= _EVAL_5;
    end
    if (_EVAL_213) begin
      _EVAL_48 <= _EVAL_18;
    end
    if (_EVAL_11) begin
      _EVAL_49 <= 4'h0;
    end else if (_EVAL_147) begin
      if (_EVAL_293) begin
        if (_EVAL_186) begin
          _EVAL_49 <= _EVAL_94;
        end else begin
          _EVAL_49 <= 4'h0;
        end
      end else begin
        _EVAL_49 <= _EVAL_78;
      end
    end
    if (_EVAL_213) begin
      _EVAL_71 <= _EVAL_4;
    end
    if (_EVAL_286) begin
      _EVAL_74 <= _EVAL_10;
    end
    if (_EVAL_286) begin
      _EVAL_80 <= _EVAL_8;
    end
    if (_EVAL_286) begin
      _EVAL_89 <= _EVAL_14;
    end
    if (_EVAL_11) begin
      _EVAL_107 <= 4'h0;
    end else if (_EVAL_217) begin
      if (_EVAL_108) begin
        if (_EVAL_75) begin
          _EVAL_107 <= _EVAL_310;
        end else begin
          _EVAL_107 <= 4'h0;
        end
      end else begin
        _EVAL_107 <= _EVAL_246;
      end
    end
    if (_EVAL_11) begin
      _EVAL_148 <= 32'h0;
    end else if (_EVAL_268) begin
      _EVAL_148 <= 32'h0;
    end else begin
      _EVAL_148 <= _EVAL_76;
    end
    if (_EVAL_11) begin
      _EVAL_194 <= 4'h0;
    end else if (_EVAL_147) begin
      if (_EVAL_205) begin
        if (_EVAL_186) begin
          _EVAL_194 <= _EVAL_94;
        end else begin
          _EVAL_194 <= 4'h0;
        end
      end else begin
        _EVAL_194 <= _EVAL_39;
      end
    end
    if (_EVAL_11) begin
      _EVAL_209 <= 4'h0;
    end else if (_EVAL_217) begin
      if (_EVAL_189) begin
        if (_EVAL_75) begin
          _EVAL_209 <= _EVAL_310;
        end else begin
          _EVAL_209 <= 4'h0;
        end
      end else begin
        _EVAL_209 <= _EVAL_54;
      end
    end
    if (_EVAL_213) begin
      _EVAL_227 <= _EVAL_1;
    end
    if (_EVAL_11) begin
      _EVAL_244 <= 18'h0;
    end else begin
      _EVAL_244 <= _EVAL_124;
    end
    if (_EVAL_213) begin
      _EVAL_247 <= _EVAL_6;
    end
    if (_EVAL_286) begin
      _EVAL_253 <= _EVAL_12;
    end
    if (_EVAL_213) begin
      _EVAL_272 <= _EVAL_0;
    end
    if (_EVAL_286) begin
      _EVAL_274 <= _EVAL_13;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_297) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8511366d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_302) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21d22f63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5daa0c22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d02c6f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_82) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_91) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_125 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b8fba4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a418621b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_86) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4876c31f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(163eca24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b82adea8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee4c901c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f302751f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d4ef079)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6174b75b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_297) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_52) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49091f92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee1a58cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_313) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d42834e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa5a9e2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34afdc24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b4b658c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c50ba1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(796b6f9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(994dfc52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5be892de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b352bfb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22fe522)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e1736a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(601dd246)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_70) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4eedcdd3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c47e6b1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_302) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(364a800a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(854952e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db55e2dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32131e37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3 & _EVAL_284) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf763808)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_212) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d788c4a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ac03027)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc249c75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f466f2f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db1db333)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_63 & _EVAL_86) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(820e378e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(942b6c96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_264) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a171b1f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(584e0880)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_82) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42d82d5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96628356)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e1736a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4526ca79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33c3102e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61ea17c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32566319)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5c7557d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43b7a47d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_291) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58e92c24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(374b3043)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_163) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b917b5b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_313) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23c05b08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(726362c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5fa21c2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_127) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b10a64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_291) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17ad5215)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98136390)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_177) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24b3c96f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3415335e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a667175)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf3107e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8950cde)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(648b2cff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5241695b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b63e18b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_305) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e47ccd94)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_191) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d589030)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_127) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7901ed44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35e89537)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89a1945d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1605db99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_305) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(746c7e4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af8463bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_60) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(668965a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f53a66b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_276) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6da1188)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_264) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(401389d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acc40d74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13330877)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_70) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53d5d707)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_163) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5979940a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9274a69e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_161 & _EVAL_191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26c0d121)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10f4890c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_60) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6fe2bdd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_171 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f87c2ef8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a6baff8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61e11f5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_52) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36 & _EVAL_276) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8d2a4e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_212) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64d7b289)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_168 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_45 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_210 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42753c52)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_42 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f160cab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_177) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_3 & _EVAL_284) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_303 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_35 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_48 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_49 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_71 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_74 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_80 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_89 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_107 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_148 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_194 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_209 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_227 = _RAND_11[30:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_244 = _RAND_12[17:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_247 = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_253 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_272 = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_274 = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
