//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_3(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  output [3:0]  _EVAL_2,
  output        _EVAL_3,
  output [3:0]  _EVAL_4,
  input  [3:0]  _EVAL_5,
  input  [3:0]  _EVAL_6,
  output        _EVAL_7,
  output [31:0] _EVAL_8,
  input  [2:0]  _EVAL_9,
  input         _EVAL_10,
  input  [2:0]  _EVAL_11,
  output        _EVAL_12,
  output        _EVAL_13,
  input         _EVAL_14,
  output [2:0]  _EVAL_15,
  input  [31:0] _EVAL_16,
  output [31:0] _EVAL_17,
  input  [31:0] _EVAL_18,
  output [2:0]  _EVAL_19,
  input  [2:0]  _EVAL_20,
  input  [1:0]  _EVAL_21,
  output        _EVAL_22,
  output [31:0] _EVAL_23,
  output        _EVAL_24,
  output [31:0] _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  output        _EVAL_28,
  input  [3:0]  _EVAL_29,
  input         _EVAL_30,
  input  [1:0]  _EVAL_31,
  input         _EVAL_32,
  output        _EVAL_33,
  input         _EVAL_34,
  output        _EVAL_35,
  input         _EVAL_36,
  output        _EVAL_37,
  output [4:0]  _EVAL_38,
  input         _EVAL_39,
  output [2:0]  _EVAL_40,
  output        _EVAL_41,
  input         _EVAL_42,
  input         _EVAL_43,
  output        _EVAL_44,
  output        _EVAL_45,
  output        _EVAL_46,
  output [30:0] _EVAL_47,
  input         _EVAL_48,
  output        _EVAL_49,
  input  [4:0]  _EVAL_50,
  output [2:0]  _EVAL_51,
  input  [4:0]  _EVAL_52,
  input  [31:0] _EVAL_53,
  input  [2:0]  _EVAL_54,
  output        _EVAL_55,
  input  [2:0]  _EVAL_56,
  input         _EVAL_57,
  input  [2:0]  _EVAL_58,
  output        _EVAL_59,
  output [3:0]  _EVAL_60,
  input         _EVAL_61,
  output        _EVAL_62,
  output        _EVAL_63,
  input         _EVAL_64,
  output        _EVAL_65,
  output [2:0]  _EVAL_66,
  output        _EVAL_67,
  input         _EVAL_68,
  input         _EVAL_69,
  input  [3:0]  _EVAL_70,
  input         _EVAL_71,
  input         _EVAL_72,
  output [1:0]  _EVAL_73,
  input         _EVAL_74,
  input         _EVAL_75,
  output [3:0]  _EVAL_76,
  input         _EVAL_77,
  input  [2:0]  _EVAL_78,
  output [31:0] _EVAL_79,
  input  [3:0]  _EVAL_80,
  output [2:0]  _EVAL_81,
  input  [31:0] _EVAL_82,
  output        _EVAL_83,
  output [2:0]  _EVAL_84,
  output [3:0]  _EVAL_85,
  output        _EVAL_86,
  input         _EVAL_87,
  output [4:0]  _EVAL_88,
  input         _EVAL_89,
  output        _EVAL_90,
  input  [3:0]  _EVAL_91,
  output [1:0]  _EVAL_92,
  output        _EVAL_93,
  input  [31:0] _EVAL_94,
  output [3:0]  _EVAL_95,
  input  [31:0] _EVAL_96
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  wire [3:0] _EVAL_97;
  wire [3:0] _EVAL_99;
  wire [3:0] _EVAL_100;
  wire [32:0] _EVAL_102;
  wire  _EVAL_103;
  wire [3:0] _EVAL_105;
  wire [5:0] _EVAL_106;
  wire  _EVAL_107;
  wire [1:0] _EVAL_109;
  wire  _EVAL_110;
  wire [7:0] _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire [6:0] _EVAL_116;
  wire [32:0] _EVAL_117;
  wire [2:0] _EVAL_119;
  wire [1:0] _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire [1:0] _EVAL_124;
  wire [3:0] _EVAL_126;
  wire [7:0] _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_130;
  wire [6:0] _EVAL_131;
  wire [1:0] _EVAL_135;
  wire [31:0] _EVAL_136;
  wire [3:0] _EVAL_139;
  reg  _EVAL_140;
  wire [2:0] _EVAL_141;
  wire [2:0] _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire [31:0] _EVAL_145;
  wire [1:0] _EVAL_146;
  wire [4:0] _EVAL_147;
  wire  _EVAL_148;
  wire [31:0] _EVAL_149;
  wire [2:0] _EVAL_150;
  wire [3:0] _EVAL_151;
  wire [2:0] _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire [1:0] _EVAL_159;
  wire [1:0] _EVAL_160;
  wire  _EVAL_161;
  reg [1:0] _EVAL_162;
  reg [5:0] _EVAL_163;
  wire [2:0] _EVAL_164;
  wire [32:0] _EVAL_165;
  wire [32:0] _EVAL_166;
  wire  _EVAL_167;
  wire [3:0] _EVAL_168;
  wire [3:0] _EVAL_169;
  wire [5:0] _EVAL_170;
  wire [3:0] _EVAL_171;
  wire  _EVAL_172;
  wire [4:0] _EVAL_173;
  wire  _EVAL_174;
  wire [4:0] _EVAL_175;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire [2:0] _EVAL_181;
  wire [31:0] _EVAL_183;
  wire [3:0] _EVAL_185;
  wire [4:0] _EVAL_186;
  wire [1:0] _EVAL_187;
  wire [4:0] _EVAL_188;
  wire [1:0] _EVAL_189;
  wire  _EVAL_190;
  wire [6:0] _EVAL_191;
  wire [1:0] _EVAL_192;
  wire  _EVAL_193;
  wire [1:0] _EVAL_194;
  wire  _EVAL_195;
  wire [3:0] _EVAL_196;
  wire  _EVAL_197;
  reg  _EVAL_198;
  wire [1:0] _EVAL_199;
  wire [3:0] _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire [2:0] _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_208;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire [5:0] _EVAL_213;
  wire [5:0] _EVAL_214;
  wire  _EVAL_215;
  wire [5:0] _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire [31:0] _EVAL_221;
  wire [3:0] _EVAL_222;
  wire  _EVAL_223;
  wire [3:0] _EVAL_224;
  wire [5:0] _EVAL_225;
  wire  _EVAL_227;
  wire [3:0] _EVAL_229;
  wire [3:0] _EVAL_230;
  wire [3:0] _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire [32:0] _EVAL_234;
  wire  _EVAL_236;
  wire [5:0] _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  reg [1:0] _EVAL_240;
  wire [5:0] _EVAL_241;
  wire [3:0] _EVAL_242;
  wire [3:0] _EVAL_243;
  wire [3:0] _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire [31:0] _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire [7:0] _EVAL_250;
  wire [1:0] _EVAL_251;
  wire [1:0] _EVAL_252;
  wire [3:0] _EVAL_254;
  wire  _EVAL_255;
  wire [5:0] _EVAL_256;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire [5:0] _EVAL_262;
  wire [3:0] _EVAL_263;
  wire  _EVAL_264;
  wire [2:0] _EVAL_265;
  wire [31:0] _EVAL_266;
  wire [5:0] _EVAL_267;
  wire  _EVAL_268;
  wire [4:0] _EVAL_269;
  wire  _EVAL_270;
  wire [1:0] _EVAL_271;
  wire  _EVAL_272;
  reg [1:0] _EVAL_273;
  wire  _EVAL_275;
  wire [5:0] _EVAL_276;
  wire [1:0] _EVAL_277;
  wire [7:0] _EVAL_279;
  wire [5:0] _EVAL_281;
  wire [1:0] _EVAL_282;
  wire [5:0] _EVAL_283;
  wire  _EVAL_284;
  wire [2:0] _EVAL_287;
  wire [4:0] _EVAL_288;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire [5:0] _EVAL_294;
  wire [3:0] _EVAL_296;
  wire  _EVAL_297;
  reg [5:0] _EVAL_298;
  reg  _EVAL_299;
  wire [1:0] _EVAL_300;
  wire  _EVAL_301;
  wire [31:0] _EVAL_303;
  wire [5:0] _EVAL_304;
  wire [31:0] _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_307;
  wire [2:0] _EVAL_308;
  wire [32:0] _EVAL_309;
  wire  _EVAL_310;
  wire  _EVAL_311;
  wire  _EVAL_312;
  wire [3:0] _EVAL_313;
  wire  _EVAL_314;
  wire [4:0] _EVAL_315;
  wire [3:0] _EVAL_316;
  wire  _EVAL_317;
  wire [1:0] _EVAL_318;
  wire [3:0] _EVAL_319;
  wire  _EVAL_320;
  reg [5:0] _EVAL_321;
  wire [1:0] _EVAL_322;
  wire [7:0] _EVAL_323;
  wire [31:0] _EVAL_324;
  wire [1:0] _EVAL_325;
  wire [4:0] _EVAL_326;
  wire [6:0] _EVAL_329;
  wire  _EVAL_330;
  wire [3:0] _EVAL_331;
  wire  _EVAL_332;
  wire [5:0] _EVAL_333;
  wire  _EVAL_334;
  wire [1:0] _EVAL_335;
  wire [2:0] _EVAL_336;
  wire [2:0] _EVAL_337;
  reg [1:0] _EVAL_338;
  wire [2:0] _EVAL_339;
  wire  _EVAL_340;
  wire [3:0] _EVAL_341;
  wire  _EVAL_342;
  wire [32:0] _EVAL_343;
  wire [1:0] _EVAL_345;
  wire [1:0] _EVAL_346;
  wire [7:0] _EVAL_347;
  reg  _EVAL_348;
  wire [5:0] _EVAL_349;
  wire  _EVAL_351;
  wire [1:0] _EVAL_352;
  wire  _EVAL_354;
  wire [1:0] _EVAL_356;
  wire  _EVAL_357;
  wire  _EVAL_358;
  wire [20:0] _EVAL_359;
  wire  _EVAL_361;
  wire  _EVAL_363;
  wire [2:0] _EVAL_364;
  wire  _EVAL_365;
  wire  _EVAL_366;
  wire  _EVAL_367;
  wire  _EVAL_368;
  wire [3:0] _EVAL_369;
  wire  _EVAL_370;
  wire  _EVAL_371;
  wire [22:0] _EVAL_372;
  wire [3:0] _EVAL_373;
  wire [1:0] _EVAL_374;
  wire [1:0] _EVAL_375;
  wire [5:0] _EVAL_376;
  wire [1:0] _EVAL_377;
  wire [4:0] _EVAL_378;
  wire [31:0] _EVAL_379;
  wire  _EVAL_380;
  wire  _EVAL_381;
  wire  _EVAL_382;
  wire [2:0] _EVAL_383;
  wire  _EVAL_384;
  wire  _EVAL_385;
  wire [5:0] _EVAL_386;
  wire  _EVAL_388;
  wire [1:0] _EVAL_389;
  wire [5:0] _EVAL_391;
  wire  _EVAL_392;
  wire  _EVAL_394;
  reg [5:0] _EVAL_395;
  reg  _EVAL_396;
  wire  _EVAL_397;
  wire  _EVAL_398;
  wire [22:0] _EVAL_399;
  wire [1:0] _EVAL_400;
  wire  _EVAL_401;
  wire [31:0] _EVAL_402;
  wire  _EVAL_403;
  wire [31:0] _EVAL_405;
  wire  _EVAL_406;
  wire [2:0] _EVAL_407;
  wire  _EVAL_408;
  wire [1:0] _EVAL_409;
  wire [1:0] _EVAL_412;
  wire [2:0] _EVAL_414;
  wire [3:0] _EVAL_415;
  reg  _EVAL_416;
  wire  _EVAL_417;
  wire [5:0] _EVAL_418;
  wire [31:0] _EVAL_419;
  wire [2:0] _EVAL_421;
  wire  _EVAL_422;
  wire [32:0] _EVAL_423;
  wire  _EVAL_424;
  wire  _EVAL_425;
  wire [2:0] _EVAL_426;
  wire [5:0] _EVAL_427;
  wire  _EVAL_428;
  wire  _EVAL_429;
  wire [1:0] _EVAL_430;
  wire  _EVAL_431;
  wire [1:0] _EVAL_433;
  wire  _EVAL_434;
  wire [5:0] _EVAL_435;
  wire [4:0] _EVAL_436;
  wire [3:0] _EVAL_437;
  wire [22:0] _EVAL_438;
  wire [32:0] _EVAL_439;
  wire  _EVAL_440;
  wire [5:0] _EVAL_441;
  wire  _EVAL_443;
  wire [3:0] _EVAL_444;
  wire  _EVAL_445;
  wire [3:0] _EVAL_447;
  wire [3:0] _EVAL_448;
  wire  _EVAL_449;
  wire [32:0] _EVAL_450;
  wire [3:0] _EVAL_451;
  wire [5:0] _EVAL_452;
  wire  _EVAL_453;
  wire  _EVAL_454;
  wire  _EVAL_455;
  wire [32:0] _EVAL_456;
  wire [31:0] _EVAL_457;
  wire [3:0] _EVAL_458;
  wire [4:0] _EVAL_459;
  wire  _EVAL_460;
  wire [1:0] _EVAL_461;
  wire [1:0] _EVAL_462;
  wire [3:0] _EVAL_463;
  wire  _EVAL_465;
  wire  _EVAL_466;
  wire [4:0] _EVAL_467;
  wire [3:0] _EVAL_468;
  wire  _EVAL_469;
  wire  _EVAL_470;
  wire [5:0] _EVAL_471;
  wire [2:0] _EVAL_472;
  wire [5:0] _EVAL_473;
  wire [1:0] _EVAL_474;
  reg  _EVAL_475;
  wire [2:0] _EVAL_476;
  wire [1:0] _EVAL_477;
  wire [3:0] _EVAL_478;
  reg  _EVAL_479;
  wire  _EVAL_480;
  wire [1:0] _EVAL_481;
  wire  _EVAL_482;
  wire  _EVAL_483;
  wire  _EVAL_484;
  wire  _EVAL_485;
  wire [32:0] _EVAL_486;
  wire  _EVAL_487;
  wire [3:0] _EVAL_488;
  wire  _EVAL_489;
  wire  _EVAL_490;
  wire [1:0] _EVAL_491;
  wire  _EVAL_492;
  wire [2:0] _EVAL_493;
  wire [3:0] _EVAL_496;
  wire [1:0] _EVAL_498;
  wire  _EVAL_499;
  wire  _EVAL_500;
  wire [3:0] _EVAL_501;
  wire  _EVAL_502;
  wire [1:0] _EVAL_503;
  wire [2:0] _EVAL_504;
  wire  _EVAL_505;
  wire  _EVAL_506;
  wire  _EVAL_507;
  wire [1:0] _EVAL_508;
  wire  _EVAL_509;
  wire  _EVAL_510;
  assign _EVAL_2 = _EVAL_448 | _EVAL_415;
  assign _EVAL_86 = _EVAL_179 | _EVAL_128;
  assign _EVAL_156 = _EVAL_284 ? _EVAL_232 : _EVAL_429;
  assign _EVAL_227 = _EVAL_507 | _EVAL_445;
  assign _EVAL_144 = _EVAL_203 & _EVAL_77;
  assign _EVAL_458 = {{1'd0}, _EVAL_152};
  assign _EVAL_347 = ~_EVAL_250;
  assign _EVAL_249 = _EVAL_367 ? _EVAL_492 : _EVAL_416;
  assign _EVAL_181 = _EVAL_203 ? _EVAL_58 : 3'h0;
  assign _EVAL_488 = _EVAL_485 ? _EVAL_80 : 4'h0;
  assign _EVAL_277 = _EVAL_187 | _EVAL_430;
  assign _EVAL_254 = _EVAL_99 | _EVAL_341;
  assign _EVAL_324 = _EVAL_408 ? _EVAL_82 : 32'h0;
  assign _EVAL_304 = {{2'd0}, _EVAL_463};
  assign _EVAL_206 = _EVAL_121 & _EVAL_246;
  assign _EVAL_45 = _EVAL_422 | _EVAL_434;
  assign _EVAL_46 = _EVAL_307 | _EVAL_197;
  assign _EVAL_239 = _EVAL_311 & _EVAL_490;
  assign _EVAL_503 = _EVAL_468[1:0];
  assign _EVAL_272 = _EVAL_284 ? _EVAL_121 : _EVAL_198;
  assign _EVAL_84 = _EVAL_308 | _EVAL_493;
  assign _EVAL_232 = _EVAL_394 | _EVAL_246;
  assign _EVAL_208 = _EVAL_26 & _EVAL_215;
  assign _EVAL_28 = _EVAL_233 | _EVAL_483;
  assign _EVAL_510 = $signed(_EVAL_439) == 33'sh0;
  assign _EVAL_213 = _EVAL_492 ? _EVAL_281 : 6'h0;
  assign _EVAL_368 = _EVAL_112 & _EVAL_71;
  assign _EVAL_122 = _EVAL_148 & _EVAL_71;
  assign _EVAL_294 = _EVAL_111[7:2];
  assign _EVAL_135 = _EVAL_148 ? _EVAL_21 : 2'h0;
  assign _EVAL_367 = _EVAL_298 == 6'h0;
  assign _EVAL_454 = ~_EVAL_260;
  assign _EVAL_225 = {{5'd0}, _EVAL_238};
  assign _EVAL_301 = _EVAL_245 & _EVAL_113;
  assign _EVAL_484 = _EVAL_27 & _EVAL_174;
  assign _EVAL_243 = {_EVAL_325,_EVAL_202,_EVAL_489};
  assign _EVAL_41 = _EVAL_220 ? _EVAL_264 : _EVAL_330;
  assign _EVAL_234 = {1'b0,$signed(_EVAL_145)};
  assign _EVAL_508 = _EVAL_478[1:0];
  assign _EVAL_22 = _EVAL_431 | _EVAL_223;
  assign _EVAL_424 = _EVAL_193 & _EVAL_87;
  assign _EVAL_429 = _EVAL_354 | _EVAL_317;
  assign _EVAL_223 = _EVAL_312 & _EVAL_30;
  assign _EVAL_308 = _EVAL_485 ? _EVAL_78 : 3'h0;
  assign _EVAL_419 = _EVAL_203 ? _EVAL_16 : 32'h0;
  assign _EVAL_474 = {_EVAL_484,_EVAL_465};
  assign _EVAL_427 = _EVAL_167 ? _EVAL_294 : 6'h0;
  assign _EVAL_158 = |_EVAL_409;
  assign _EVAL_23 = _EVAL_402 | _EVAL_379;
  assign _EVAL_25 = _EVAL_303 | _EVAL_183;
  assign _EVAL_109 = {_EVAL_202,_EVAL_489};
  assign _EVAL_40 = _EVAL_414 | _EVAL_119;
  assign _EVAL_486 = $signed(_EVAL_165) & 33'sh40000000;
  assign _EVAL_160 = _EVAL_474 & _EVAL_345;
  assign _EVAL_303 = _EVAL_193 ? _EVAL_96 : 32'h0;
  assign _EVAL_216 = _EVAL_267 | _EVAL_304;
  assign _EVAL_333 = _EVAL_347[7:2];
  assign _EVAL_287 = {_EVAL_199, 1'h0};
  assign _EVAL_88 = _EVAL_188 | _EVAL_175;
  assign _EVAL_340 = _EVAL_475 & _EVAL_465;
  assign _EVAL_248 = _EVAL_367 ? _EVAL_365 : _EVAL_416;
  assign _EVAL_349 = _EVAL_201 ? _EVAL_471 : 6'h0;
  assign _EVAL_244 = _EVAL_52[4:1];
  assign _EVAL_307 = _EVAL_193 & _EVAL_48;
  assign _EVAL_363 = _EVAL_477[0];
  assign _EVAL_461 = _EVAL_196[3:2];
  assign _EVAL_496 = _EVAL_437 | _EVAL_319;
  assign _EVAL_292 = _EVAL_284 & _EVAL_64;
  assign _EVAL_212 = _EVAL_180 & _EVAL_489;
  assign _EVAL_498 = _EVAL_193 ? _EVAL_31 : 2'h0;
  assign _EVAL_205 = {_EVAL_187, 1'h0};
  assign _EVAL_359 = 21'h3f << _EVAL_451;
  assign _EVAL_185 = {_EVAL_240, 2'h0};
  assign _EVAL_501 = _EVAL_241[5:2];
  assign _EVAL_102 = _EVAL_117;
  assign _EVAL_269 = _EVAL_312 ? _EVAL_467 : 5'h0;
  assign _EVAL_250 = _EVAL_438[7:0];
  assign _EVAL_378 = _EVAL_485 ? _EVAL_52 : 5'h0;
  assign _EVAL_168 = {{1'd0}, _EVAL_426};
  assign _EVAL_431 = _EVAL_203 & _EVAL_74;
  assign _EVAL_468 = _EVAL_126 | _EVAL_185;
  assign _EVAL_389 = _EVAL_352 | _EVAL_481;
  assign _EVAL_92 = _EVAL_374 | _EVAL_135;
  assign _EVAL_236 = _EVAL_9[2];
  assign _EVAL_259 = _EVAL_252[1];
  assign _EVAL_245 = $signed(_EVAL_102) == 33'sh0;
  assign _EVAL_241 = ~_EVAL_473;
  assign _EVAL_124 = _EVAL_496[1:0];
  assign _EVAL_315 = _EVAL_378 | _EVAL_147;
  assign _EVAL_265 = _EVAL_112 ? _EVAL_56 : 3'h0;
  assign _EVAL_472 = _EVAL_408 ? _EVAL_58 : 3'h0;
  assign _EVAL_377 = ~_EVAL_240;
  assign _EVAL_388 = $signed(_EVAL_456) == 33'sh0;
  assign _EVAL_3 = _EVAL_315[0];
  assign _EVAL_487 = |_EVAL_474;
  assign _EVAL_443 = _EVAL_64 & _EVAL_480;
  assign _EVAL_51 = _EVAL_171[2:0];
  assign _EVAL_112 = _EVAL_220 ? _EVAL_290 : _EVAL_348;
  assign _EVAL_270 = _EVAL_408 & _EVAL_14;
  assign _EVAL_449 = _EVAL_335[1];
  assign _EVAL_33 = _EVAL_157 | _EVAL_122;
  assign _EVAL_17 = _EVAL_419 | _EVAL_136;
  assign _EVAL_376 = _EVAL_106 | _EVAL_170;
  assign _EVAL_116 = _EVAL_395 - _EVAL_225;
  assign _EVAL_471 = _EVAL_279[7:2];
  assign _EVAL_175 = _EVAL_249 ? _EVAL_467 : 5'h0;
  assign _EVAL_12 = _EVAL_239 | _EVAL_110;
  assign _EVAL_352 = _EVAL_477 & _EVAL_409;
  assign _EVAL_371 = _EVAL_50[4];
  assign _EVAL_105 = _EVAL_408 ? _EVAL_70 : 4'h0;
  assign _EVAL_361 = _EVAL_252[0];
  assign _EVAL_507 = _EVAL_396 & _EVAL_275;
  assign _EVAL_142 = _EVAL_193 ? _EVAL_78 : 3'h0;
  assign _EVAL_131 = _EVAL_298 - _EVAL_237;
  assign _EVAL_399 = 23'hff << _EVAL_80;
  assign _EVAL_351 = _EVAL_249 & _EVAL_0;
  assign _EVAL_149 = _EVAL_408 ? _EVAL_16 : 32'h0;
  assign _EVAL_238 = _EVAL_39 & _EVAL_161;
  assign _EVAL_462 = _EVAL_196[1:0];
  assign _EVAL_106 = _EVAL_506 ? _EVAL_349 : 6'h0;
  assign _EVAL_430 = _EVAL_205[1:0];
  assign _EVAL_247 = _EVAL_249 ? _EVAL_18 : 32'h0;
  assign _EVAL_193 = _EVAL_220 ? _EVAL_332 : _EVAL_475;
  assign _EVAL_414 = _EVAL_408 ? _EVAL_9 : 3'h0;
  assign _EVAL_358 = _EVAL_408 & _EVAL_69;
  assign _EVAL_146 = _EVAL_364[1:0];
  assign _EVAL_314 = _EVAL_482 ? _EVAL_449 : _EVAL_140;
  assign _EVAL_334 = _EVAL_220 ? _EVAL_259 : _EVAL_348;
  assign _EVAL_275 = _EVAL_61 & _EVAL_245;
  assign _EVAL_436 = _EVAL_112 ? _EVAL_50 : 5'h0;
  assign _EVAL_222 = _EVAL_139 | _EVAL_458;
  assign _EVAL_49 = _EVAL_258 | _EVAL_153;
  assign _EVAL_47 = _EVAL_305[30:0];
  assign _EVAL_335 = ~_EVAL_433;
  assign _EVAL_103 = _EVAL_220 ? _EVAL_361 : _EVAL_475;
  assign _EVAL_279 = ~_EVAL_323;
  assign _EVAL_394 = _EVAL_72 & _EVAL_403;
  assign _EVAL_434 = _EVAL_312 & _EVAL_32;
  assign _EVAL_407 = _EVAL_243[3:1];
  assign _EVAL_143 = _EVAL_312 & _EVAL_0;
  assign _EVAL_342 = |_EVAL_159;
  assign _EVAL_490 = _EVAL_64 & _EVAL_272;
  assign _EVAL_139 = {_EVAL_160,_EVAL_484,_EVAL_465};
  assign _EVAL_8 = _EVAL_324 | _EVAL_457;
  assign _EVAL_332 = _EVAL_361 & _EVAL_465;
  assign _EVAL_153 = _EVAL_112 & _EVAL_42;
  assign _EVAL_300 = _EVAL_375 & _EVAL_503;
  assign _EVAL_375 = _EVAL_468[3:2];
  assign _EVAL_231 = _EVAL_249 ? _EVAL_29 : 4'h0;
  assign _EVAL_466 = _EVAL_403 & _EVAL_443;
  assign _EVAL_343 = {1'b0,$signed(_EVAL_266)};
  assign _EVAL_506 = _EVAL_363 & _EVAL_394;
  assign _EVAL_435 = _EVAL_212 ? _EVAL_427 : 6'h0;
  assign _EVAL_447 = _EVAL_203 ? _EVAL_5 : 4'h0;
  assign _EVAL_169 = _EVAL_312 ? _EVAL_91 : 4'h0;
  assign _EVAL_417 = _EVAL_440 & _EVAL_342;
  assign _EVAL_317 = _EVAL_198 & _EVAL_246;
  assign _EVAL_67 = _EVAL_270 | _EVAL_306;
  assign _EVAL_408 = _EVAL_367 ? _EVAL_177 : _EVAL_396;
  assign _EVAL_319 = {_EVAL_273, 2'h0};
  assign _EVAL_426 = _EVAL_100[3:1];
  assign _EVAL_356 = ~_EVAL_162;
  assign _EVAL_400 = _EVAL_287[1:0];
  assign _EVAL_465 = _EVAL_72 & _EVAL_454;
  assign _EVAL_428 = _EVAL_320 | _EVAL_509;
  assign _EVAL_297 = _EVAL_388 & _EVAL_107;
  assign _EVAL_330 = _EVAL_340 | _EVAL_406;
  assign _EVAL_504 = _EVAL_99[3:1];
  assign _EVAL_305 = _EVAL_149 | _EVAL_247;
  assign _EVAL_415 = _EVAL_312 ? _EVAL_29 : 4'h0;
  assign _EVAL_433 = _EVAL_461 & _EVAL_462;
  assign _EVAL_418 = _EVAL_435 | _EVAL_386;
  assign _EVAL_93 = _EVAL_172 | _EVAL_255;
  assign _EVAL_230 = {_EVAL_162, 2'h0};
  assign _EVAL_197 = _EVAL_112 & _EVAL_34;
  assign _EVAL_337 = _EVAL_313[3:1];
  assign _EVAL_159 = {_EVAL_453,_EVAL_275};
  assign _EVAL_341 = {{1'd0}, _EVAL_504};
  assign _EVAL_369 = {{1'd0}, _EVAL_421};
  assign _EVAL_425 = _EVAL_502 & _EVAL_487;
  assign _EVAL_165 = {1'b0,$signed(_EVAL_16)};
  assign _EVAL_310 = _EVAL_249 & _EVAL_1;
  assign _EVAL_438 = 23'hff << _EVAL_29;
  assign _EVAL_492 = _EVAL_365 & _EVAL_453;
  assign _EVAL_260 = _EVAL_52[4];
  assign _EVAL_120 = _EVAL_159 & _EVAL_356;
  assign _EVAL_224 = _EVAL_193 ? _EVAL_80 : 4'h0;
  assign _EVAL_117 = $signed(_EVAL_343) & 33'sh40000000;
  assign _EVAL_372 = 23'hff << _EVAL_70;
  assign _EVAL_509 = _EVAL_140 & _EVAL_202;
  assign _EVAL_199 = _EVAL_189 & _EVAL_159;
  assign _EVAL_166 = _EVAL_309;
  assign _EVAL_90 = _EVAL_466 | _EVAL_460;
  assign _EVAL_157 = _EVAL_485 & _EVAL_87;
  assign _EVAL_451 = {{1'd0}, _EVAL_20};
  assign _EVAL_489 = _EVAL_61 & _EVAL_510;
  assign _EVAL_441 = _EVAL_191[5:0];
  assign _EVAL_179 = _EVAL_203 & _EVAL_69;
  assign _EVAL_476 = {_EVAL_352, 1'h0};
  assign _EVAL_380 = _EVAL_485 & _EVAL_48;
  assign _EVAL_194 = _EVAL_199 | _EVAL_400;
  assign _EVAL_312 = _EVAL_482 ? _EVAL_384 : _EVAL_140;
  assign _EVAL_148 = _EVAL_284 ? _EVAL_206 : _EVAL_198;
  assign _EVAL_66 = _EVAL_141 | _EVAL_383;
  assign _EVAL_85 = _EVAL_326[3:0];
  assign _EVAL_325 = _EVAL_109 & _EVAL_251;
  assign _EVAL_4 = _EVAL_331 | _EVAL_444;
  assign _EVAL_306 = _EVAL_249 & _EVAL_32;
  assign _EVAL_290 = _EVAL_259 & _EVAL_484;
  assign _EVAL_167 = ~_EVAL_236;
  assign _EVAL_423 = $signed(_EVAL_450) & 33'sh40000000;
  assign _EVAL_467 = {{1'd0}, _EVAL_6};
  assign _EVAL_453 = _EVAL_75 & _EVAL_381;
  assign _EVAL_201 = _EVAL_78[0];
  assign _EVAL_214 = _EVAL_116[5:0];
  assign _EVAL_63 = _EVAL_358 | _EVAL_310;
  assign _EVAL_79 = _EVAL_221 | _EVAL_405;
  assign _EVAL_444 = _EVAL_249 ? _EVAL_91 : 4'h0;
  assign _EVAL_401 = _EVAL_189[0];
  assign _EVAL_384 = _EVAL_449 & _EVAL_202;
  assign _EVAL_99 = {_EVAL_120,_EVAL_453,_EVAL_275};
  assign _EVAL_316 = _EVAL_112 ? _EVAL_451 : 4'h0;
  assign _EVAL_374 = _EVAL_485 ? _EVAL_31 : 2'h0;
  assign _EVAL_379 = _EVAL_148 ? _EVAL_53 : 32'h0;
  assign _EVAL_398 = _EVAL_367 ? _EVAL_401 : _EVAL_396;
  assign _EVAL_276 = _EVAL_131[5:0];
  assign _EVAL_38 = _EVAL_459 | _EVAL_269;
  assign _EVAL_445 = _EVAL_416 & _EVAL_453;
  assign _EVAL_233 = _EVAL_203 & _EVAL_36;
  assign _EVAL_409 = {_EVAL_246,_EVAL_394};
  assign _EVAL_456 = _EVAL_423;
  assign _EVAL_392 = _EVAL_510 & _EVAL_115;
  assign _EVAL_323 = _EVAL_399[7:0];
  assign _EVAL_365 = _EVAL_189[1];
  assign _EVAL_481 = _EVAL_476[1:0];
  assign _EVAL_141 = _EVAL_203 ? _EVAL_9 : 3'h0;
  assign _EVAL_171 = _EVAL_105 | _EVAL_231;
  assign _EVAL_24 = _EVAL_366 | _EVAL_178;
  assign _EVAL_383 = _EVAL_312 ? _EVAL_11 : 3'h0;
  assign _EVAL_493 = _EVAL_148 ? _EVAL_56 : 3'h0;
  assign _EVAL_282 = _EVAL_112 ? _EVAL_21 : 2'h0;
  assign _EVAL_256 = _EVAL_329[5:0];
  assign _EVAL_262 = {{5'd0}, _EVAL_208};
  assign _EVAL_19 = _EVAL_181 | _EVAL_336;
  assign _EVAL_7 = _EVAL_367 ? _EVAL_114 : _EVAL_227;
  assign _EVAL_172 = _EVAL_408 & _EVAL_36;
  assign _EVAL_97 = _EVAL_50[4:1];
  assign _EVAL_402 = _EVAL_485 ? _EVAL_96 : 32'h0;
  assign _EVAL_126 = {{1'd0}, _EVAL_150};
  assign _EVAL_220 = _EVAL_395 == 6'h0;
  assign _EVAL_237 = {{5'd0}, _EVAL_397};
  assign _EVAL_147 = _EVAL_148 ? _EVAL_50 : 5'h0;
  assign _EVAL_450 = {1'b0,$signed(_EVAL_18)};
  assign _EVAL_219 = _EVAL_482 ? _EVAL_180 : _EVAL_479;
  assign _EVAL_482 = _EVAL_163 == 6'h0;
  assign _EVAL_485 = _EVAL_284 ? _EVAL_506 : _EVAL_299;
  assign _EVAL_403 = _EVAL_244 == 4'h8;
  assign _EVAL_258 = _EVAL_193 & _EVAL_57;
  assign _EVAL_264 = _EVAL_465 | _EVAL_484;
  assign _EVAL_370 = _EVAL_249 & _EVAL_30;
  assign _EVAL_397 = _EVAL_68 & _EVAL_455;
  assign _EVAL_281 = _EVAL_505 ? _EVAL_333 : 6'h0;
  assign _EVAL_127 = _EVAL_372[7:0];
  assign _EVAL_183 = _EVAL_112 ? _EVAL_53 : 32'h0;
  assign _EVAL_192 = _EVAL_412 & _EVAL_124;
  assign _EVAL_252 = ~_EVAL_192;
  assign _EVAL_502 = _EVAL_220 & _EVAL_39;
  assign _EVAL_406 = _EVAL_348 & _EVAL_484;
  assign _EVAL_83 = _EVAL_380 | _EVAL_123;
  assign _EVAL_150 = _EVAL_151[3:1];
  assign _EVAL_288 = {{4'd0}, _EVAL_89};
  assign _EVAL_187 = _EVAL_335 & _EVAL_109;
  assign _EVAL_211 = _EVAL_408 & _EVAL_74;
  assign _EVAL_463 = _EVAL_290 ? _EVAL_200 : 4'h0;
  assign _EVAL_200 = _EVAL_499 ? _EVAL_501 : 4'h0;
  assign _EVAL_130 = _EVAL_64 & _EVAL_156;
  assign _EVAL_15 = _EVAL_142 | _EVAL_265;
  assign _EVAL_391 = _EVAL_177 ? _EVAL_427 : 6'h0;
  assign _EVAL_246 = _EVAL_27 & _EVAL_311;
  assign _EVAL_217 = _EVAL_68 & _EVAL_248;
  assign _EVAL_180 = _EVAL_335[0];
  assign _EVAL_421 = _EVAL_254[3:1];
  assign _EVAL_385 = _EVAL_39 & _EVAL_334;
  assign _EVAL_478 = _EVAL_369 | _EVAL_230;
  assign _EVAL_457 = _EVAL_249 ? _EVAL_94 : 32'h0;
  assign _EVAL_470 = _EVAL_292 & _EVAL_158;
  assign _EVAL_59 = _EVAL_284 ? _EVAL_232 : _EVAL_429;
  assign _EVAL_189 = ~_EVAL_491;
  assign _EVAL_177 = _EVAL_401 & _EVAL_275;
  assign _EVAL_366 = _EVAL_485 & _EVAL_57;
  assign _EVAL_318 = _EVAL_478[3:2];
  assign _EVAL_128 = _EVAL_312 & _EVAL_1;
  assign _EVAL_500 = |_EVAL_109;
  assign _EVAL_284 = _EVAL_321 == 6'h0;
  assign _EVAL_114 = _EVAL_275 | _EVAL_453;
  assign _EVAL_268 = _EVAL_381 & _EVAL_217;
  assign _EVAL_329 = _EVAL_163 - _EVAL_262;
  assign _EVAL_81 = _EVAL_472 | _EVAL_164;
  assign _EVAL_119 = _EVAL_249 ? _EVAL_11 : 3'h0;
  assign _EVAL_145 = _EVAL_18 ^ 32'h40000000;
  assign _EVAL_123 = _EVAL_148 & _EVAL_34;
  assign _EVAL_190 = _EVAL_408 & _EVAL_77;
  assign _EVAL_422 = _EVAL_203 & _EVAL_14;
  assign _EVAL_354 = _EVAL_299 & _EVAL_394;
  assign _EVAL_121 = _EVAL_477[1];
  assign _EVAL_113 = _EVAL_68 & _EVAL_398;
  assign _EVAL_296 = _EVAL_148 ? _EVAL_451 : 4'h0;
  assign _EVAL_35 = _EVAL_144 | _EVAL_143;
  assign _EVAL_178 = _EVAL_148 & _EVAL_42;
  assign _EVAL_100 = {_EVAL_346,_EVAL_246,_EVAL_394};
  assign _EVAL_188 = _EVAL_408 ? _EVAL_186 : 5'h0;
  assign _EVAL_483 = _EVAL_312 & _EVAL_43;
  assign _EVAL_161 = _EVAL_220 ? _EVAL_264 : _EVAL_330;
  assign _EVAL_336 = _EVAL_312 ? _EVAL_54 : 3'h0;
  assign _EVAL_173 = _EVAL_193 ? _EVAL_52 : 5'h0;
  assign _EVAL_55 = _EVAL_482 ? _EVAL_382 : _EVAL_428;
  assign _EVAL_339 = _EVAL_222[3:1];
  assign _EVAL_437 = {{1'd0}, _EVAL_339};
  assign _EVAL_309 = $signed(_EVAL_234) & 33'sh40000000;
  assign _EVAL_460 = _EVAL_454 & _EVAL_357;
  assign _EVAL_73 = _EVAL_498 | _EVAL_282;
  assign _EVAL_440 = _EVAL_367 & _EVAL_68;
  assign _EVAL_326 = _EVAL_173 | _EVAL_436;
  assign _EVAL_229 = {{1'd0}, _EVAL_337};
  assign _EVAL_283 = {{5'd0}, _EVAL_130};
  assign _EVAL_95 = _EVAL_447 | _EVAL_169;
  assign _EVAL_382 = _EVAL_489 | _EVAL_202;
  assign _EVAL_203 = _EVAL_482 ? _EVAL_212 : _EVAL_479;
  assign _EVAL_110 = _EVAL_174 & _EVAL_385;
  assign _EVAL_251 = ~_EVAL_338;
  assign _EVAL_37 = _EVAL_392 | _EVAL_301;
  assign _EVAL_469 = _EVAL_195 & _EVAL_500;
  assign _EVAL_480 = _EVAL_284 ? _EVAL_363 : _EVAL_299;
  assign _EVAL_381 = $signed(_EVAL_166) == 33'sh0;
  assign _EVAL_473 = _EVAL_359[5:0];
  assign _EVAL_195 = _EVAL_482 & _EVAL_26;
  assign _EVAL_13 = _EVAL_424 | _EVAL_368;
  assign _EVAL_111 = ~_EVAL_127;
  assign _EVAL_170 = {{2'd0}, _EVAL_373};
  assign _EVAL_331 = _EVAL_408 ? _EVAL_5 : 4'h0;
  assign _EVAL_499 = _EVAL_56[0];
  assign _EVAL_477 = ~_EVAL_300;
  assign _EVAL_196 = _EVAL_229 | _EVAL_263;
  assign _EVAL_174 = ~_EVAL_371;
  assign _EVAL_136 = _EVAL_312 ? _EVAL_18 : 32'h0;
  assign _EVAL_115 = _EVAL_26 & _EVAL_219;
  assign _EVAL_164 = _EVAL_249 ? _EVAL_54 : 3'h0;
  assign _EVAL_405 = _EVAL_312 ? _EVAL_94 : 32'h0;
  assign _EVAL_448 = _EVAL_203 ? _EVAL_70 : 4'h0;
  assign _EVAL_107 = _EVAL_26 & _EVAL_314;
  assign _EVAL_491 = _EVAL_318 & _EVAL_508;
  assign _EVAL_152 = _EVAL_139[3:1];
  assign _EVAL_202 = _EVAL_75 & _EVAL_388;
  assign _EVAL_439 = _EVAL_486;
  assign _EVAL_313 = _EVAL_243 | _EVAL_242;
  assign _EVAL_505 = ~_EVAL_291;
  assign _EVAL_452 = _EVAL_391 | _EVAL_213;
  assign _EVAL_271 = _EVAL_252 & _EVAL_474;
  assign _EVAL_60 = _EVAL_488 | _EVAL_296;
  assign _EVAL_373 = _EVAL_206 ? _EVAL_200 : 4'h0;
  assign _EVAL_44 = _EVAL_190 | _EVAL_351;
  assign _EVAL_455 = _EVAL_367 ? _EVAL_114 : _EVAL_227;
  assign _EVAL_386 = _EVAL_384 ? _EVAL_281 : 6'h0;
  assign _EVAL_255 = _EVAL_249 & _EVAL_43;
  assign _EVAL_346 = _EVAL_409 & _EVAL_377;
  assign _EVAL_65 = _EVAL_297 | _EVAL_268;
  assign _EVAL_186 = _EVAL_288 | 5'h10;
  assign _EVAL_215 = _EVAL_482 ? _EVAL_382 : _EVAL_428;
  assign _EVAL_357 = _EVAL_39 & _EVAL_103;
  assign _EVAL_291 = _EVAL_11[2];
  assign _EVAL_412 = _EVAL_496[3:2];
  assign _EVAL_151 = _EVAL_100 | _EVAL_168;
  assign _EVAL_62 = _EVAL_211 | _EVAL_370;
  assign _EVAL_221 = _EVAL_203 ? _EVAL_82 : 32'h0;
  assign _EVAL_242 = {{1'd0}, _EVAL_407};
  assign _EVAL_311 = _EVAL_97 == 4'h8;
  assign _EVAL_345 = ~_EVAL_273;
  assign _EVAL_191 = _EVAL_321 - _EVAL_283;
  assign _EVAL_459 = _EVAL_203 ? _EVAL_186 : 5'h0;
  assign _EVAL_263 = {_EVAL_338, 2'h0};
  assign _EVAL_76 = _EVAL_224 | _EVAL_316;
  assign _EVAL_322 = _EVAL_271 | _EVAL_146;
  assign _EVAL_267 = _EVAL_332 ? _EVAL_349 : 6'h0;
  assign _EVAL_320 = _EVAL_479 & _EVAL_489;
  assign _EVAL_266 = _EVAL_16 ^ 32'h40000000;
  assign _EVAL_364 = {_EVAL_271, 1'h0};
  always @(posedge _EVAL_10) begin
    if (_EVAL) begin
      _EVAL_140 <= 1'h0;
    end else if (_EVAL_482) begin
      _EVAL_140 <= _EVAL_384;
    end
    if (_EVAL) begin
      _EVAL_162 <= 2'h3;
    end else if (_EVAL_417) begin
      _EVAL_162 <= _EVAL_194;
    end
    if (_EVAL) begin
      _EVAL_163 <= 6'h0;
    end else if (_EVAL_195) begin
      _EVAL_163 <= _EVAL_418;
    end else begin
      _EVAL_163 <= _EVAL_256;
    end
    if (_EVAL) begin
      _EVAL_198 <= 1'h0;
    end else if (_EVAL_284) begin
      _EVAL_198 <= _EVAL_206;
    end
    if (_EVAL) begin
      _EVAL_240 <= 2'h3;
    end else if (_EVAL_470) begin
      _EVAL_240 <= _EVAL_389;
    end
    if (_EVAL) begin
      _EVAL_273 <= 2'h3;
    end else if (_EVAL_425) begin
      _EVAL_273 <= _EVAL_322;
    end
    if (_EVAL) begin
      _EVAL_298 <= 6'h0;
    end else if (_EVAL_440) begin
      _EVAL_298 <= _EVAL_452;
    end else begin
      _EVAL_298 <= _EVAL_276;
    end
    if (_EVAL) begin
      _EVAL_299 <= 1'h0;
    end else if (_EVAL_284) begin
      _EVAL_299 <= _EVAL_506;
    end
    if (_EVAL) begin
      _EVAL_321 <= 6'h0;
    end else if (_EVAL_292) begin
      _EVAL_321 <= _EVAL_376;
    end else begin
      _EVAL_321 <= _EVAL_441;
    end
    if (_EVAL) begin
      _EVAL_338 <= 2'h3;
    end else if (_EVAL_469) begin
      _EVAL_338 <= _EVAL_277;
    end
    if (_EVAL) begin
      _EVAL_348 <= 1'h0;
    end else if (_EVAL_220) begin
      _EVAL_348 <= _EVAL_290;
    end
    if (_EVAL) begin
      _EVAL_395 <= 6'h0;
    end else if (_EVAL_502) begin
      _EVAL_395 <= _EVAL_216;
    end else begin
      _EVAL_395 <= _EVAL_214;
    end
    if (_EVAL) begin
      _EVAL_396 <= 1'h0;
    end else if (_EVAL_367) begin
      _EVAL_396 <= _EVAL_177;
    end
    if (_EVAL) begin
      _EVAL_416 <= 1'h0;
    end else if (_EVAL_367) begin
      _EVAL_416 <= _EVAL_492;
    end
    if (_EVAL) begin
      _EVAL_475 <= 1'h0;
    end else if (_EVAL_220) begin
      _EVAL_475 <= _EVAL_332;
    end
    if (_EVAL) begin
      _EVAL_479 <= 1'h0;
    end else if (_EVAL_482) begin
      _EVAL_479 <= _EVAL_212;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_140 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_162 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_163 = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_198 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_240 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_273 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_298 = _RAND_6[5:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_299 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_321 = _RAND_8[5:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_338 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_348 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_395 = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_396 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_416 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_475 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_479 = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
