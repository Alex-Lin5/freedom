//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_124(
  output [29:0] _EVAL,
  output        _EVAL_0,
  output [1:0]  _EVAL_1,
  output [29:0] _EVAL_2,
  input  [31:0] _EVAL_3,
  output        _EVAL_4,
  output [29:0] _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  output [31:0] _EVAL_8,
  output        _EVAL_9,
  output        _EVAL_10,
  input  [1:0]  _EVAL_11,
  input         _EVAL_12,
  output        _EVAL_13,
  output        _EVAL_14,
  output        _EVAL_15,
  output        _EVAL_16,
  output        _EVAL_17,
  output        _EVAL_18,
  input  [29:0] _EVAL_19,
  output [1:0]  _EVAL_20,
  input         _EVAL_21,
  output        _EVAL_22,
  output        _EVAL_23,
  output        _EVAL_24,
  output        _EVAL_25,
  input         _EVAL_26,
  output        _EVAL_27,
  output        _EVAL_28,
  input         _EVAL_29,
  output        _EVAL_30,
  output        _EVAL_31,
  output        _EVAL_32,
  output        _EVAL_33,
  input  [1:0]  _EVAL_34,
  input         _EVAL_35,
  output        _EVAL_36,
  output        _EVAL_37,
  output        _EVAL_38,
  output [1:0]  _EVAL_39,
  output [29:0] _EVAL_40,
  input  [31:0] _EVAL_41,
  output        _EVAL_42,
  input         _EVAL_43,
  output [31:0] _EVAL_44,
  input         _EVAL_45,
  input         _EVAL_46,
  input         _EVAL_47,
  input  [29:0] _EVAL_48,
  input  [1:0]  _EVAL_49,
  input  [29:0] _EVAL_50,
  output        _EVAL_51,
  output        _EVAL_52,
  output        _EVAL_53,
  input  [1:0]  _EVAL_54,
  input         _EVAL_55,
  input         _EVAL_56,
  output        _EVAL_57,
  output        _EVAL_58,
  output        _EVAL_59,
  input         _EVAL_60,
  input  [1:0]  _EVAL_61,
  output        _EVAL_62,
  output [31:0] _EVAL_63,
  output [31:0] _EVAL_64,
  input  [29:0] _EVAL_65,
  input         _EVAL_66,
  input         _EVAL_67,
  output        _EVAL_68,
  output [29:0] _EVAL_69,
  input         _EVAL_70,
  input  [31:0] _EVAL_71,
  input         _EVAL_72,
  output        _EVAL_73,
  output [1:0]  _EVAL_74,
  output [29:0] _EVAL_75,
  output        _EVAL_76,
  output [29:0] _EVAL_77,
  output [31:0] _EVAL_78,
  output        _EVAL_79,
  output        _EVAL_80,
  output [1:0]  _EVAL_81,
  input  [29:0] _EVAL_82,
  output        _EVAL_83,
  output        _EVAL_84,
  input         _EVAL_85,
  output        _EVAL_86,
  input  [31:0] _EVAL_87,
  output        _EVAL_88,
  input  [31:0] _EVAL_89,
  input  [31:0] _EVAL_90,
  output        _EVAL_91,
  input  [1:0]  _EVAL_92,
  output [1:0]  _EVAL_93,
  input  [31:0] _EVAL_94,
  output [1:0]  _EVAL_95,
  output        _EVAL_96,
  output [29:0] _EVAL_97,
  output        _EVAL_98,
  output        _EVAL_99,
  input  [1:0]  _EVAL_100,
  input  [29:0] _EVAL_101,
  input         _EVAL_102,
  output [31:0] _EVAL_103,
  input         _EVAL_104,
  output [1:0]  _EVAL_105,
  output [29:0] _EVAL_106,
  input         _EVAL_107,
  output [1:0]  _EVAL_108,
  input         _EVAL_109,
  output [1:0]  _EVAL_110,
  output [31:0] _EVAL_111,
  output [1:0]  _EVAL_112,
  output [31:0] _EVAL_113,
  input         _EVAL_114,
  output [1:0]  _EVAL_115,
  output        _EVAL_116,
  output        _EVAL_117,
  output [31:0] _EVAL_118,
  input         _EVAL_119,
  input  [31:0] _EVAL_120,
  output [29:0] _EVAL_121,
  input  [1:0]  _EVAL_122,
  output        _EVAL_123,
  output        _EVAL_124,
  output [29:0] _EVAL_125,
  output [31:0] _EVAL_126,
  output        _EVAL_127,
  output        _EVAL_128,
  input  [29:0] _EVAL_129,
  output        _EVAL_130,
  input         _EVAL_131,
  output [1:0]  _EVAL_132,
  output        _EVAL_133,
  output [29:0] _EVAL_134,
  output        _EVAL_135,
  output        _EVAL_136,
  output [29:0] _EVAL_137,
  output [29:0] _EVAL_138,
  output [1:0]  _EVAL_139,
  input  [29:0] _EVAL_140,
  output        _EVAL_141,
  input         _EVAL_142,
  output [31:0] _EVAL_143,
  input         _EVAL_144,
  output        _EVAL_145,
  output        _EVAL_146,
  output [31:0] _EVAL_147,
  output        _EVAL_148,
  input  [1:0]  _EVAL_149,
  output        _EVAL_150,
  output [29:0] _EVAL_151,
  output        _EVAL_152,
  output [31:0] _EVAL_153,
  output        _EVAL_154,
  output        _EVAL_155,
  input  [31:0] _EVAL_156,
  output [29:0] _EVAL_157,
  output        _EVAL_158,
  output [31:0] _EVAL_159,
  output        _EVAL_160,
  output        _EVAL_161,
  output [1:0]  _EVAL_162,
  output [31:0] _EVAL_163,
  output        _EVAL_164,
  output [1:0]  _EVAL_165,
  input         _EVAL_166,
  input         _EVAL_167,
  output [31:0] _EVAL_168,
  input         _EVAL_169,
  input         _EVAL_170,
  output        _EVAL_171,
  output [1:0]  _EVAL_172,
  output        _EVAL_173,
  output [31:0] _EVAL_174,
  input         _EVAL_175,
  output        _EVAL_176,
  output [31:0] _EVAL_177,
  input  [1:0]  _EVAL_178,
  output        _EVAL_179,
  output        _EVAL_180,
  input         _EVAL_181,
  output [1:0]  _EVAL_182,
  output [31:0] _EVAL_183,
  input  [31:0] _EVAL_184,
  input         _EVAL_185,
  input         _EVAL_186,
  output        _EVAL_187
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire [31:0] _EVAL_197;
  wire  _EVAL_198;
  wire [31:0] _EVAL_199;
  wire [15:0] _EVAL_200;
  wire  _EVAL_201;
  wire [9:0] _EVAL_202;
  wire [31:0] _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire [25:0] _EVAL_207;
  wire  _EVAL_208;
  wire [9:0] _EVAL_209;
  wire  _EVAL_210;
  wire [31:0] _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire [19:0] _EVAL_218;
  wire [32:0] _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire [31:0] _EVAL_229;
  wire [31:0] _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire [31:0] _EVAL_233;
  wire [26:0] _EVAL_234;
  wire [19:0] _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire [31:0] _EVAL_240;
  wire  _EVAL_241;
  wire [31:0] _EVAL_243;
  wire [31:0] _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire [31:0] _EVAL_248;
  wire [31:0] _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire [31:0] _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire [19:0] _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire [31:0] _EVAL_264;
  wire  _EVAL_265;
  wire [31:0] _EVAL_266;
  wire  _EVAL_267;
  wire [14:0] _EVAL_268;
  wire [31:0] _EVAL_269;
  wire [31:0] _EVAL_270;
  wire [30:0] _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire [31:0] _EVAL_278;
  wire  _EVAL_279;
  wire  _EVAL_281;
  wire [28:0] _EVAL_282;
  wire  _EVAL_283;
  wire [28:0] _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire [30:0] _EVAL_287;
  wire  _EVAL_288;
  wire [2:0] state_barrier__EVAL;
  wire [2:0] state_barrier__EVAL_0;
  wire [31:0] _EVAL_289;
  wire  _EVAL_290;
  wire [25:0] _EVAL_291;
  wire [31:0] _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_294;
  wire  _EVAL_295;
  wire  _EVAL_296;
  wire  _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire [32:0] _EVAL_300;
  wire  _EVAL_302;
  wire  _EVAL_303;
  wire [31:0] _EVAL_304;
  wire  _EVAL_305;
  wire [25:0] _EVAL_306;
  wire  _EVAL_308;
  wire  _EVAL_309;
  wire  _EVAL_310;
  wire [14:0] _EVAL_311;
  wire  _EVAL_312;
  wire [30:0] _EVAL_313;
  wire  _EVAL_314;
  wire [2:0] _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_317;
  wire [31:0] _EVAL_318;
  wire  _EVAL_319;
  wire [31:0] _EVAL_320;
  wire  _EVAL_321;
  wire [31:0] _EVAL_322;
  wire [19:0] _EVAL_323;
  wire  _EVAL_324;
  wire  _EVAL_325;
  wire  _EVAL_326;
  wire [19:0] _EVAL_327;
  wire  _EVAL_328;
  wire [19:0] _EVAL_329;
  wire  _EVAL_330;
  wire  _EVAL_331;
  wire [31:0] _EVAL_332;
  wire  _EVAL_333;
  wire  _EVAL_335;
  wire  _EVAL_336;
  wire  _EVAL_337;
  wire  _EVAL_338;
  wire [31:0] _EVAL_339;
  wire  _EVAL_340;
  wire  _EVAL_341;
  wire  _EVAL_342;
  wire  _EVAL_343;
  wire  _EVAL_344;
  wire  _EVAL_345;
  wire [9:0] _EVAL_346;
  wire  _EVAL_347;
  wire  _EVAL_348;
  wire  _EVAL_349;
  wire  _EVAL_350;
  wire [31:0] _EVAL_351;
  wire  _EVAL_352;
  wire  _EVAL_353;
  wire  _EVAL_354;
  wire  _EVAL_355;
  wire [32:0] _EVAL_356;
  reg [2:0] _EVAL_357;
  wire  _EVAL_358;
  wire [19:0] _EVAL_359;
  wire  _EVAL_360;
  wire  _EVAL_361;
  wire  _EVAL_362;
  wire [31:0] _EVAL_363;
  wire  _EVAL_364;
  wire [14:0] _EVAL_365;
  wire  _EVAL_366;
  wire  _EVAL_367;
  wire [31:0] _EVAL_368;
  wire  _EVAL_369;
  wire [2:0] _EVAL_370;
  wire [31:0] _EVAL_371;
  wire [31:0] _EVAL_372;
  wire  _EVAL_373;
  wire  _EVAL_374;
  wire  arb__EVAL;
  wire  arb__EVAL_0;
  wire  arb__EVAL_1;
  wire  _EVAL_375;
  wire  _EVAL_376;
  wire [31:0] _EVAL_377;
  wire  _EVAL_378;
  wire [31:0] _EVAL_379;
  wire [19:0] _EVAL_380;
  wire [31:0] _EVAL_381;
  wire  _EVAL_382;
  wire  _EVAL_383;
  wire [31:0] _EVAL_384;
  wire  _EVAL_385;
  wire  _EVAL_386;
  wire  _EVAL_387;
  wire  _EVAL_388;
  wire  _EVAL_389;
  wire  _EVAL_390;
  wire [31:0] _EVAL_391;
  wire [31:0] _EVAL_392;
  wire [2:0] _EVAL_393;
  wire [31:0] _EVAL_394;
  wire  _EVAL_395;
  wire [15:0] _EVAL_396;
  wire  _EVAL_397;
  wire  _EVAL_398;
  wire  _EVAL_399;
  wire  _EVAL_400;
  wire  _EVAL_401;
  wire  _EVAL_402;
  wire [31:0] _EVAL_403;
  wire [31:0] _EVAL_404;
  wire  _EVAL_405;
  wire  _EVAL_406;
  wire  _EVAL_407;
  wire [1:0] _EVAL_408;
  wire  _EVAL_409;
  wire  _EVAL_410;
  wire [9:0] _EVAL_411;
  wire [2:0] _EVAL_412;
  wire  _EVAL_413;
  wire  _EVAL_414;
  wire  _EVAL_415;
  wire [9:0] _EVAL_416;
  wire  _EVAL_417;
  wire  _EVAL_418;
  wire [31:0] _EVAL_419;
  wire  _EVAL_420;
  wire [31:0] _EVAL_421;
  wire  _EVAL_422;
  wire [15:0] _EVAL_423;
  wire [9:0] _EVAL_424;
  wire  _EVAL_425;
  wire  _EVAL_426;
  wire  _EVAL_427;
  wire  _EVAL_428;
  wire [31:0] _EVAL_429;
  wire  _EVAL_430;
  wire [31:0] _EVAL_431;
  wire  _EVAL_432;
  wire  _EVAL_433;
  wire  _EVAL_434;
  wire [26:0] _EVAL_435;
  wire  _EVAL_436;
  wire  _EVAL_437;
  wire  _EVAL_438;
  wire  _EVAL_439;
  wire  _EVAL_440;
  wire [9:0] _EVAL_441;
  wire  _EVAL_442;
  wire  _EVAL_443;
  wire  _EVAL_444;
  reg  _EVAL_445;
  wire  _EVAL_446;
  wire  _EVAL_447;
  wire  _EVAL_448;
  wire  _EVAL_449;
  wire  _EVAL_450;
  wire  _EVAL_451;
  wire  _EVAL_452;
  wire [26:0] _EVAL_453;
  wire  _EVAL_454;
  wire  _EVAL_455;
  wire  _EVAL_456;
  wire [9:0] _EVAL_457;
  wire [28:0] _EVAL_458;
  wire  _EVAL_459;
  wire  _EVAL_460;
  wire  _EVAL_461;
  _EVAL_123 state_barrier (
    ._EVAL(state_barrier__EVAL),
    ._EVAL_0(state_barrier__EVAL_0)
  );
  _EVAL_122 arb (
    ._EVAL(arb__EVAL),
    ._EVAL_0(arb__EVAL_0),
    ._EVAL_1(arb__EVAL_1)
  );
  assign _EVAL_369 = _EVAL_218 != 20'h0;
  assign _EVAL_449 = ~_EVAL_314;
  assign _EVAL_52 = _EVAL_186;
  assign _EVAL_30 = _EVAL_131;
  assign _EVAL_288 = $signed(_EVAL_453) == 27'sh0;
  assign _EVAL_154 = _EVAL_170;
  assign _EVAL_397 = _EVAL_122[0];
  assign _EVAL_386 = _EVAL_54[1];
  assign _EVAL_146 = _EVAL_43;
  assign _EVAL_40 = _EVAL_48;
  assign _EVAL_314 = 32'h0 < _EVAL_320;
  assign _EVAL_359 = _EVAL_244[31:12];
  assign _EVAL_115 = _EVAL_149;
  assign _EVAL_141 = _EVAL_45;
  assign _EVAL_348 = _EVAL_100[0];
  assign _EVAL_309 = $signed(_EVAL_458) == 29'sh0;
  assign _EVAL_297 = _EVAL_444 | _EVAL_288;
  assign _EVAL_59 = _EVAL_7;
  assign _EVAL_298 = 32'h0 < _EVAL_199;
  assign _EVAL_160 = _EVAL_104;
  assign _EVAL_361 = _EVAL_61[1];
  assign _EVAL_203 = ~_EVAL_233;
  assign _EVAL_206 = _EVAL_445 ? _EVAL_428 : _EVAL_433;
  assign _EVAL_393 = _EVAL_213 ? 3'h1 : _EVAL_412;
  assign _EVAL_258 = _EVAL_355 | _EVAL_430;
  assign _EVAL_253 = 3'h2 == _EVAL_357;
  assign _EVAL_433 = _EVAL_156[21];
  assign _EVAL_124 = _EVAL_70;
  assign _EVAL_438 = _EVAL_344 | _EVAL_239;
  assign _EVAL_286 = _EVAL_90[21];
  assign _EVAL_374 = _EVAL_336 & _EVAL_345;
  assign _EVAL_159 = _EVAL_184;
  assign _EVAL_231 = _EVAL_308 & _EVAL_456;
  assign _EVAL_389 = _EVAL_34[0];
  assign _EVAL_10 = _EVAL_114;
  assign _EVAL_299 = _EVAL_388 ? _EVAL_275 : _EVAL_442;
  assign _EVAL_387 = _EVAL_87[21];
  assign _EVAL_332 = _EVAL_384 | 32'h3;
  assign _EVAL_222 = _EVAL_92[0];
  assign _EVAL_163 = _EVAL_71;
  assign _EVAL_337 = _EVAL_89[11];
  assign _EVAL_191 = ~_EVAL_276;
  assign _EVAL_367 = _EVAL_188 | _EVAL_333;
  assign _EVAL_226 = _EVAL_202 != 10'h0;
  assign _EVAL_304 = {_EVAL_48, 2'h0};
  assign _EVAL_382 = _EVAL_90[11];
  assign _EVAL_326 = _EVAL_386 ? _EVAL_195 : _EVAL_205;
  assign _EVAL_155 = _EVAL_56;
  assign _EVAL_74 = _EVAL_54;
  assign _EVAL_113 = _EVAL_3;
  assign _EVAL_443 = _EVAL_445 ? _EVAL_319 : _EVAL_387;
  assign _EVAL_164 = _EVAL_107;
  assign _EVAL_260 = $signed(_EVAL_291) == 26'sh0;
  assign _EVAL_145 = _EVAL_26;
  assign _EVAL_264 = _EVAL_270 | 32'h3;
  assign _EVAL_83 = _EVAL_167;
  assign _EVAL_428 = _EVAL_156[11];
  assign _EVAL_192 = _EVAL_206 | _EVAL_461;
  assign _EVAL_135 = _EVAL_26;
  assign _EVAL_190 = _EVAL_257 | _EVAL_321;
  assign _EVAL_416 = _EVAL_266[31:22];
  assign _EVAL_234 = {1'b0,$signed(26'h2000000)};
  assign _EVAL_383 = _EVAL_411 != 10'h0;
  assign _EVAL_362 = _EVAL_273 & _EVAL_210;
  assign _EVAL_350 = ~_EVAL_348;
  assign _EVAL_323 = _EVAL_254[31:12];
  assign _EVAL_424 = _EVAL_244[31:22];
  assign _EVAL_418 = _EVAL_438 | _EVAL_335;
  assign _EVAL_422 = ~_EVAL_389;
  assign _EVAL_408 = {1'b0,$signed(1'h0)};
  assign _EVAL_207 = $signed(_EVAL_306) & -26'sh4000;
  assign _EVAL_401 = 32'h0 < _EVAL_197;
  assign _EVAL_413 = _EVAL_347 ? _EVAL_272 : _EVAL_265;
  assign _EVAL_373 = _EVAL_191 | _EVAL_398;
  assign _EVAL_345 = _EVAL_417 ? _EVAL_252 : _EVAL_258;
  assign _EVAL_95 = _EVAL_122;
  assign _EVAL_454 = _EVAL_359 != 20'h0;
  assign _EVAL_205 = _EVAL_450 | _EVAL_316;
  assign _EVAL_293 = ~_EVAL_325;
  assign _EVAL_230 = _EVAL_243 & _EVAL_377;
  assign _EVAL_37 = _EVAL_119;
  assign _EVAL_243 = ~_EVAL_248;
  assign _EVAL_165 = _EVAL_49;
  assign _EVAL_42 = arb__EVAL_1;
  assign _EVAL_204 = _EVAL_261 != 20'h0;
  assign _EVAL_195 = _EVAL_414 | _EVAL_194;
  assign _EVAL_287 = {1'b0,$signed(30'h20000000)};
  assign _EVAL_32 = _EVAL_12;
  assign _EVAL_187 = _EVAL_66;
  assign _EVAL_434 = _EVAL_445 ? _EVAL_454 : _EVAL_328;
  assign _EVAL_431 = ~_EVAL_421;
  assign _EVAL_134 = _EVAL_140;
  assign _EVAL_125 = _EVAL_129;
  assign _EVAL_392 = _EVAL_431 | 32'h3;
  assign _EVAL_437 = _EVAL_448 ? _EVAL_256 : _EVAL_352;
  assign _EVAL_458 = _EVAL_284;
  assign _EVAL_429 = $signed(_EVAL_322) & -32'sh2000;
  assign _EVAL_436 = 32'h0 < _EVAL_372;
  assign _EVAL_402 = _EVAL_303 | _EVAL_409;
  assign _EVAL_148 = _EVAL_12;
  assign _EVAL_415 = 32'h0 < _EVAL_254;
  assign _EVAL_76 = _EVAL_85;
  assign _EVAL_232 = _EVAL_241 & _EVAL_349;
  assign _EVAL_399 = _EVAL_407 & _EVAL_420;
  assign _EVAL_197 = ~_EVAL_278;
  assign _EVAL_121 = _EVAL_129;
  assign _EVAL_199 = ~_EVAL_289;
  assign _EVAL_202 = _EVAL_320[31:22];
  assign _EVAL_39 = _EVAL_100;
  assign _EVAL_240 = _EVAL_254 & _EVAL_377;
  assign _EVAL_78 = _EVAL_89;
  assign _EVAL_320 = ~_EVAL_332;
  assign _EVAL_174 = _EVAL_41;
  assign _EVAL_270 = ~_EVAL_304;
  assign _EVAL_138 = _EVAL_82;
  assign _EVAL_266 = ~_EVAL_392;
  assign _EVAL_18 = _EVAL_60;
  assign _EVAL_171 = _EVAL_169;
  assign _EVAL_259 = _EVAL_460 | _EVAL_302;
  assign _EVAL_223 = _EVAL_297 | _EVAL_309;
  assign _EVAL_451 = 32'h0 < _EVAL_244;
  assign _EVAL_233 = {_EVAL_140, 2'h0};
  assign _EVAL_330 = _EVAL_178[1];
  assign _EVAL_417 = _EVAL_149[1];
  assign _EVAL_22 = _EVAL_186;
  assign _EVAL_17 = _EVAL_167;
  assign _EVAL_136 = _EVAL_85;
  assign _EVAL_404 = {_EVAL_129, 2'h0};
  assign _EVAL_457 = _EVAL_197[31:22];
  assign _EVAL_112 = _EVAL_11;
  assign _EVAL_360 = 32'h0 < _EVAL_363;
  assign _EVAL_453 = _EVAL_435;
  assign _EVAL_346 = _EVAL_243[31:22];
  assign _EVAL_244 = ~_EVAL_264;
  assign _EVAL_128 = _EVAL_175;
  assign _EVAL_372 = ~_EVAL_381;
  assign _EVAL_4 = _EVAL_144;
  assign _EVAL_255 = _EVAL_445 ? _EVAL_406 : _EVAL_447;
  assign _EVAL_425 = _EVAL_445 ? _EVAL_337 : _EVAL_459;
  assign _EVAL_105 = _EVAL_61;
  assign _EVAL_409 = $signed(_EVAL_268) == 15'sh0;
  assign _EVAL_363 = _EVAL_199 & _EVAL_377;
  assign _EVAL_364 = $signed(_EVAL_271) == 31'sh0;
  assign _EVAL_173 = _EVAL_142;
  assign _EVAL_365 = $signed(_EVAL_311) & -15'sh1000;
  assign _EVAL_209 = _EVAL_372[31:22];
  assign _EVAL_117 = _EVAL_60;
  assign _EVAL_168 = _EVAL_87;
  assign _EVAL_276 = _EVAL_178[0];
  assign _EVAL_249 = ~_EVAL_292;
  assign _EVAL_25 = _EVAL_70;
  assign _EVAL_318 = {_EVAL_65, 2'h0};
  assign _EVAL_254 = ~_EVAL_269;
  assign _EVAL_447 = _EVAL_184[21];
  assign _EVAL_398 = _EVAL_367 | _EVAL_426;
  assign _EVAL_84 = _EVAL_102;
  assign _EVAL_444 = _EVAL_402 | _EVAL_260;
  assign _EVAL_51 = arb__EVAL;
  assign _EVAL_306 = {1'b0,$signed(25'h1800000)};
  assign _EVAL_69 = _EVAL_19;
  assign _EVAL_375 = 32'h0 < _EVAL_379;
  assign _EVAL_282 = {1'b0,$signed(28'hc000000)};
  assign _EVAL_14 = _EVAL_109;
  assign _EVAL_290 = _EVAL_333 & _EVAL_360;
  assign _EVAL_257 = ~_EVAL_277;
  assign _EVAL_335 = $signed(_EVAL_300) == 33'sh0;
  assign _EVAL_261 = _EVAL_199[31:12];
  assign _EVAL_180 = _EVAL_109;
  assign _EVAL_24 = _EVAL_46;
  assign _EVAL_211 = _EVAL_244 & _EVAL_377;
  assign _EVAL_296 = ~_EVAL_222;
  assign _EVAL_151 = _EVAL_19;
  assign _EVAL_96 = _EVAL_55;
  assign _EVAL_133 = _EVAL_45;
  assign _EVAL_331 = _EVAL_149[0];
  assign _EVAL_241 = ~_EVAL_451;
  assign _EVAL_292 = {_EVAL_82, 2'h0};
  assign _EVAL_291 = _EVAL_207;
  assign _EVAL_278 = _EVAL_419 | 32'h3;
  assign _EVAL_172 = _EVAL_34;
  assign _EVAL_396 = $signed(_EVAL_423) & -16'sh5000;
  assign _EVAL_456 = _EVAL_361 ? _EVAL_263 : _EVAL_190;
  assign _EVAL_8 = _EVAL_94;
  assign _EVAL_99 = _EVAL_47;
  assign _EVAL_214 = _EVAL_231 & _EVAL_413;
  assign _EVAL_400 = _EVAL_310 ? _EVAL_366 : _EVAL_281;
  assign _EVAL_158 = _EVAL_181;
  assign _EVAL_31 = _EVAL_46;
  assign _EVAL_150 = _EVAL_21;
  assign _EVAL_176 = _EVAL_6;
  assign _EVAL_325 = 32'h0 < _EVAL_266;
  assign _EVAL_305 = _EVAL_3[11];
  assign _EVAL_137 = _EVAL_82;
  assign _EVAL_423 = {{14{_EVAL_408[1]}},_EVAL_408};
  assign _EVAL_5 = _EVAL_50;
  assign _EVAL_81 = _EVAL_61;
  assign _EVAL_118 = _EVAL_87;
  assign _EVAL_441 = _EVAL_254[31:22];
  assign _EVAL_126 = _EVAL_94;
  assign _EVAL_385 = _EVAL_445 ? _EVAL_238 : _EVAL_245;
  assign _EVAL_227 = _EVAL_327 != 20'h0;
  assign _EVAL_273 = ~_EVAL_250;
  assign _EVAL_201 = _EVAL_295 | _EVAL_445;
  assign _EVAL_442 = _EVAL_224 | _EVAL_198;
  assign _EVAL_455 = _EVAL_213 ? 1'h0 : _EVAL_440;
  assign _EVAL_358 = 3'h7 == _EVAL_357;
  assign _EVAL_229 = _EVAL_320 & _EVAL_377;
  assign _EVAL_440 = _EVAL_253 ? 1'h0 : _EVAL_225;
  assign _EVAL_339 = _EVAL_197 & _EVAL_377;
  assign _EVAL_295 = ~_EVAL_189;
  assign _EVAL_188 = 32'h0 < _EVAL_229;
  assign _EVAL_127 = _EVAL_6;
  assign _EVAL_221 = _EVAL_346 != 10'h0;
  assign _EVAL_333 = ~_EVAL_415;
  assign _EVAL_220 = _EVAL_262 & _EVAL_375;
  assign _EVAL_57 = _EVAL_67;
  assign _EVAL_88 = _EVAL_247 ? 1'h0 : _EVAL_455;
  assign _EVAL_430 = _EVAL_446 | _EVAL_232;
  assign _EVAL_391 = ~_EVAL_371;
  assign _EVAL_75 = _EVAL_48;
  assign _EVAL_317 = _EVAL_209 != 10'h0;
  assign _EVAL_403 = {_EVAL_19, 2'h0};
  assign _EVAL_80 = _EVAL_47;
  assign _EVAL_321 = _EVAL_216 | _EVAL_220;
  assign _EVAL_366 = _EVAL_255 | _EVAL_434;
  assign _EVAL_338 = _EVAL_94[21];
  assign _EVAL_189 = _EVAL_432 & _EVAL_353;
  assign _EVAL_53 = _EVAL_166;
  assign _EVAL_405 = _EVAL_445 ? _EVAL_274 : _EVAL_410;
  assign _EVAL_432 = _EVAL_445 ? _EVAL_418 : _EVAL_309;
  assign _EVAL_250 = 32'h0 < _EVAL_243;
  assign _EVAL_420 = 32'h0 < _EVAL_211;
  assign _EVAL_15 = _EVAL_56;
  assign _EVAL_91 = _EVAL_107;
  assign _EVAL_289 = _EVAL_351 | 32'h3;
  assign _EVAL_208 = _EVAL_330 ? _EVAL_192 : _EVAL_373;
  assign _EVAL_13 = _EVAL_170;
  assign _EVAL_108 = _EVAL_149;
  assign _EVAL_38 = _EVAL_7;
  assign _EVAL_62 = _EVAL_55;
  assign _EVAL_153 = _EVAL_120;
  assign _EVAL_351 = ~_EVAL_403;
  assign _EVAL_376 = _EVAL_445 ? _EVAL_382 : _EVAL_286;
  assign _EVAL_450 = ~_EVAL_452;
  assign _EVAL_212 = _EVAL_41[21];
  assign _EVAL_460 = _EVAL_375 | _EVAL_407;
  assign _EVAL_316 = _EVAL_324 | _EVAL_290;
  assign _EVAL_461 = _EVAL_445 ? _EVAL_294 : _EVAL_217;
  assign _EVAL_64 = _EVAL_3;
  assign state_barrier__EVAL_0 = _EVAL_247 ? _EVAL_357 : _EVAL_393;
  assign _EVAL_352 = _EVAL_422 | _EVAL_395;
  assign _EVAL_328 = _EVAL_424 != 10'h0;
  assign _EVAL_210 = 32'h0 < _EVAL_394;
  assign _EVAL_324 = _EVAL_267 | _EVAL_262;
  assign _EVAL_239 = $signed(_EVAL_368) == 32'sh0;
  assign _EVAL_427 = _EVAL_341 | _EVAL_399;
  assign _EVAL_459 = _EVAL_89[21];
  assign _EVAL_284 = $signed(_EVAL_282) & -29'sh400000;
  assign _EVAL_275 = _EVAL_390 | _EVAL_340;
  assign _EVAL_182 = _EVAL_178;
  assign _EVAL_193 = _EVAL_445 ? _EVAL_285 : _EVAL_338;
  assign _EVAL_200 = _EVAL_396;
  assign _EVAL_315 = _EVAL_342 ? 3'h5 : _EVAL_370;
  assign _EVAL_435 = $signed(_EVAL_234) & -27'sh10000;
  assign _EVAL_370 = _EVAL_358 ? 3'h0 : _EVAL_357;
  assign _EVAL_224 = ~_EVAL_397;
  assign _EVAL_421 = {_EVAL_50, 2'h0};
  assign _EVAL_281 = _EVAL_296 | _EVAL_427;
  assign _EVAL_380 = _EVAL_266[31:12];
  assign _EVAL_354 = _EVAL_445 ? _EVAL_369 : _EVAL_317;
  assign _EVAL_68 = _EVAL_185;
  assign _EVAL_407 = ~_EVAL_401;
  assign _EVAL_274 = _EVAL_329 != 20'h0;
  assign _EVAL_238 = _EVAL_380 != 20'h0;
  assign _EVAL_371 = {_EVAL_101, 2'h0};
  assign _EVAL_23 = _EVAL_166;
  assign _EVAL_198 = _EVAL_449 | _EVAL_188;
  assign _EVAL_277 = _EVAL_61[0];
  assign _EVAL_406 = _EVAL_184[11];
  assign _EVAL_179 = _EVAL_21;
  assign _EVAL_300 = _EVAL_219;
  assign _EVAL_439 = _EVAL_299 & _EVAL_208;
  assign _EVAL_343 = ~_EVAL_436;
  assign _EVAL_228 = _EVAL_445 < 1'h1;
  assign _EVAL_379 = _EVAL_266 & _EVAL_377;
  assign _EVAL_353 = _EVAL_374 & _EVAL_437;
  assign _EVAL_217 = _EVAL_441 != 10'h0;
  assign _EVAL_294 = _EVAL_323 != 20'h0;
  assign _EVAL_412 = _EVAL_253 ? 3'h4 : _EVAL_315;
  assign _EVAL_426 = _EVAL_449 & _EVAL_267;
  assign _EVAL_1 = _EVAL_178;
  assign _EVAL_28 = _EVAL_29;
  assign _EVAL_36 = 1'h0;
  assign _EVAL_247 = 3'h0 == _EVAL_357;
  assign _EVAL_9 = _EVAL_66;
  assign _EVAL_256 = _EVAL_425 | _EVAL_354;
  assign _EVAL_329 = _EVAL_197[31:12];
  assign _EVAL_73 = _EVAL_181;
  assign _EVAL_132 = _EVAL_92;
  assign _EVAL_123 = _EVAL_114;
  assign _EVAL_20 = _EVAL_34;
  assign _EVAL_103 = _EVAL_184;
  assign _EVAL_110 = _EVAL_92;
  assign _EVAL_310 = _EVAL_92[1];
  assign _EVAL_268 = _EVAL_365;
  assign _EVAL_384 = ~_EVAL_318;
  assign _EVAL_279 = _EVAL_41[11];
  assign _EVAL_216 = _EVAL_360 | _EVAL_293;
  assign _EVAL_63 = _EVAL_90;
  assign _EVAL_147 = _EVAL_71;
  assign _EVAL_452 = _EVAL_54[0];
  assign _EVAL_271 = _EVAL_313;
  assign _EVAL_143 = _EVAL_156;
  assign _EVAL_262 = ~_EVAL_298;
  assign _EVAL_340 = _EVAL_445 ? _EVAL_196 : _EVAL_226;
  assign _EVAL_394 = _EVAL_372 & _EVAL_377;
  assign _EVAL_215 = _EVAL_445 ? _EVAL_227 : _EVAL_221;
  assign _EVAL_448 = _EVAL_34[1];
  assign _EVAL_252 = _EVAL_443 | _EVAL_215;
  assign _EVAL_161 = _EVAL_102;
  assign _EVAL_355 = ~_EVAL_331;
  assign _EVAL_313 = $signed(_EVAL_287) & -31'sh2000;
  assign _EVAL_196 = _EVAL_237 != 20'h0;
  assign _EVAL_381 = _EVAL_249 | 32'h3;
  assign _EVAL_388 = _EVAL_122[1];
  assign _EVAL_327 = _EVAL_243[31:12];
  assign _EVAL_308 = _EVAL_439 & _EVAL_326;
  assign _EVAL_263 = _EVAL_376 | _EVAL_385;
  assign _EVAL_377 = _EVAL_445 ? 32'hfffff000 : 32'hffc00000;
  assign _EVAL_97 = _EVAL_101;
  assign _EVAL_116 = _EVAL_131;
  assign _EVAL_225 = _EVAL_342 & _EVAL_228;
  assign _EVAL_285 = _EVAL_94[11];
  assign _EVAL_213 = 3'h1 == _EVAL_357;
  assign _EVAL_130 = _EVAL_119;
  assign _EVAL_269 = _EVAL_391 | 32'h3;
  assign _EVAL_341 = _EVAL_283 | _EVAL_241;
  assign _EVAL_33 = _EVAL_67;
  assign _EVAL_390 = _EVAL_445 ? _EVAL_305 : _EVAL_246;
  assign _EVAL_419 = ~_EVAL_404;
  assign _EVAL_347 = _EVAL_100[1];
  assign _EVAL_368 = _EVAL_429;
  assign _EVAL_272 = _EVAL_193 | _EVAL_405;
  assign _EVAL_411 = _EVAL_199[31:22];
  assign _EVAL_2 = _EVAL_140;
  assign _EVAL_77 = _EVAL_50;
  assign _EVAL_349 = 32'h0 < _EVAL_230;
  assign _EVAL_219 = $signed(_EVAL_356) & -33'sh4000;
  assign _EVAL_218 = _EVAL_372[31:12];
  assign _EVAL_248 = _EVAL_203 | 32'h3;
  assign _EVAL_79 = _EVAL_169;
  assign _EVAL_312 = _EVAL_358 ? _EVAL_201 : _EVAL_445;
  assign _EVAL_27 = _EVAL_142;
  assign _EVAL_139 = _EVAL_100;
  assign _EVAL_183 = _EVAL_41;
  assign _EVAL_98 = _EVAL_175;
  assign _EVAL_245 = _EVAL_416 != 10'h0;
  assign _EVAL_111 = _EVAL_89;
  assign arb__EVAL_0 = _EVAL_357 == 3'h0;
  assign _EVAL_177 = _EVAL_90;
  assign _EVAL_378 = _EVAL_349 | _EVAL_343;
  assign _EVAL_356 = {1'b0,$signed(32'h80000000)};
  assign _EVAL_106 = _EVAL_65;
  assign _EVAL_342 = 3'h4 == _EVAL_357;
  assign _EVAL_322 = {1'b0,$signed(31'h40000000)};
  assign _EVAL_162 = _EVAL_122;
  assign _EVAL_152 = _EVAL_144;
  assign _EVAL_311 = {1'b0,$signed(14'h3000)};
  assign _EVAL_410 = _EVAL_457 != 10'h0;
  assign _EVAL_319 = _EVAL_87[11];
  assign _EVAL_237 = _EVAL_320[31:12];
  assign _EVAL_302 = _EVAL_293 & _EVAL_283;
  assign _EVAL_58 = 1'h0;
  assign _EVAL_0 = _EVAL_185;
  assign _EVAL_344 = _EVAL_223 | _EVAL_364;
  assign _EVAL_267 = 32'h0 < _EVAL_240;
  assign _EVAL_246 = _EVAL_3[21];
  assign _EVAL_446 = _EVAL_420 | _EVAL_273;
  assign _EVAL_86 = _EVAL_104;
  assign _EVAL_303 = $signed(_EVAL_200) == 16'sh0;
  assign _EVAL_395 = _EVAL_378 | _EVAL_362;
  assign _EVAL_194 = _EVAL_445 ? _EVAL_204 : _EVAL_383;
  assign _EVAL = _EVAL_101;
  assign _EVAL_93 = _EVAL_54;
  assign _EVAL_157 = _EVAL_65;
  assign _EVAL_44 = _EVAL_156;
  assign _EVAL_283 = 32'h0 < _EVAL_339;
  assign _EVAL_16 = _EVAL_29;
  assign _EVAL_265 = _EVAL_350 | _EVAL_259;
  assign _EVAL_414 = _EVAL_445 ? _EVAL_279 : _EVAL_212;
  assign _EVAL_336 = _EVAL_214 & _EVAL_400;
  always @(posedge _EVAL_72) begin
    if (_EVAL_35) begin
      _EVAL_357 <= 3'h0;
    end else begin
      _EVAL_357 <= state_barrier__EVAL;
    end
    if (_EVAL_247) begin
      _EVAL_445 <= 1'h0;
    end else if (!(_EVAL_213)) begin
      if (!(_EVAL_253)) begin
        if (!(_EVAL_342)) begin
          _EVAL_445 <= _EVAL_312;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_357 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_445 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
