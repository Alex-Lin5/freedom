//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_135_assert(
  input         _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [31:0] _EVAL_2,
  input         _EVAL_3,
  input  [2:0]  _EVAL_4,
  input  [3:0]  _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input  [1:0]  _EVAL_8,
  input         _EVAL_9,
  input  [3:0]  _EVAL_10,
  input  [2:0]  _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input  [3:0]  _EVAL_14,
  input  [3:0]  _EVAL_15,
  input  [3:0]  _EVAL_16,
  input  [2:0]  _EVAL_17,
  input         _EVAL_18
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire [5:0] _EVAL_23;
  reg [5:0] _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire [31:0] _EVAL_46;
  wire [2:0] _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire [32:0] _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire [5:0] _EVAL_60;
  wire  _EVAL_61;
  wire [32:0] _EVAL_62;
  wire [6:0] _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  reg [2:0] _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire [32:0] _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  reg  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire [3:0] _EVAL_86;
  wire  _EVAL_87;
  wire [31:0] _EVAL_88;
  wire [6:0] _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire [3:0] _EVAL_98;
  wire [31:0] _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  reg [1:0] _EVAL_107;
  wire  _EVAL_108;
  wire [31:0] _EVAL_109;
  wire [32:0] _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire [32:0] _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_117;
  wire [32:0] _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire [8:0] _EVAL_124;
  wire  _EVAL_125;
  reg  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire [32:0] _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire [5:0] _EVAL_135;
  wire [32:0] _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire [31:0] _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire [32:0] _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire [5:0] _EVAL_153;
  wire  _EVAL_154;
  wire [32:0] _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_158;
  wire [32:0] _EVAL_159;
  wire  _EVAL_160;
  wire [32:0] _EVAL_161;
  wire  _EVAL_162;
  reg [5:0] _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire [32:0] _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire [32:0] _EVAL_171;
  wire [32:0] _EVAL_172;
  reg [5:0] _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire [6:0] _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  reg [8:0] _EVAL_185;
  wire  _EVAL_186;
  reg [3:0] _EVAL_187;
  wire [15:0] _EVAL_188;
  reg [31:0] _EVAL_189;
  wire  _EVAL_190;
  wire [8:0] _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire [32:0] _EVAL_200;
  wire  _EVAL_201;
  reg [2:0] _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire [8:0] _EVAL_212;
  wire  _EVAL_213;
  wire [31:0] _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire [8:0] _EVAL_219;
  wire  _EVAL_220;
  wire [32:0] _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire [7:0] _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire [22:0] _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire [15:0] _EVAL_252;
  wire [7:0] _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire [8:0] _EVAL_256;
  wire  _EVAL_257;
  reg [3:0] _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire [32:0] _EVAL_263;
  wire [8:0] _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  reg [5:0] _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire [7:0] _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire [32:0] _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire [32:0] _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire [31:0] _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire [31:0] _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire  _EVAL_293;
  wire  _EVAL_294;
  wire [6:0] _EVAL_295;
  wire  _EVAL_296;
  wire [31:0] _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_307;
  wire [8:0] _EVAL_308;
  wire [32:0] _EVAL_309;
  wire  _EVAL_310;
  wire  _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire [15:0] _EVAL_317;
  wire  _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_320;
  wire  _EVAL_321;
  wire  _EVAL_322;
  wire  _EVAL_323;
  wire  _EVAL_324;
  wire [22:0] _EVAL_325;
  wire  _EVAL_326;
  wire [32:0] _EVAL_327;
  wire [1:0] _EVAL_328;
  wire  _EVAL_329;
  wire [32:0] _EVAL_330;
  wire [5:0] _EVAL_331;
  wire  _EVAL_332;
  wire  _EVAL_333;
  reg [31:0] _EVAL_334;
  reg [3:0] _EVAL_335;
  wire [1:0] _EVAL_336;
  wire  _EVAL_337;
  wire  _EVAL_338;
  wire  _EVAL_339;
  wire  _EVAL_340;
  wire  _EVAL_341;
  wire [32:0] _EVAL_342;
  wire  _EVAL_343;
  wire  _EVAL_344;
  wire [3:0] _EVAL_345;
  wire [32:0] _EVAL_346;
  wire  _EVAL_347;
  wire [7:0] _EVAL_348;
  wire  _EVAL_349;
  wire  _EVAL_350;
  wire [2:0] _EVAL_351;
  wire  _EVAL_352;
  wire [8:0] _EVAL_353;
  reg [3:0] _EVAL_354;
  wire  _EVAL_355;
  wire [5:0] _EVAL_356;
  wire  _EVAL_357;
  wire [3:0] _EVAL_358;
  wire [15:0] _EVAL_359;
  wire  _EVAL_360;
  wire  _EVAL_361;
  wire  _EVAL_362;
  wire [31:0] _EVAL_363;
  wire  _EVAL_364;
  wire  _EVAL_365;
  wire  _EVAL_366;
  wire  _EVAL_367;
  reg [2:0] _EVAL_369;
  wire  _EVAL_370;
  wire  _EVAL_371;
  wire  _EVAL_372;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_199 = _EVAL_256[0];
  assign _EVAL_82 = _EVAL_10 <= 4'h2;
  assign _EVAL_21 = _EVAL_0 == _EVAL_79;
  assign _EVAL_317 = 16'h1 << _EVAL_5;
  assign _EVAL_313 = ~_EVAL_7;
  assign _EVAL_245 = _EVAL & _EVAL_162;
  assign _EVAL_318 = _EVAL_4 <= 3'h2;
  assign _EVAL_211 = _EVAL_19 | _EVAL_6;
  assign _EVAL_137 = _EVAL_87 | _EVAL_76;
  assign _EVAL_268 = ~_EVAL_211;
  assign _EVAL_288 = _EVAL_310 | _EVAL_6;
  assign _EVAL_117 = _EVAL_56 | _EVAL_6;
  assign _EVAL_118 = $signed(_EVAL_74) & -33'sh10000;
  assign _EVAL_115 = ~_EVAL_42;
  assign _EVAL_155 = $signed(_EVAL_62) & -33'sh5000;
  assign _EVAL_316 = ~_EVAL_108;
  assign _EVAL_213 = ~_EVAL_324;
  assign _EVAL_349 = _EVAL_2 == _EVAL_334;
  assign _EVAL_357 = _EVAL & _EVAL_208;
  assign _EVAL_371 = _EVAL_32 | _EVAL_6;
  assign _EVAL_139 = _EVAL_2[1];
  assign _EVAL_90 = _EVAL & _EVAL_156;
  assign _EVAL_48 = _EVAL_10 >= 4'h2;
  assign _EVAL_293 = _EVAL_95 | _EVAL_360;
  assign _EVAL_224 = _EVAL_16 == 4'h8;
  assign _EVAL_161 = _EVAL_280;
  assign _EVAL_287 = _EVAL_2 ^ 32'h80000000;
  assign _EVAL_194 = ~_EVAL_301;
  assign _EVAL_244 = _EVAL_58 & _EVAL_272;
  assign _EVAL_331 = _EVAL_295[5:0];
  assign _EVAL_223 = _EVAL_11 == 3'h6;
  assign _EVAL_128 = _EVAL_239 | _EVAL_76;
  assign _EVAL_77 = ~_EVAL_100;
  assign _EVAL_159 = _EVAL_189 + 32'h1;
  assign _EVAL_370 = _EVAL_1 & _EVAL_26;
  assign _EVAL_36 = _EVAL_41 & _EVAL_367;
  assign _EVAL_97 = _EVAL_232 | _EVAL_127;
  assign _EVAL_55 = {1'b0,$signed(_EVAL_99)};
  assign _EVAL_310 = _EVAL_11 == _EVAL_67;
  assign _EVAL_109 = _EVAL_2 ^ 32'h1800000;
  assign _EVAL_135 = _EVAL_274[7:2];
  assign _EVAL_336 = 2'h1 << _EVAL_283;
  assign _EVAL_340 = _EVAL_151 | _EVAL_28;
  assign _EVAL_282 = _EVAL_12 == _EVAL_126;
  assign _EVAL_175 = $signed(_EVAL_110) == 33'sh0;
  assign _EVAL_214 = _EVAL_2 ^ 32'h40000000;
  assign _EVAL_70 = _EVAL_345 == 4'h0;
  assign _EVAL_272 = _EVAL_57 | _EVAL_229;
  assign _EVAL_89 = _EVAL_173 - 6'h1;
  assign _EVAL_34 = _EVAL_140 | _EVAL_115;
  assign _EVAL_28 = _EVAL_27 & _EVAL_73;
  assign _EVAL_176 = _EVAL & _EVAL_206;
  assign _EVAL_84 = _EVAL_87 | _EVAL_229;
  assign _EVAL_303 = _EVAL_254 & _EVAL_292;
  assign _EVAL_343 = _EVAL_5 == _EVAL_258;
  assign _EVAL_184 = _EVAL_237 | _EVAL_6;
  assign _EVAL_307 = _EVAL_17 == 3'h0;
  assign _EVAL_337 = _EVAL_273 & _EVAL_41;
  assign _EVAL_110 = _EVAL_277;
  assign _EVAL_69 = _EVAL_49 | _EVAL_6;
  assign _EVAL_253 = _EVAL_234[7:0];
  assign _EVAL_350 = _EVAL_65 | _EVAL_71;
  assign _EVAL_147 = _EVAL_27 & _EVAL_259;
  assign _EVAL_64 = _EVAL_203 & _EVAL_174;
  assign _EVAL_183 = ~_EVAL_117;
  assign _EVAL_242 = _EVAL_154 | _EVAL_6;
  assign _EVAL_237 = _EVAL_8 == 2'h0;
  assign _EVAL_302 = _EVAL_349 | _EVAL_6;
  assign _EVAL_20 = ~_EVAL_204;
  assign _EVAL_264 = _EVAL_212 >> _EVAL_16;
  assign _EVAL_345 = _EVAL_14 & _EVAL_86;
  assign _EVAL_276 = _EVAL_76 | _EVAL_296;
  assign _EVAL_198 = _EVAL_290 & _EVAL_193;
  assign _EVAL_154 = _EVAL_4 <= 3'h3;
  assign _EVAL_52 = _EVAL & _EVAL_179;
  assign _EVAL_142 = _EVAL_17 == _EVAL_202;
  assign _EVAL_326 = ~_EVAL_339;
  assign _EVAL_144 = _EVAL_232 & _EVAL_312;
  assign _EVAL_275 = ~_EVAL_362;
  assign _EVAL_367 = _EVAL_2[0];
  assign _EVAL_167 = ~_EVAL_338;
  assign _EVAL_342 = _EVAL_346;
  assign _EVAL_40 = _EVAL_250 & _EVAL_205;
  assign _EVAL_324 = _EVAL_320 | _EVAL_6;
  assign _EVAL_297 = {{24'd0}, _EVAL_274};
  assign _EVAL_95 = _EVAL_91 | _EVAL_143;
  assign _EVAL_339 = _EVAL_343 | _EVAL_6;
  assign _EVAL_295 = _EVAL_267 - 6'h1;
  assign _EVAL_218 = _EVAL_24 == 6'h0;
  assign _EVAL_257 = _EVAL_11 == 3'h2;
  assign _EVAL_314 = _EVAL_361 | _EVAL_6;
  assign _EVAL_323 = _EVAL_318 | _EVAL_6;
  assign _EVAL_205 = _EVAL_47 <= 3'h6;
  assign _EVAL_203 = _EVAL_82 & _EVAL_40;
  assign _EVAL_83 = _EVAL_5 == 4'h8;
  assign _EVAL_143 = plusarg_reader_out == 32'h0;
  assign _EVAL_243 = ~_EVAL_190;
  assign _EVAL_196 = ~_EVAL_6;
  assign _EVAL_322 = ~_EVAL_199;
  assign _EVAL_100 = _EVAL_85 | _EVAL_6;
  assign _EVAL_162 = _EVAL_17 == 3'h6;
  assign _EVAL_254 = _EVAL_10 <= 4'h8;
  assign _EVAL_148 = ~_EVAL_372;
  assign _EVAL_366 = _EVAL_240 & _EVAL_246;
  assign _EVAL_255 = _EVAL_16 == _EVAL_335;
  assign _EVAL_325 = 23'hff << _EVAL_10;
  assign _EVAL_222 = _EVAL_1 & _EVAL_43;
  assign _EVAL_75 = ~_EVAL_12;
  assign _EVAL_76 = $signed(_EVAL_136) == 33'sh0;
  assign _EVAL_263 = {1'b0,$signed(_EVAL_88)};
  assign _EVAL_149 = _EVAL_329 | _EVAL_6;
  assign _EVAL_215 = _EVAL_68 | _EVAL_6;
  assign _EVAL_141 = _EVAL_2 & _EVAL_297;
  assign _EVAL_362 = _EVAL_92 | _EVAL_6;
  assign _EVAL_32 = _EVAL_40 | _EVAL_83;
  assign _EVAL_269 = ~_EVAL_288;
  assign _EVAL_125 = _EVAL_366 | _EVAL_6;
  assign _EVAL_25 = _EVAL_238 | _EVAL_292;
  assign _EVAL_329 = _EVAL_8 == _EVAL_107;
  assign _EVAL_59 = _EVAL & _EVAL_210;
  assign _EVAL_300 = _EVAL_38 & _EVAL_83;
  assign _EVAL_216 = _EVAL_220 | _EVAL_6;
  assign _EVAL_281 = ~_EVAL_262;
  assign _EVAL_49 = _EVAL_15 >= 4'h2;
  assign _EVAL_119 = ~_EVAL_31;
  assign _EVAL_227 = ~_EVAL_253;
  assign _EVAL_85 = _EVAL_4 <= 3'h1;
  assign _EVAL_360 = _EVAL_189 < plusarg_reader_out;
  assign _EVAL_238 = $signed(_EVAL_171) == 33'sh0;
  assign _EVAL_23 = _EVAL_63[5:0];
  assign _EVAL_146 = _EVAL_180 | _EVAL_6;
  assign _EVAL_153 = _EVAL_227[7:2];
  assign _EVAL_46 = _EVAL_2 ^ 32'h3000;
  assign _EVAL_134 = ~_EVAL_69;
  assign _EVAL_166 = _EVAL_303 | _EVAL_260;
  assign _EVAL_312 = _EVAL_267 == 6'h0;
  assign _EVAL_178 = _EVAL_27 & _EVAL_36;
  assign _EVAL_182 = _EVAL_163 - 6'h1;
  assign _EVAL_217 = _EVAL_1 & _EVAL_247;
  assign _EVAL_43 = _EVAL_11 == 3'h4;
  assign _EVAL_127 = _EVAL_18 & _EVAL;
  assign _EVAL_256 = _EVAL_185 >> _EVAL_5;
  assign _EVAL_131 = _EVAL_17[0];
  assign _EVAL_192 = ~_EVAL_314;
  assign _EVAL_226 = _EVAL_70 | _EVAL_6;
  assign _EVAL_33 = ~_EVAL_225;
  assign _EVAL_71 = $signed(_EVAL_221) == 33'sh0;
  assign _EVAL_206 = ~_EVAL_61;
  assign _EVAL_61 = _EVAL_163 == 6'h0;
  assign _EVAL_114 = _EVAL_64 | _EVAL_6;
  assign _EVAL_86 = ~_EVAL_98;
  assign _EVAL_286 = _EVAL_166 | _EVAL_6;
  assign _EVAL_246 = _EVAL_82 & _EVAL_130;
  assign _EVAL_112 = ~_EVAL_114;
  assign _EVAL_315 = _EVAL_232 & _EVAL_311;
  assign _EVAL_306 = _EVAL_291 | _EVAL_224;
  assign _EVAL_44 = ~_EVAL_242;
  assign _EVAL_330 = _EVAL_145;
  assign _EVAL_101 = ~_EVAL_158;
  assign _EVAL_31 = _EVAL_313 | _EVAL_6;
  assign _EVAL_327 = {1'b0,$signed(_EVAL_109)};
  assign _EVAL_347 = ~_EVAL_146;
  assign _EVAL_130 = _EVAL_128 | _EVAL_229;
  assign _EVAL_53 = _EVAL_5[3];
  assign _EVAL_151 = _EVAL_48 | _EVAL_81;
  assign _EVAL_234 = 23'hff << _EVAL_15;
  assign _EVAL_240 = _EVAL_230 & _EVAL_40;
  assign _EVAL_352 = _EVAL_165 | _EVAL_6;
  assign _EVAL_27 = _EVAL_328[0];
  assign _EVAL_168 = {1'b0,$signed(_EVAL_214)};
  assign _EVAL_78 = ~_EVAL_54;
  assign _EVAL_120 = _EVAL_8 != 2'h2;
  assign _EVAL_358 = ~_EVAL_14;
  assign _EVAL_321 = ~_EVAL_105;
  assign _EVAL_58 = _EVAL_10 <= 4'h6;
  assign _EVAL_164 = _EVAL_4 == 3'h0;
  assign _EVAL_133 = ~_EVAL_285;
  assign _EVAL_271 = _EVAL_16[3];
  assign _EVAL_210 = _EVAL_17 == 3'h5;
  assign _EVAL_320 = _EVAL_15 == _EVAL_354;
  assign _EVAL_111 = _EVAL_25 | _EVAL_175;
  assign _EVAL_38 = 4'h6 == _EVAL_10;
  assign _EVAL_138 = _EVAL_58 & _EVAL_84;
  assign _EVAL_93 = _EVAL_14 == _EVAL_98;
  assign _EVAL_88 = _EVAL_2 ^ 32'h20000000;
  assign _EVAL_204 = _EVAL_322 | _EVAL_6;
  assign _EVAL_102 = $signed(_EVAL_330) == 33'sh0;
  assign _EVAL_291 = _EVAL_332 & _EVAL_169;
  assign _EVAL_304 = |_EVAL_185;
  assign _EVAL_177 = ~_EVAL_311;
  assign _EVAL_262 = _EVAL_51 | _EVAL_6;
  assign _EVAL_348 = _EVAL_325[7:0];
  assign _EVAL_171 = _EVAL_155;
  assign _EVAL_37 = _EVAL_48 | _EVAL_337;
  assign _EVAL_132 = _EVAL_1 & _EVAL_177;
  assign _EVAL_252 = 16'h1 << _EVAL_16;
  assign _EVAL_250 = ~_EVAL_53;
  assign _EVAL_294 = ~_EVAL_123;
  assign _EVAL_284 = _EVAL_159[31:0];
  assign _EVAL_122 = ~_EVAL_149;
  assign _EVAL_174 = _EVAL_303 | _EVAL_244;
  assign _EVAL_188 = _EVAL_198 ? _EVAL_252 : 16'h0;
  assign _EVAL_29 = ~_EVAL_216;
  assign _EVAL_190 = _EVAL_34 | _EVAL_6;
  assign _EVAL_129 = {1'b0,$signed(_EVAL_287)};
  assign _EVAL_172 = $signed(_EVAL_200) & -33'sh1000;
  assign _EVAL_179 = _EVAL_17 == 3'h1;
  assign _EVAL_19 = _EVAL_4 != 3'h0;
  assign _EVAL_56 = _EVAL_358 == 4'h0;
  assign _EVAL_42 = |_EVAL_124;
  assign _EVAL_87 = _EVAL_350 | _EVAL_102;
  assign _EVAL_124 = _EVAL_359[8:0];
  assign _EVAL_74 = {1'b0,$signed(_EVAL_363)};
  assign _EVAL_160 = _EVAL_93 | _EVAL_6;
  assign _EVAL_221 = _EVAL_118;
  assign _EVAL_105 = _EVAL_207 | _EVAL_6;
  assign _EVAL_104 = _EVAL_37 | _EVAL_178;
  assign _EVAL_47 = _EVAL_5[2:0];
  assign _EVAL_328 = _EVAL_336 | 2'h1;
  assign _EVAL_359 = _EVAL_144 ? _EVAL_317 : 16'h0;
  assign _EVAL_355 = ~_EVAL_186;
  assign _EVAL_170 = ~_EVAL_201;
  assign _EVAL_96 = _EVAL_41 & _EVAL_251;
  assign _EVAL_309 = _EVAL_172;
  assign _EVAL_277 = $signed(_EVAL_327) & -33'sh4000;
  assign _EVAL_152 = ~_EVAL_352;
  assign _EVAL_180 = _EVAL_141 == 32'h0;
  assign _EVAL_239 = _EVAL_197 | _EVAL_102;
  assign _EVAL_208 = _EVAL_17 == 3'h4;
  assign _EVAL_260 = _EVAL_58 & _EVAL_276;
  assign _EVAL_266 = _EVAL_1 & _EVAL_223;
  assign _EVAL_123 = _EVAL_48 | _EVAL_6;
  assign _EVAL_285 = _EVAL_261 | _EVAL_6;
  assign _EVAL_212 = _EVAL_124 | _EVAL_185;
  assign _EVAL_30 = _EVAL_164 | _EVAL_6;
  assign _EVAL_51 = _EVAL_203 | _EVAL_300;
  assign _EVAL_145 = $signed(_EVAL_55) & -33'sh400000;
  assign _EVAL_57 = _EVAL_137 | _EVAL_296;
  assign _EVAL_229 = $signed(_EVAL_342) == 33'sh0;
  assign _EVAL_290 = _EVAL_127 & _EVAL_218;
  assign _EVAL_106 = _EVAL & _EVAL_307;
  assign _EVAL_305 = _EVAL_151 | _EVAL_147;
  assign _EVAL_230 = 4'h2 == _EVAL_10;
  assign _EVAL_332 = ~_EVAL_271;
  assign _EVAL_91 = ~_EVAL_304;
  assign _EVAL_301 = _EVAL_142 | _EVAL_6;
  assign _EVAL_60 = _EVAL_89[5:0];
  assign _EVAL_65 = _EVAL_238 | _EVAL_175;
  assign _EVAL_54 = _EVAL_306 | _EVAL_6;
  assign _EVAL_270 = _EVAL_282 | _EVAL_6;
  assign _EVAL_68 = _EVAL_8 <= 2'h2;
  assign _EVAL_98 = {_EVAL_340,_EVAL_305,_EVAL_104,_EVAL_72};
  assign _EVAL_220 = _EVAL_10 == _EVAL_187;
  assign _EVAL_251 = ~_EVAL_367;
  assign _EVAL_62 = {1'b0,$signed(_EVAL_2)};
  assign _EVAL_259 = _EVAL_139 & _EVAL_251;
  assign _EVAL_156 = _EVAL_17 == 3'h2;
  assign _EVAL_338 = _EVAL_293 | _EVAL_6;
  assign _EVAL_22 = ~_EVAL_160;
  assign _EVAL_181 = _EVAL_35 | _EVAL_6;
  assign _EVAL_140 = _EVAL_124 != _EVAL_353;
  assign _EVAL_292 = $signed(_EVAL_309) == 33'sh0;
  assign _EVAL_280 = $signed(_EVAL_168) & -33'sh2000;
  assign _EVAL_200 = {1'b0,$signed(_EVAL_46)};
  assign _EVAL_344 = _EVAL_1 & _EVAL_235;
  assign _EVAL_94 = ~_EVAL_371;
  assign _EVAL_235 = _EVAL_11 == 3'h1;
  assign _EVAL_193 = ~_EVAL_162;
  assign _EVAL_50 = _EVAL_1 & _EVAL_341;
  assign _EVAL_279 = _EVAL_1 & _EVAL_333;
  assign _EVAL_372 = _EVAL_120 | _EVAL_6;
  assign _EVAL_274 = ~_EVAL_348;
  assign _EVAL_298 = ~_EVAL_302;
  assign _EVAL_356 = _EVAL_182[5:0];
  assign _EVAL_346 = $signed(_EVAL_129) & -33'sh4000;
  assign _EVAL_333 = _EVAL_11 == 3'h5;
  assign _EVAL_273 = _EVAL_328[1];
  assign _EVAL_169 = _EVAL_351 <= 3'h6;
  assign _EVAL_108 = _EVAL_11[2];
  assign _EVAL_361 = ~_EVAL_3;
  assign _EVAL_41 = ~_EVAL_139;
  assign _EVAL_364 = ~_EVAL_286;
  assign _EVAL_228 = _EVAL_1 & _EVAL_257;
  assign _EVAL_191 = _EVAL_185 | _EVAL_124;
  assign _EVAL_35 = _EVAL_303 | _EVAL_138;
  assign _EVAL_261 = _EVAL_75 | _EVAL_7;
  assign _EVAL_319 = _EVAL_255 | _EVAL_6;
  assign _EVAL_113 = $signed(_EVAL_263) & -33'sh2000;
  assign _EVAL_353 = _EVAL_188[8:0];
  assign _EVAL_197 = _EVAL_111 | _EVAL_71;
  assign _EVAL_249 = ~_EVAL_215;
  assign _EVAL_365 = ~_EVAL_226;
  assign _EVAL_103 = ~_EVAL_270;
  assign _EVAL_136 = _EVAL_113;
  assign _EVAL_26 = _EVAL_11 == 3'h3;
  assign _EVAL_195 = ~_EVAL_184;
  assign _EVAL_278 = _EVAL_127 & _EVAL_61;
  assign _EVAL_39 = ~_EVAL_125;
  assign _EVAL_63 = _EVAL_24 - 6'h1;
  assign _EVAL_283 = _EVAL_10[0];
  assign _EVAL_248 = _EVAL_27 & _EVAL_96;
  assign _EVAL_311 = _EVAL_173 == 6'h0;
  assign _EVAL_92 = _EVAL_17 <= 3'h6;
  assign _EVAL_296 = $signed(_EVAL_161) == 33'sh0;
  assign _EVAL_265 = ~_EVAL_181;
  assign _EVAL_99 = _EVAL_2 ^ 32'hc000000;
  assign _EVAL_232 = _EVAL_13 & _EVAL_1;
  assign _EVAL_225 = _EVAL_75 | _EVAL_6;
  assign _EVAL_80 = _EVAL_4 == _EVAL_369;
  assign _EVAL_73 = _EVAL_139 & _EVAL_367;
  assign _EVAL_158 = _EVAL_174 | _EVAL_6;
  assign _EVAL_72 = _EVAL_37 | _EVAL_248;
  assign _EVAL_81 = _EVAL_273 & _EVAL_139;
  assign _EVAL_201 = _EVAL_21 | _EVAL_6;
  assign _EVAL_241 = ~_EVAL_30;
  assign _EVAL_186 = _EVAL_80 | _EVAL_6;
  assign _EVAL_219 = _EVAL_191 & _EVAL_308;
  assign _EVAL_165 = _EVAL_4 <= 3'h4;
  assign _EVAL_236 = ~_EVAL_323;
  assign _EVAL_351 = _EVAL_16[2:0];
  assign _EVAL_341 = _EVAL_11 == 3'h7;
  assign _EVAL_308 = ~_EVAL_353;
  assign _EVAL_247 = _EVAL_11 == 3'h0;
  assign _EVAL_207 = _EVAL_264[0];
  assign _EVAL_231 = ~_EVAL_319;
  assign _EVAL_363 = _EVAL_2 ^ 32'h2000000;
  always @(posedge _EVAL_9) begin
    if (_EVAL_6) begin
      _EVAL_24 <= 6'h0;
    end else if (_EVAL_127) begin
      if (_EVAL_218) begin
        if (_EVAL_131) begin
          _EVAL_24 <= _EVAL_153;
        end else begin
          _EVAL_24 <= 6'h0;
        end
      end else begin
        _EVAL_24 <= _EVAL_23;
      end
    end
    if (_EVAL_315) begin
      _EVAL_67 <= _EVAL_11;
    end
    if (_EVAL_278) begin
      _EVAL_79 <= _EVAL_0;
    end
    if (_EVAL_278) begin
      _EVAL_107 <= _EVAL_8;
    end
    if (_EVAL_278) begin
      _EVAL_126 <= _EVAL_12;
    end
    if (_EVAL_6) begin
      _EVAL_163 <= 6'h0;
    end else if (_EVAL_127) begin
      if (_EVAL_61) begin
        if (_EVAL_131) begin
          _EVAL_163 <= _EVAL_153;
        end else begin
          _EVAL_163 <= 6'h0;
        end
      end else begin
        _EVAL_163 <= _EVAL_356;
      end
    end
    if (_EVAL_6) begin
      _EVAL_173 <= 6'h0;
    end else if (_EVAL_232) begin
      if (_EVAL_311) begin
        if (_EVAL_316) begin
          _EVAL_173 <= _EVAL_135;
        end else begin
          _EVAL_173 <= 6'h0;
        end
      end else begin
        _EVAL_173 <= _EVAL_60;
      end
    end
    if (_EVAL_6) begin
      _EVAL_185 <= 9'h0;
    end else begin
      _EVAL_185 <= _EVAL_219;
    end
    if (_EVAL_315) begin
      _EVAL_187 <= _EVAL_10;
    end
    if (_EVAL_6) begin
      _EVAL_189 <= 32'h0;
    end else if (_EVAL_97) begin
      _EVAL_189 <= 32'h0;
    end else begin
      _EVAL_189 <= _EVAL_284;
    end
    if (_EVAL_278) begin
      _EVAL_202 <= _EVAL_17;
    end
    if (_EVAL_315) begin
      _EVAL_258 <= _EVAL_5;
    end
    if (_EVAL_6) begin
      _EVAL_267 <= 6'h0;
    end else if (_EVAL_232) begin
      if (_EVAL_312) begin
        if (_EVAL_316) begin
          _EVAL_267 <= _EVAL_135;
        end else begin
          _EVAL_267 <= 6'h0;
        end
      end else begin
        _EVAL_267 <= _EVAL_331;
      end
    end
    if (_EVAL_315) begin
      _EVAL_334 <= _EVAL_2;
    end
    if (_EVAL_278) begin
      _EVAL_335 <= _EVAL_16;
    end
    if (_EVAL_278) begin
      _EVAL_354 <= _EVAL_15;
    end
    if (_EVAL_315) begin
      _EVAL_369 <= _EVAL_4;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eaa3103a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67ebbbca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_347) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9519c0d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL & _EVAL_275) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55485b40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_370 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a86633c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_265) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6dd8beb6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e5b5a1c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_279 & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_321) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99fbb7c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0a9cac6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_279 & _EVAL_347) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d5e5dd1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee41712d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10b717b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_236) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_357 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f59fd1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46d99b0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_294) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5834691f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee41712d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4640b5c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_321) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb547259)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL & _EVAL_275) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_279 & _EVAL_364) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6251a551)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_294) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_183) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_298) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_279 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3a4a8cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_347) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49c34e02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_357 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22401708)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_370 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5902bcbc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_347) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12c5a6a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_279 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11706b8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_279 & _EVAL_347) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(827566c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5ca23f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_279 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_279 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ae588fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_268) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_279 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cbad70ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9bdb8dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_357 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_370 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc8fcc62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_347) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(929043b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1723fb7e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_355) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b21e4d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_298) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b6ba24f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8758287)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_370 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_347) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_281) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_269) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d57cc519)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_112) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_357 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b938816a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_347) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28bdf861)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3788c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b9584e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_326) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d854495)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_279 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee80d0d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_268) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8264d8c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_347) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9db79c0b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_365) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_357 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2967af9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a2c3fa8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29b4270a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab2c2a9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_265) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8739fa9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e77f022)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_370 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14ca317d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c35707e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10a38d4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5864a3b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_236) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3e7a266)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_281) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a653170)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb8dfe9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_134) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24382ad1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d58d5bdc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7103c34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4b8465f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_167) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bce3eb99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdb122da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_357 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23d17dba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_279 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_355) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_357 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d99995cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_370 & _EVAL_347) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a4ee769)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_152) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_183) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf43e39d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_152) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28446467)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_357 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_279 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8ad87b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8fb4e951)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_370 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d984ef1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_357 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9e2047b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_347) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0e7af38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_347) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9dbbf1c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74cdbec6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_144 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_347) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c18d74cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_294) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_195) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(def2ad62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_357 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_269) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_357 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6bad9fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_294) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(deeb006c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_357 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91155d42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_370 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(717bd96d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_347) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_59 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e109d7be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd2dec62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_195) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8561a5b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8799821a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_279 & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82538676)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b83f58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_365) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d7c32ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_279 & _EVAL_364) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_347) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73db08d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_228 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3510675d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_326) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ec335d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_370 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_112) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f5e8ecd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_370 & _EVAL_347) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc978fbd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_245 & _EVAL_134) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_24 = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_67 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_79 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_107 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_126 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_163 = _RAND_5[5:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_173 = _RAND_6[5:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_185 = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_187 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_189 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_202 = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_258 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_267 = _RAND_12[5:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_334 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_335 = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_354 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_369 = _RAND_16[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
