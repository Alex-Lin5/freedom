//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_94(
  output [31:0] _EVAL,
  output [31:0] _EVAL_0,
  output [31:0] _EVAL_1,
  output [4:0]  _EVAL_2,
  output        _EVAL_3,
  input  [2:0]  _EVAL_4,
  input  [4:0]  _EVAL_5,
  output [2:0]  _EVAL_6,
  output [1:0]  _EVAL_7,
  output [11:0] _EVAL_8,
  input  [1:0]  _EVAL_9,
  output [1:0]  _EVAL_10,
  input         _EVAL_11,
  output [3:0]  _EVAL_12,
  output        _EVAL_13,
  output [31:0] _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  output        _EVAL_17,
  input         _EVAL_18,
  input  [31:0] _EVAL_19,
  output [3:0]  _EVAL_20,
  output [9:0]  _EVAL_21,
  output [1:0]  _EVAL_22,
  input  [2:0]  _EVAL_23,
  input  [31:0] _EVAL_24,
  output [1:0]  _EVAL_25,
  input  [3:0]  _EVAL_26,
  input         _EVAL_27,
  input  [2:0]  _EVAL_28,
  output [2:0]  _EVAL_29,
  input  [2:0]  _EVAL_30,
  output [2:0]  _EVAL_31,
  input  [31:0] _EVAL_32,
  output [9:0]  _EVAL_33,
  input  [4:0]  _EVAL_34,
  input         _EVAL_35,
  input  [31:0] _EVAL_36,
  output [2:0]  _EVAL_37,
  output [2:0]  _EVAL_38,
  output        _EVAL_39,
  input         _EVAL_40,
  output [2:0]  _EVAL_41,
  input  [2:0]  _EVAL_42,
  output        _EVAL_43,
  output [4:0]  _EVAL_44,
  output [14:0] _EVAL_45,
  output        _EVAL_46,
  output        _EVAL_47,
  output [2:0]  _EVAL_48,
  input  [31:0] _EVAL_49,
  input         _EVAL_50,
  input  [9:0]  _EVAL_51,
  output [3:0]  _EVAL_52,
  output [9:0]  _EVAL_53,
  output [2:0]  _EVAL_54,
  input         _EVAL_55,
  input         _EVAL_56,
  output [1:0]  _EVAL_57,
  output        _EVAL_58,
  input         _EVAL_59,
  input  [1:0]  _EVAL_60,
  input  [3:0]  _EVAL_61,
  input  [1:0]  _EVAL_62,
  input  [2:0]  _EVAL_63,
  output        _EVAL_64,
  output        _EVAL_65,
  output        _EVAL_66,
  input  [2:0]  _EVAL_67,
  input  [31:0] _EVAL_68,
  output [4:0]  _EVAL_69,
  input         _EVAL_70,
  output        _EVAL_71,
  output [1:0]  _EVAL_72,
  output [1:0]  _EVAL_73,
  input  [9:0]  _EVAL_74,
  input         _EVAL_75,
  input         _EVAL_76,
  output [25:0] _EVAL_77,
  output        _EVAL_78,
  output [31:0] _EVAL_79,
  input         _EVAL_80,
  output [27:0] _EVAL_81,
  input         _EVAL_82,
  input  [31:0] _EVAL_83,
  output [3:0]  _EVAL_84,
  input  [4:0]  _EVAL_85,
  output        _EVAL_86,
  output [2:0]  _EVAL_87,
  output [2:0]  _EVAL_88,
  output        _EVAL_89,
  output [2:0]  _EVAL_90,
  output        _EVAL_91,
  output [31:0] _EVAL_92,
  output [3:0]  _EVAL_93,
  input  [2:0]  _EVAL_94,
  output        _EVAL_95,
  input         _EVAL_96,
  output        _EVAL_97,
  input  [1:0]  _EVAL_98,
  output        _EVAL_99,
  output [2:0]  _EVAL_100,
  output [31:0] _EVAL_101,
  output        _EVAL_102,
  output [31:0] _EVAL_103,
  input  [1:0]  _EVAL_104,
  output [29:0] _EVAL_105,
  output [1:0]  _EVAL_106,
  input  [1:0]  _EVAL_107,
  output [2:0]  _EVAL_108,
  output        _EVAL_109,
  output [31:0] _EVAL_110,
  output [2:0]  _EVAL_111,
  output        _EVAL_112,
  input         _EVAL_113,
  input  [2:0]  _EVAL_114,
  output [31:0] _EVAL_115,
  output [2:0]  _EVAL_116,
  output [3:0]  _EVAL_117,
  input  [9:0]  _EVAL_118,
  input  [31:0] _EVAL_119,
  input         _EVAL_120,
  output [3:0]  _EVAL_121,
  input  [2:0]  _EVAL_122,
  input  [9:0]  _EVAL_123,
  output [9:0]  _EVAL_124,
  output        _EVAL_125,
  input  [31:0] _EVAL_126,
  output [3:0]  _EVAL_127,
  input         _EVAL_128,
  output        _EVAL_129,
  output        _EVAL_130,
  output [2:0]  _EVAL_131,
  output        _EVAL_132,
  input         _EVAL_133
);
  wire [31:0] _EVAL_134;
  wire [2:0] atomics__EVAL;
  wire [2:0] atomics__EVAL_0;
  wire  atomics__EVAL_1;
  wire [4:0] atomics__EVAL_2;
  wire [1:0] atomics__EVAL_3;
  wire  atomics__EVAL_4;
  wire [4:0] atomics__EVAL_5;
  wire [3:0] atomics__EVAL_6;
  wire  atomics__EVAL_7;
  wire  atomics__EVAL_8;
  wire [31:0] atomics__EVAL_9;
  wire [31:0] atomics__EVAL_10;
  wire  atomics__EVAL_11;
  wire [2:0] atomics__EVAL_12;
  wire [2:0] atomics__EVAL_13;
  wire [2:0] atomics__EVAL_14;
  wire  atomics__EVAL_15;
  wire  atomics__EVAL_16;
  wire  atomics__EVAL_17;
  wire [2:0] atomics__EVAL_18;
  wire  atomics__EVAL_19;
  wire  atomics__EVAL_20;
  wire  atomics__EVAL_21;
  wire [3:0] atomics__EVAL_22;
  wire [31:0] atomics__EVAL_23;
  wire  atomics__EVAL_24;
  wire [31:0] atomics__EVAL_25;
  wire  atomics__EVAL_26;
  wire  atomics__EVAL_27;
  wire [1:0] atomics__EVAL_28;
  wire [4:0] atomics__EVAL_29;
  wire [3:0] atomics__EVAL_30;
  wire  atomics__EVAL_31;
  wire [3:0] atomics__EVAL_32;
  wire  atomics__EVAL_33;
  wire  atomics__EVAL_34;
  wire  atomics__EVAL_35;
  wire [31:0] atomics__EVAL_36;
  wire [4:0] atomics__EVAL_37;
  wire  atomics__EVAL_38;
  wire  atomics__EVAL_39;
  wire  atomics__EVAL_40;
  wire [31:0] atomics__EVAL_41;
  wire  atomics__EVAL_42;
  wire  atomics__EVAL_43;
  wire  atomics__EVAL_44;
  wire [3:0] atomics__EVAL_45;
  wire [3:0] atomics__EVAL_46;
  wire  atomics__EVAL_47;
  wire  atomics__EVAL_48;
  wire [4:0] _EVAL_135;
  wire [2:0] coupler_to_clint__EVAL;
  wire [2:0] coupler_to_clint__EVAL_0;
  wire [3:0] coupler_to_clint__EVAL_1;
  wire [2:0] coupler_to_clint__EVAL_2;
  wire  coupler_to_clint__EVAL_3;
  wire [4:0] coupler_to_clint__EVAL_4;
  wire  coupler_to_clint__EVAL_5;
  wire [9:0] coupler_to_clint__EVAL_6;
  wire  coupler_to_clint__EVAL_7;
  wire [2:0] coupler_to_clint__EVAL_8;
  wire  coupler_to_clint__EVAL_9;
  wire  coupler_to_clint__EVAL_10;
  wire [2:0] coupler_to_clint__EVAL_11;
  wire [31:0] coupler_to_clint__EVAL_12;
  wire  coupler_to_clint__EVAL_13;
  wire [31:0] coupler_to_clint__EVAL_14;
  wire  coupler_to_clint__EVAL_15;
  wire [31:0] coupler_to_clint__EVAL_16;
  wire [2:0] coupler_to_clint__EVAL_17;
  wire [2:0] coupler_to_clint__EVAL_18;
  wire [31:0] coupler_to_clint__EVAL_19;
  wire  coupler_to_clint__EVAL_20;
  wire  coupler_to_clint__EVAL_21;
  wire [3:0] coupler_to_clint__EVAL_22;
  wire [2:0] coupler_to_clint__EVAL_23;
  wire [1:0] coupler_to_clint__EVAL_24;
  wire [4:0] coupler_to_clint__EVAL_25;
  wire  coupler_to_clint__EVAL_26;
  wire [1:0] coupler_to_clint__EVAL_27;
  wire  coupler_to_clint__EVAL_28;
  wire [9:0] coupler_to_clint__EVAL_29;
  wire [25:0] coupler_to_clint__EVAL_30;
  wire [25:0] coupler_to_clint__EVAL_31;
  wire  coupler_to_clint__EVAL_32;
  wire  wrapped_error_device__EVAL;
  wire [3:0] wrapped_error_device__EVAL_0;
  wire [13:0] wrapped_error_device__EVAL_1;
  wire [2:0] wrapped_error_device__EVAL_2;
  wire [3:0] wrapped_error_device__EVAL_3;
  wire [3:0] wrapped_error_device__EVAL_4;
  wire  wrapped_error_device__EVAL_5;
  wire [31:0] wrapped_error_device__EVAL_6;
  wire [4:0] wrapped_error_device__EVAL_7;
  wire [1:0] wrapped_error_device__EVAL_8;
  wire [2:0] wrapped_error_device__EVAL_9;
  wire [2:0] wrapped_error_device__EVAL_10;
  wire  wrapped_error_device__EVAL_11;
  wire  wrapped_error_device__EVAL_12;
  wire  wrapped_error_device__EVAL_13;
  wire  wrapped_error_device__EVAL_14;
  wire  wrapped_error_device__EVAL_15;
  wire [4:0] wrapped_error_device__EVAL_16;
  wire  wrapped_error_device__EVAL_17;
  wire  wrapped_error_device__EVAL_18;
  wire  wrapped_error_device__EVAL_19;
  wire  _EVAL_136;
  wire [4:0] _EVAL_137;
  wire  _EVAL_138;
  wire [31:0] coupler_to_tile__EVAL;
  wire [2:0] coupler_to_tile__EVAL_0;
  wire [1:0] coupler_to_tile__EVAL_1;
  wire  coupler_to_tile__EVAL_2;
  wire [4:0] coupler_to_tile__EVAL_3;
  wire [31:0] coupler_to_tile__EVAL_4;
  wire [2:0] coupler_to_tile__EVAL_5;
  wire [2:0] coupler_to_tile__EVAL_6;
  wire [4:0] coupler_to_tile__EVAL_7;
  wire [2:0] coupler_to_tile__EVAL_8;
  wire  coupler_to_tile__EVAL_9;
  wire [4:0] coupler_to_tile__EVAL_10;
  wire [3:0] coupler_to_tile__EVAL_11;
  wire [2:0] coupler_to_tile__EVAL_12;
  wire [4:0] coupler_to_tile__EVAL_13;
  wire [1:0] coupler_to_tile__EVAL_14;
  wire  coupler_to_tile__EVAL_15;
  wire  coupler_to_tile__EVAL_16;
  wire  coupler_to_tile__EVAL_17;
  wire [2:0] coupler_to_tile__EVAL_18;
  wire [4:0] coupler_to_tile__EVAL_19;
  wire [31:0] coupler_to_tile__EVAL_20;
  wire  coupler_to_tile__EVAL_21;
  wire [3:0] coupler_to_tile__EVAL_22;
  wire [31:0] coupler_to_tile__EVAL_23;
  wire [3:0] coupler_to_tile__EVAL_24;
  wire [31:0] coupler_to_tile__EVAL_25;
  wire  coupler_to_tile__EVAL_26;
  wire [31:0] coupler_to_tile__EVAL_27;
  wire [31:0] coupler_to_tile__EVAL_28;
  wire [2:0] coupler_to_tile__EVAL_29;
  wire [2:0] coupler_to_tile__EVAL_30;
  wire  coupler_to_tile__EVAL_31;
  wire [31:0] coupler_to_tile__EVAL_32;
  wire [2:0] coupler_to_tile__EVAL_33;
  wire [1:0] coupler_to_tile__EVAL_34;
  wire  coupler_to_tile__EVAL_35;
  wire [2:0] coupler_to_tile__EVAL_36;
  wire [31:0] coupler_to_tile__EVAL_37;
  wire [2:0] coupler_to_tile__EVAL_38;
  wire [2:0] coupler_to_tile__EVAL_39;
  wire [2:0] coupler_to_tile__EVAL_40;
  wire [1:0] coupler_to_tile__EVAL_41;
  wire  coupler_to_tile__EVAL_42;
  wire [2:0] coupler_to_tile__EVAL_43;
  wire [4:0] coupler_to_tile__EVAL_44;
  wire [2:0] coupler_to_tile__EVAL_45;
  wire [2:0] _EVAL_139;
  wire [2:0] _EVAL_140;
  wire  _EVAL_141;
  wire [2:0] _EVAL_142;
  wire [3:0] buffer__EVAL;
  wire  buffer__EVAL_0;
  wire  buffer__EVAL_1;
  wire  buffer__EVAL_2;
  wire  buffer__EVAL_3;
  wire  buffer__EVAL_4;
  wire [4:0] buffer__EVAL_5;
  wire  buffer__EVAL_6;
  wire [4:0] buffer__EVAL_7;
  wire  buffer__EVAL_8;
  wire  buffer__EVAL_9;
  wire [3:0] buffer__EVAL_10;
  wire [31:0] buffer__EVAL_11;
  wire  buffer__EVAL_12;
  wire [2:0] buffer__EVAL_13;
  wire [1:0] buffer__EVAL_14;
  wire  buffer__EVAL_15;
  wire  buffer__EVAL_16;
  wire [4:0] buffer__EVAL_17;
  wire  buffer__EVAL_18;
  wire [2:0] buffer__EVAL_19;
  wire [2:0] buffer__EVAL_20;
  wire [31:0] buffer__EVAL_21;
  wire  buffer__EVAL_22;
  wire  buffer__EVAL_23;
  wire  buffer__EVAL_24;
  wire  buffer__EVAL_25;
  wire  buffer__EVAL_26;
  wire [3:0] buffer__EVAL_27;
  wire [4:0] buffer__EVAL_28;
  wire  buffer__EVAL_29;
  wire [31:0] buffer__EVAL_30;
  wire  buffer__EVAL_31;
  wire  buffer__EVAL_32;
  wire [31:0] buffer__EVAL_33;
  wire [2:0] buffer__EVAL_34;
  wire  buffer__EVAL_35;
  wire  buffer__EVAL_36;
  wire [1:0] buffer__EVAL_37;
  wire [2:0] buffer__EVAL_38;
  wire [3:0] buffer__EVAL_39;
  wire [31:0] buffer__EVAL_40;
  wire  buffer__EVAL_41;
  wire [3:0] buffer__EVAL_42;
  wire  buffer__EVAL_43;
  wire  buffer__EVAL_44;
  wire [3:0] buffer__EVAL_45;
  wire [2:0] buffer__EVAL_46;
  wire [31:0] buffer__EVAL_47;
  wire  buffer__EVAL_48;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire [3:0] _EVAL_147;
  wire [3:0] _EVAL_148;
  wire  _EVAL_149;
  wire [2:0] _EVAL_150;
  wire [2:0] _EVAL_151;
  wire  _EVAL_152;
  wire [31:0] _EVAL_153;
  wire [2:0] _EVAL_154;
  wire [3:0] _EVAL_155;
  wire [4:0] _EVAL_156;
  wire [2:0] _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire [4:0] _EVAL_161;
  wire  out_xbar__EVAL;
  wire [2:0] out_xbar__EVAL_0;
  wire  out_xbar__EVAL_1;
  wire [3:0] out_xbar__EVAL_2;
  wire  out_xbar__EVAL_3;
  wire [11:0] out_xbar__EVAL_4;
  wire [2:0] out_xbar__EVAL_5;
  wire [4:0] out_xbar__EVAL_6;
  wire  out_xbar__EVAL_7;
  wire [3:0] out_xbar__EVAL_8;
  wire [4:0] out_xbar__EVAL_9;
  wire  out_xbar__EVAL_10;
  wire [2:0] out_xbar__EVAL_11;
  wire [31:0] out_xbar__EVAL_12;
  wire [14:0] out_xbar__EVAL_13;
  wire [4:0] out_xbar__EVAL_14;
  wire [1:0] out_xbar__EVAL_15;
  wire [2:0] out_xbar__EVAL_16;
  wire [31:0] out_xbar__EVAL_17;
  wire  out_xbar__EVAL_18;
  wire  out_xbar__EVAL_19;
  wire  out_xbar__EVAL_20;
  wire [31:0] out_xbar__EVAL_21;
  wire  out_xbar__EVAL_22;
  wire  out_xbar__EVAL_23;
  wire [31:0] out_xbar__EVAL_24;
  wire  out_xbar__EVAL_25;
  wire  out_xbar__EVAL_26;
  wire [3:0] out_xbar__EVAL_27;
  wire [1:0] out_xbar__EVAL_28;
  wire  out_xbar__EVAL_29;
  wire [4:0] out_xbar__EVAL_30;
  wire  out_xbar__EVAL_31;
  wire [4:0] out_xbar__EVAL_32;
  wire  out_xbar__EVAL_33;
  wire [2:0] out_xbar__EVAL_34;
  wire  out_xbar__EVAL_35;
  wire [1:0] out_xbar__EVAL_36;
  wire  out_xbar__EVAL_37;
  wire  out_xbar__EVAL_38;
  wire [2:0] out_xbar__EVAL_39;
  wire  out_xbar__EVAL_40;
  wire  out_xbar__EVAL_41;
  wire [25:0] out_xbar__EVAL_42;
  wire [3:0] out_xbar__EVAL_43;
  wire  out_xbar__EVAL_44;
  wire  out_xbar__EVAL_45;
  wire [2:0] out_xbar__EVAL_46;
  wire [2:0] out_xbar__EVAL_47;
  wire  out_xbar__EVAL_48;
  wire [3:0] out_xbar__EVAL_49;
  wire  out_xbar__EVAL_50;
  wire [2:0] out_xbar__EVAL_51;
  wire  out_xbar__EVAL_52;
  wire [31:0] out_xbar__EVAL_53;
  wire  out_xbar__EVAL_54;
  wire  out_xbar__EVAL_55;
  wire [2:0] out_xbar__EVAL_56;
  wire [2:0] out_xbar__EVAL_57;
  wire  out_xbar__EVAL_58;
  wire [2:0] out_xbar__EVAL_59;
  wire  out_xbar__EVAL_60;
  wire  out_xbar__EVAL_61;
  wire [2:0] out_xbar__EVAL_62;
  wire [3:0] out_xbar__EVAL_63;
  wire [3:0] out_xbar__EVAL_64;
  wire [31:0] out_xbar__EVAL_65;
  wire  out_xbar__EVAL_66;
  wire  out_xbar__EVAL_67;
  wire  out_xbar__EVAL_68;
  wire [2:0] out_xbar__EVAL_69;
  wire  out_xbar__EVAL_70;
  wire  out_xbar__EVAL_71;
  wire [4:0] out_xbar__EVAL_72;
  wire [27:0] out_xbar__EVAL_73;
  wire [31:0] out_xbar__EVAL_74;
  wire  out_xbar__EVAL_75;
  wire  out_xbar__EVAL_76;
  wire [31:0] out_xbar__EVAL_77;
  wire [2:0] out_xbar__EVAL_78;
  wire [2:0] out_xbar__EVAL_79;
  wire  out_xbar__EVAL_80;
  wire [4:0] out_xbar__EVAL_81;
  wire  out_xbar__EVAL_82;
  wire [2:0] out_xbar__EVAL_83;
  wire  out_xbar__EVAL_84;
  wire  out_xbar__EVAL_85;
  wire  out_xbar__EVAL_86;
  wire [31:0] out_xbar__EVAL_87;
  wire  out_xbar__EVAL_88;
  wire [2:0] out_xbar__EVAL_89;
  wire  out_xbar__EVAL_90;
  wire [31:0] out_xbar__EVAL_91;
  wire [2:0] out_xbar__EVAL_92;
  wire [4:0] out_xbar__EVAL_93;
  wire [2:0] out_xbar__EVAL_94;
  wire [2:0] out_xbar__EVAL_95;
  wire [2:0] out_xbar__EVAL_96;
  wire  out_xbar__EVAL_97;
  wire  out_xbar__EVAL_98;
  wire [31:0] out_xbar__EVAL_99;
  wire  out_xbar__EVAL_100;
  wire [2:0] out_xbar__EVAL_101;
  wire [2:0] out_xbar__EVAL_102;
  wire  out_xbar__EVAL_103;
  wire [4:0] out_xbar__EVAL_104;
  wire [31:0] out_xbar__EVAL_105;
  wire [2:0] out_xbar__EVAL_106;
  wire [2:0] out_xbar__EVAL_107;
  wire [3:0] out_xbar__EVAL_108;
  wire  out_xbar__EVAL_109;
  wire [4:0] out_xbar__EVAL_110;
  wire [2:0] out_xbar__EVAL_111;
  wire [31:0] out_xbar__EVAL_112;
  wire [3:0] out_xbar__EVAL_113;
  wire [3:0] out_xbar__EVAL_114;
  wire [2:0] out_xbar__EVAL_115;
  wire [4:0] out_xbar__EVAL_116;
  wire [2:0] out_xbar__EVAL_117;
  wire [2:0] out_xbar__EVAL_118;
  wire [4:0] out_xbar__EVAL_119;
  wire  out_xbar__EVAL_120;
  wire [2:0] out_xbar__EVAL_121;
  wire  out_xbar__EVAL_122;
  wire [2:0] out_xbar__EVAL_123;
  wire [4:0] out_xbar__EVAL_124;
  wire  out_xbar__EVAL_125;
  wire [13:0] out_xbar__EVAL_126;
  wire [2:0] out_xbar__EVAL_127;
  wire  out_xbar__EVAL_128;
  wire [29:0] out_xbar__EVAL_129;
  wire [3:0] out_xbar__EVAL_130;
  wire [4:0] out_xbar__EVAL_131;
  wire  out_xbar__EVAL_132;
  wire  out_xbar__EVAL_133;
  wire [2:0] out_xbar__EVAL_134;
  wire [3:0] out_xbar__EVAL_135;
  wire [2:0] out_xbar__EVAL_136;
  wire [4:0] out_xbar__EVAL_137;
  wire [31:0] out_xbar__EVAL_138;
  wire [31:0] out_xbar__EVAL_139;
  wire  out_xbar__EVAL_140;
  wire [4:0] out_xbar__EVAL_141;
  wire [2:0] out_xbar__EVAL_142;
  wire  out_xbar__EVAL_143;
  wire [31:0] out_xbar__EVAL_144;
  wire [31:0] out_xbar__EVAL_145;
  wire  out_xbar__EVAL_146;
  wire  _EVAL_162;
  wire [31:0] _EVAL_163;
  wire [2:0] _EVAL_164;
  wire  _EVAL_165;
  wire [31:0] _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire [2:0] _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire [31:0] _EVAL_172;
  wire  _EVAL_173;
  wire [3:0] _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire [31:0] _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire [31:0] _EVAL_181;
  wire [2:0] _EVAL_182;
  wire [31:0] _EVAL_183;
  wire  _EVAL_184;
  wire  coupler_to_debug__EVAL;
  wire [2:0] coupler_to_debug__EVAL_0;
  wire  coupler_to_debug__EVAL_1;
  wire [2:0] coupler_to_debug__EVAL_2;
  wire [2:0] coupler_to_debug__EVAL_3;
  wire  coupler_to_debug__EVAL_4;
  wire  coupler_to_debug__EVAL_5;
  wire [9:0] coupler_to_debug__EVAL_6;
  wire  coupler_to_debug__EVAL_7;
  wire [1:0] coupler_to_debug__EVAL_8;
  wire  coupler_to_debug__EVAL_9;
  wire [31:0] coupler_to_debug__EVAL_10;
  wire [2:0] coupler_to_debug__EVAL_11;
  wire  coupler_to_debug__EVAL_12;
  wire [2:0] coupler_to_debug__EVAL_13;
  wire [4:0] coupler_to_debug__EVAL_14;
  wire  coupler_to_debug__EVAL_15;
  wire [1:0] coupler_to_debug__EVAL_16;
  wire  coupler_to_debug__EVAL_17;
  wire [2:0] coupler_to_debug__EVAL_18;
  wire [3:0] coupler_to_debug__EVAL_19;
  wire [11:0] coupler_to_debug__EVAL_20;
  wire [4:0] coupler_to_debug__EVAL_21;
  wire  coupler_to_debug__EVAL_22;
  wire  coupler_to_debug__EVAL_23;
  wire [2:0] coupler_to_debug__EVAL_24;
  wire [31:0] coupler_to_debug__EVAL_25;
  wire [31:0] coupler_to_debug__EVAL_26;
  wire [11:0] coupler_to_debug__EVAL_27;
  wire [2:0] coupler_to_debug__EVAL_28;
  wire [31:0] coupler_to_debug__EVAL_29;
  wire [3:0] coupler_to_debug__EVAL_30;
  wire  coupler_to_debug__EVAL_31;
  wire [9:0] coupler_to_debug__EVAL_32;
  wire  fixedClockNode__EVAL;
  wire  fixedClockNode__EVAL_0;
  wire  fixedClockNode__EVAL_1;
  wire  fixedClockNode__EVAL_2;
  wire  fixedClockNode__EVAL_3;
  wire  fixedClockNode__EVAL_4;
  wire  fixedClockNode__EVAL_5;
  wire  fixedClockNode__EVAL_6;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire [3:0] _EVAL_188;
  wire  _EVAL_189;
  wire  coupler_to_port_named_ahb_periph_port__EVAL;
  wire [2:0] coupler_to_port_named_ahb_periph_port__EVAL_0;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_1;
  wire [29:0] coupler_to_port_named_ahb_periph_port__EVAL_2;
  wire [3:0] coupler_to_port_named_ahb_periph_port__EVAL_3;
  wire [2:0] coupler_to_port_named_ahb_periph_port__EVAL_4;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_5;
  wire [31:0] coupler_to_port_named_ahb_periph_port__EVAL_6;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_7;
  wire [2:0] coupler_to_port_named_ahb_periph_port__EVAL_8;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_9;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_10;
  wire [4:0] coupler_to_port_named_ahb_periph_port__EVAL_11;
  wire [31:0] coupler_to_port_named_ahb_periph_port__EVAL_12;
  wire [2:0] coupler_to_port_named_ahb_periph_port__EVAL_13;
  wire [2:0] coupler_to_port_named_ahb_periph_port__EVAL_14;
  wire [1:0] coupler_to_port_named_ahb_periph_port__EVAL_15;
  wire [4:0] coupler_to_port_named_ahb_periph_port__EVAL_16;
  wire [31:0] coupler_to_port_named_ahb_periph_port__EVAL_17;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_18;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_19;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_20;
  wire [29:0] coupler_to_port_named_ahb_periph_port__EVAL_21;
  wire [3:0] coupler_to_port_named_ahb_periph_port__EVAL_22;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_23;
  wire [1:0] coupler_to_port_named_ahb_periph_port__EVAL_24;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_25;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_26;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_27;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_28;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_29;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_30;
  wire [31:0] coupler_to_port_named_ahb_periph_port__EVAL_31;
  wire [2:0] coupler_to_port_named_ahb_periph_port__EVAL_32;
  wire  coupler_to_port_named_ahb_periph_port__EVAL_33;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire [31:0] _EVAL_196;
  wire [3:0] _EVAL_197;
  wire [3:0] fixer__EVAL;
  wire [31:0] fixer__EVAL_0;
  wire  fixer__EVAL_1;
  wire  fixer__EVAL_2;
  wire  fixer__EVAL_3;
  wire  fixer__EVAL_4;
  wire  fixer__EVAL_5;
  wire [1:0] fixer__EVAL_6;
  wire  fixer__EVAL_7;
  wire  fixer__EVAL_8;
  wire [3:0] fixer__EVAL_9;
  wire [2:0] fixer__EVAL_10;
  wire  fixer__EVAL_11;
  wire  fixer__EVAL_12;
  wire [3:0] fixer__EVAL_13;
  wire  fixer__EVAL_14;
  wire  fixer__EVAL_15;
  wire [31:0] fixer__EVAL_16;
  wire [4:0] fixer__EVAL_17;
  wire [31:0] fixer__EVAL_18;
  wire  fixer__EVAL_19;
  wire [4:0] fixer__EVAL_20;
  wire [31:0] fixer__EVAL_21;
  wire  fixer__EVAL_22;
  wire  fixer__EVAL_23;
  wire [31:0] fixer__EVAL_24;
  wire [2:0] fixer__EVAL_25;
  wire [2:0] fixer__EVAL_26;
  wire [4:0] fixer__EVAL_27;
  wire  fixer__EVAL_28;
  wire [3:0] fixer__EVAL_29;
  wire [2:0] fixer__EVAL_30;
  wire [2:0] fixer__EVAL_31;
  wire [31:0] fixer__EVAL_32;
  wire [3:0] fixer__EVAL_33;
  wire  fixer__EVAL_34;
  wire  fixer__EVAL_35;
  wire  fixer__EVAL_36;
  wire  fixer__EVAL_37;
  wire [1:0] fixer__EVAL_38;
  wire  fixer__EVAL_39;
  wire  fixer__EVAL_40;
  wire  fixer__EVAL_41;
  wire [3:0] fixer__EVAL_42;
  wire  fixer__EVAL_43;
  wire  fixer__EVAL_44;
  wire  fixer__EVAL_45;
  wire [4:0] fixer__EVAL_46;
  wire [2:0] fixer__EVAL_47;
  wire  fixer__EVAL_48;
  wire  _EVAL_198;
  wire [3:0] _EVAL_199;
  wire [1:0] _EVAL_200;
  wire  _EVAL_201;
  wire [4:0] _EVAL_202;
  wire [1:0] _EVAL_203;
  wire [2:0] _EVAL_204;
  wire  _EVAL_205;
  wire [3:0] _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire [4:0] _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  coupler_to_testIndicator__EVAL;
  wire [2:0] coupler_to_testIndicator__EVAL_0;
  wire [3:0] coupler_to_testIndicator__EVAL_1;
  wire [1:0] coupler_to_testIndicator__EVAL_2;
  wire [31:0] coupler_to_testIndicator__EVAL_3;
  wire  coupler_to_testIndicator__EVAL_4;
  wire  coupler_to_testIndicator__EVAL_5;
  wire  coupler_to_testIndicator__EVAL_6;
  wire [2:0] coupler_to_testIndicator__EVAL_7;
  wire  coupler_to_testIndicator__EVAL_8;
  wire  coupler_to_testIndicator__EVAL_9;
  wire [31:0] coupler_to_testIndicator__EVAL_10;
  wire  coupler_to_testIndicator__EVAL_11;
  wire [14:0] coupler_to_testIndicator__EVAL_12;
  wire [2:0] coupler_to_testIndicator__EVAL_13;
  wire [4:0] coupler_to_testIndicator__EVAL_14;
  wire [14:0] coupler_to_testIndicator__EVAL_15;
  wire  coupler_to_testIndicator__EVAL_16;
  wire [9:0] coupler_to_testIndicator__EVAL_17;
  wire  coupler_to_testIndicator__EVAL_18;
  wire [4:0] coupler_to_testIndicator__EVAL_19;
  wire [2:0] coupler_to_testIndicator__EVAL_20;
  wire [2:0] coupler_to_testIndicator__EVAL_21;
  wire [3:0] coupler_to_testIndicator__EVAL_22;
  wire  coupler_to_testIndicator__EVAL_23;
  wire [31:0] coupler_to_testIndicator__EVAL_24;
  wire [9:0] coupler_to_testIndicator__EVAL_25;
  wire [2:0] coupler_to_testIndicator__EVAL_26;
  wire [31:0] coupler_to_testIndicator__EVAL_27;
  wire [2:0] coupler_to_testIndicator__EVAL_28;
  wire  coupler_to_testIndicator__EVAL_29;
  wire [2:0] coupler_to_testIndicator__EVAL_30;
  wire [1:0] coupler_to_testIndicator__EVAL_31;
  wire  coupler_to_testIndicator__EVAL_32;
  wire [1:0] _EVAL_212;
  wire [2:0] _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire [4:0] _EVAL_217;
  wire  _EVAL_218;
  wire [4:0] _EVAL_219;
  wire [31:0] _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire [3:0] _EVAL_223;
  wire  _EVAL_224;
  wire  coupler_to_plic__EVAL;
  wire [9:0] coupler_to_plic__EVAL_0;
  wire  coupler_to_plic__EVAL_1;
  wire  coupler_to_plic__EVAL_2;
  wire [31:0] coupler_to_plic__EVAL_3;
  wire  coupler_to_plic__EVAL_4;
  wire [2:0] coupler_to_plic__EVAL_5;
  wire [27:0] coupler_to_plic__EVAL_6;
  wire [2:0] coupler_to_plic__EVAL_7;
  wire [31:0] coupler_to_plic__EVAL_8;
  wire [2:0] coupler_to_plic__EVAL_9;
  wire [9:0] coupler_to_plic__EVAL_10;
  wire [3:0] coupler_to_plic__EVAL_11;
  wire [1:0] coupler_to_plic__EVAL_12;
  wire [2:0] coupler_to_plic__EVAL_13;
  wire [2:0] coupler_to_plic__EVAL_14;
  wire [2:0] coupler_to_plic__EVAL_15;
  wire  coupler_to_plic__EVAL_16;
  wire [2:0] coupler_to_plic__EVAL_17;
  wire [2:0] coupler_to_plic__EVAL_18;
  wire [31:0] coupler_to_plic__EVAL_19;
  wire [31:0] coupler_to_plic__EVAL_20;
  wire  coupler_to_plic__EVAL_21;
  wire [1:0] coupler_to_plic__EVAL_22;
  wire  coupler_to_plic__EVAL_23;
  wire  coupler_to_plic__EVAL_24;
  wire [4:0] coupler_to_plic__EVAL_25;
  wire [27:0] coupler_to_plic__EVAL_26;
  wire  coupler_to_plic__EVAL_27;
  wire [3:0] coupler_to_plic__EVAL_28;
  wire  coupler_to_plic__EVAL_29;
  wire [4:0] coupler_to_plic__EVAL_30;
  wire  coupler_to_plic__EVAL_31;
  wire  coupler_to_plic__EVAL_32;
  wire [31:0] _EVAL_225;
  wire [3:0] _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire [31:0] _EVAL_230;
  wire [3:0] _EVAL_231;
  wire [3:0] _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire [1:0] _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  _EVAL_52 atomics (
    ._EVAL(atomics__EVAL),
    ._EVAL_0(atomics__EVAL_0),
    ._EVAL_1(atomics__EVAL_1),
    ._EVAL_2(atomics__EVAL_2),
    ._EVAL_3(atomics__EVAL_3),
    ._EVAL_4(atomics__EVAL_4),
    ._EVAL_5(atomics__EVAL_5),
    ._EVAL_6(atomics__EVAL_6),
    ._EVAL_7(atomics__EVAL_7),
    ._EVAL_8(atomics__EVAL_8),
    ._EVAL_9(atomics__EVAL_9),
    ._EVAL_10(atomics__EVAL_10),
    ._EVAL_11(atomics__EVAL_11),
    ._EVAL_12(atomics__EVAL_12),
    ._EVAL_13(atomics__EVAL_13),
    ._EVAL_14(atomics__EVAL_14),
    ._EVAL_15(atomics__EVAL_15),
    ._EVAL_16(atomics__EVAL_16),
    ._EVAL_17(atomics__EVAL_17),
    ._EVAL_18(atomics__EVAL_18),
    ._EVAL_19(atomics__EVAL_19),
    ._EVAL_20(atomics__EVAL_20),
    ._EVAL_21(atomics__EVAL_21),
    ._EVAL_22(atomics__EVAL_22),
    ._EVAL_23(atomics__EVAL_23),
    ._EVAL_24(atomics__EVAL_24),
    ._EVAL_25(atomics__EVAL_25),
    ._EVAL_26(atomics__EVAL_26),
    ._EVAL_27(atomics__EVAL_27),
    ._EVAL_28(atomics__EVAL_28),
    ._EVAL_29(atomics__EVAL_29),
    ._EVAL_30(atomics__EVAL_30),
    ._EVAL_31(atomics__EVAL_31),
    ._EVAL_32(atomics__EVAL_32),
    ._EVAL_33(atomics__EVAL_33),
    ._EVAL_34(atomics__EVAL_34),
    ._EVAL_35(atomics__EVAL_35),
    ._EVAL_36(atomics__EVAL_36),
    ._EVAL_37(atomics__EVAL_37),
    ._EVAL_38(atomics__EVAL_38),
    ._EVAL_39(atomics__EVAL_39),
    ._EVAL_40(atomics__EVAL_40),
    ._EVAL_41(atomics__EVAL_41),
    ._EVAL_42(atomics__EVAL_42),
    ._EVAL_43(atomics__EVAL_43),
    ._EVAL_44(atomics__EVAL_44),
    ._EVAL_45(atomics__EVAL_45),
    ._EVAL_46(atomics__EVAL_46),
    ._EVAL_47(atomics__EVAL_47),
    ._EVAL_48(atomics__EVAL_48)
  );
  _EVAL_67 coupler_to_clint (
    ._EVAL(coupler_to_clint__EVAL),
    ._EVAL_0(coupler_to_clint__EVAL_0),
    ._EVAL_1(coupler_to_clint__EVAL_1),
    ._EVAL_2(coupler_to_clint__EVAL_2),
    ._EVAL_3(coupler_to_clint__EVAL_3),
    ._EVAL_4(coupler_to_clint__EVAL_4),
    ._EVAL_5(coupler_to_clint__EVAL_5),
    ._EVAL_6(coupler_to_clint__EVAL_6),
    ._EVAL_7(coupler_to_clint__EVAL_7),
    ._EVAL_8(coupler_to_clint__EVAL_8),
    ._EVAL_9(coupler_to_clint__EVAL_9),
    ._EVAL_10(coupler_to_clint__EVAL_10),
    ._EVAL_11(coupler_to_clint__EVAL_11),
    ._EVAL_12(coupler_to_clint__EVAL_12),
    ._EVAL_13(coupler_to_clint__EVAL_13),
    ._EVAL_14(coupler_to_clint__EVAL_14),
    ._EVAL_15(coupler_to_clint__EVAL_15),
    ._EVAL_16(coupler_to_clint__EVAL_16),
    ._EVAL_17(coupler_to_clint__EVAL_17),
    ._EVAL_18(coupler_to_clint__EVAL_18),
    ._EVAL_19(coupler_to_clint__EVAL_19),
    ._EVAL_20(coupler_to_clint__EVAL_20),
    ._EVAL_21(coupler_to_clint__EVAL_21),
    ._EVAL_22(coupler_to_clint__EVAL_22),
    ._EVAL_23(coupler_to_clint__EVAL_23),
    ._EVAL_24(coupler_to_clint__EVAL_24),
    ._EVAL_25(coupler_to_clint__EVAL_25),
    ._EVAL_26(coupler_to_clint__EVAL_26),
    ._EVAL_27(coupler_to_clint__EVAL_27),
    ._EVAL_28(coupler_to_clint__EVAL_28),
    ._EVAL_29(coupler_to_clint__EVAL_29),
    ._EVAL_30(coupler_to_clint__EVAL_30),
    ._EVAL_31(coupler_to_clint__EVAL_31),
    ._EVAL_32(coupler_to_clint__EVAL_32)
  );
  _EVAL_59 wrapped_error_device (
    ._EVAL(wrapped_error_device__EVAL),
    ._EVAL_0(wrapped_error_device__EVAL_0),
    ._EVAL_1(wrapped_error_device__EVAL_1),
    ._EVAL_2(wrapped_error_device__EVAL_2),
    ._EVAL_3(wrapped_error_device__EVAL_3),
    ._EVAL_4(wrapped_error_device__EVAL_4),
    ._EVAL_5(wrapped_error_device__EVAL_5),
    ._EVAL_6(wrapped_error_device__EVAL_6),
    ._EVAL_7(wrapped_error_device__EVAL_7),
    ._EVAL_8(wrapped_error_device__EVAL_8),
    ._EVAL_9(wrapped_error_device__EVAL_9),
    ._EVAL_10(wrapped_error_device__EVAL_10),
    ._EVAL_11(wrapped_error_device__EVAL_11),
    ._EVAL_12(wrapped_error_device__EVAL_12),
    ._EVAL_13(wrapped_error_device__EVAL_13),
    ._EVAL_14(wrapped_error_device__EVAL_14),
    ._EVAL_15(wrapped_error_device__EVAL_15),
    ._EVAL_16(wrapped_error_device__EVAL_16),
    ._EVAL_17(wrapped_error_device__EVAL_17),
    ._EVAL_18(wrapped_error_device__EVAL_18),
    ._EVAL_19(wrapped_error_device__EVAL_19)
  );
  _EVAL_77 coupler_to_tile (
    ._EVAL(coupler_to_tile__EVAL),
    ._EVAL_0(coupler_to_tile__EVAL_0),
    ._EVAL_1(coupler_to_tile__EVAL_1),
    ._EVAL_2(coupler_to_tile__EVAL_2),
    ._EVAL_3(coupler_to_tile__EVAL_3),
    ._EVAL_4(coupler_to_tile__EVAL_4),
    ._EVAL_5(coupler_to_tile__EVAL_5),
    ._EVAL_6(coupler_to_tile__EVAL_6),
    ._EVAL_7(coupler_to_tile__EVAL_7),
    ._EVAL_8(coupler_to_tile__EVAL_8),
    ._EVAL_9(coupler_to_tile__EVAL_9),
    ._EVAL_10(coupler_to_tile__EVAL_10),
    ._EVAL_11(coupler_to_tile__EVAL_11),
    ._EVAL_12(coupler_to_tile__EVAL_12),
    ._EVAL_13(coupler_to_tile__EVAL_13),
    ._EVAL_14(coupler_to_tile__EVAL_14),
    ._EVAL_15(coupler_to_tile__EVAL_15),
    ._EVAL_16(coupler_to_tile__EVAL_16),
    ._EVAL_17(coupler_to_tile__EVAL_17),
    ._EVAL_18(coupler_to_tile__EVAL_18),
    ._EVAL_19(coupler_to_tile__EVAL_19),
    ._EVAL_20(coupler_to_tile__EVAL_20),
    ._EVAL_21(coupler_to_tile__EVAL_21),
    ._EVAL_22(coupler_to_tile__EVAL_22),
    ._EVAL_23(coupler_to_tile__EVAL_23),
    ._EVAL_24(coupler_to_tile__EVAL_24),
    ._EVAL_25(coupler_to_tile__EVAL_25),
    ._EVAL_26(coupler_to_tile__EVAL_26),
    ._EVAL_27(coupler_to_tile__EVAL_27),
    ._EVAL_28(coupler_to_tile__EVAL_28),
    ._EVAL_29(coupler_to_tile__EVAL_29),
    ._EVAL_30(coupler_to_tile__EVAL_30),
    ._EVAL_31(coupler_to_tile__EVAL_31),
    ._EVAL_32(coupler_to_tile__EVAL_32),
    ._EVAL_33(coupler_to_tile__EVAL_33),
    ._EVAL_34(coupler_to_tile__EVAL_34),
    ._EVAL_35(coupler_to_tile__EVAL_35),
    ._EVAL_36(coupler_to_tile__EVAL_36),
    ._EVAL_37(coupler_to_tile__EVAL_37),
    ._EVAL_38(coupler_to_tile__EVAL_38),
    ._EVAL_39(coupler_to_tile__EVAL_39),
    ._EVAL_40(coupler_to_tile__EVAL_40),
    ._EVAL_41(coupler_to_tile__EVAL_41),
    ._EVAL_42(coupler_to_tile__EVAL_42),
    ._EVAL_43(coupler_to_tile__EVAL_43),
    ._EVAL_44(coupler_to_tile__EVAL_44),
    ._EVAL_45(coupler_to_tile__EVAL_45)
  );
  _EVAL_50 buffer (
    ._EVAL(buffer__EVAL),
    ._EVAL_0(buffer__EVAL_0),
    ._EVAL_1(buffer__EVAL_1),
    ._EVAL_2(buffer__EVAL_2),
    ._EVAL_3(buffer__EVAL_3),
    ._EVAL_4(buffer__EVAL_4),
    ._EVAL_5(buffer__EVAL_5),
    ._EVAL_6(buffer__EVAL_6),
    ._EVAL_7(buffer__EVAL_7),
    ._EVAL_8(buffer__EVAL_8),
    ._EVAL_9(buffer__EVAL_9),
    ._EVAL_10(buffer__EVAL_10),
    ._EVAL_11(buffer__EVAL_11),
    ._EVAL_12(buffer__EVAL_12),
    ._EVAL_13(buffer__EVAL_13),
    ._EVAL_14(buffer__EVAL_14),
    ._EVAL_15(buffer__EVAL_15),
    ._EVAL_16(buffer__EVAL_16),
    ._EVAL_17(buffer__EVAL_17),
    ._EVAL_18(buffer__EVAL_18),
    ._EVAL_19(buffer__EVAL_19),
    ._EVAL_20(buffer__EVAL_20),
    ._EVAL_21(buffer__EVAL_21),
    ._EVAL_22(buffer__EVAL_22),
    ._EVAL_23(buffer__EVAL_23),
    ._EVAL_24(buffer__EVAL_24),
    ._EVAL_25(buffer__EVAL_25),
    ._EVAL_26(buffer__EVAL_26),
    ._EVAL_27(buffer__EVAL_27),
    ._EVAL_28(buffer__EVAL_28),
    ._EVAL_29(buffer__EVAL_29),
    ._EVAL_30(buffer__EVAL_30),
    ._EVAL_31(buffer__EVAL_31),
    ._EVAL_32(buffer__EVAL_32),
    ._EVAL_33(buffer__EVAL_33),
    ._EVAL_34(buffer__EVAL_34),
    ._EVAL_35(buffer__EVAL_35),
    ._EVAL_36(buffer__EVAL_36),
    ._EVAL_37(buffer__EVAL_37),
    ._EVAL_38(buffer__EVAL_38),
    ._EVAL_39(buffer__EVAL_39),
    ._EVAL_40(buffer__EVAL_40),
    ._EVAL_41(buffer__EVAL_41),
    ._EVAL_42(buffer__EVAL_42),
    ._EVAL_43(buffer__EVAL_43),
    ._EVAL_44(buffer__EVAL_44),
    ._EVAL_45(buffer__EVAL_45),
    ._EVAL_46(buffer__EVAL_46),
    ._EVAL_47(buffer__EVAL_47),
    ._EVAL_48(buffer__EVAL_48)
  );
  _EVAL_46 out_xbar (
    ._EVAL(out_xbar__EVAL),
    ._EVAL_0(out_xbar__EVAL_0),
    ._EVAL_1(out_xbar__EVAL_1),
    ._EVAL_2(out_xbar__EVAL_2),
    ._EVAL_3(out_xbar__EVAL_3),
    ._EVAL_4(out_xbar__EVAL_4),
    ._EVAL_5(out_xbar__EVAL_5),
    ._EVAL_6(out_xbar__EVAL_6),
    ._EVAL_7(out_xbar__EVAL_7),
    ._EVAL_8(out_xbar__EVAL_8),
    ._EVAL_9(out_xbar__EVAL_9),
    ._EVAL_10(out_xbar__EVAL_10),
    ._EVAL_11(out_xbar__EVAL_11),
    ._EVAL_12(out_xbar__EVAL_12),
    ._EVAL_13(out_xbar__EVAL_13),
    ._EVAL_14(out_xbar__EVAL_14),
    ._EVAL_15(out_xbar__EVAL_15),
    ._EVAL_16(out_xbar__EVAL_16),
    ._EVAL_17(out_xbar__EVAL_17),
    ._EVAL_18(out_xbar__EVAL_18),
    ._EVAL_19(out_xbar__EVAL_19),
    ._EVAL_20(out_xbar__EVAL_20),
    ._EVAL_21(out_xbar__EVAL_21),
    ._EVAL_22(out_xbar__EVAL_22),
    ._EVAL_23(out_xbar__EVAL_23),
    ._EVAL_24(out_xbar__EVAL_24),
    ._EVAL_25(out_xbar__EVAL_25),
    ._EVAL_26(out_xbar__EVAL_26),
    ._EVAL_27(out_xbar__EVAL_27),
    ._EVAL_28(out_xbar__EVAL_28),
    ._EVAL_29(out_xbar__EVAL_29),
    ._EVAL_30(out_xbar__EVAL_30),
    ._EVAL_31(out_xbar__EVAL_31),
    ._EVAL_32(out_xbar__EVAL_32),
    ._EVAL_33(out_xbar__EVAL_33),
    ._EVAL_34(out_xbar__EVAL_34),
    ._EVAL_35(out_xbar__EVAL_35),
    ._EVAL_36(out_xbar__EVAL_36),
    ._EVAL_37(out_xbar__EVAL_37),
    ._EVAL_38(out_xbar__EVAL_38),
    ._EVAL_39(out_xbar__EVAL_39),
    ._EVAL_40(out_xbar__EVAL_40),
    ._EVAL_41(out_xbar__EVAL_41),
    ._EVAL_42(out_xbar__EVAL_42),
    ._EVAL_43(out_xbar__EVAL_43),
    ._EVAL_44(out_xbar__EVAL_44),
    ._EVAL_45(out_xbar__EVAL_45),
    ._EVAL_46(out_xbar__EVAL_46),
    ._EVAL_47(out_xbar__EVAL_47),
    ._EVAL_48(out_xbar__EVAL_48),
    ._EVAL_49(out_xbar__EVAL_49),
    ._EVAL_50(out_xbar__EVAL_50),
    ._EVAL_51(out_xbar__EVAL_51),
    ._EVAL_52(out_xbar__EVAL_52),
    ._EVAL_53(out_xbar__EVAL_53),
    ._EVAL_54(out_xbar__EVAL_54),
    ._EVAL_55(out_xbar__EVAL_55),
    ._EVAL_56(out_xbar__EVAL_56),
    ._EVAL_57(out_xbar__EVAL_57),
    ._EVAL_58(out_xbar__EVAL_58),
    ._EVAL_59(out_xbar__EVAL_59),
    ._EVAL_60(out_xbar__EVAL_60),
    ._EVAL_61(out_xbar__EVAL_61),
    ._EVAL_62(out_xbar__EVAL_62),
    ._EVAL_63(out_xbar__EVAL_63),
    ._EVAL_64(out_xbar__EVAL_64),
    ._EVAL_65(out_xbar__EVAL_65),
    ._EVAL_66(out_xbar__EVAL_66),
    ._EVAL_67(out_xbar__EVAL_67),
    ._EVAL_68(out_xbar__EVAL_68),
    ._EVAL_69(out_xbar__EVAL_69),
    ._EVAL_70(out_xbar__EVAL_70),
    ._EVAL_71(out_xbar__EVAL_71),
    ._EVAL_72(out_xbar__EVAL_72),
    ._EVAL_73(out_xbar__EVAL_73),
    ._EVAL_74(out_xbar__EVAL_74),
    ._EVAL_75(out_xbar__EVAL_75),
    ._EVAL_76(out_xbar__EVAL_76),
    ._EVAL_77(out_xbar__EVAL_77),
    ._EVAL_78(out_xbar__EVAL_78),
    ._EVAL_79(out_xbar__EVAL_79),
    ._EVAL_80(out_xbar__EVAL_80),
    ._EVAL_81(out_xbar__EVAL_81),
    ._EVAL_82(out_xbar__EVAL_82),
    ._EVAL_83(out_xbar__EVAL_83),
    ._EVAL_84(out_xbar__EVAL_84),
    ._EVAL_85(out_xbar__EVAL_85),
    ._EVAL_86(out_xbar__EVAL_86),
    ._EVAL_87(out_xbar__EVAL_87),
    ._EVAL_88(out_xbar__EVAL_88),
    ._EVAL_89(out_xbar__EVAL_89),
    ._EVAL_90(out_xbar__EVAL_90),
    ._EVAL_91(out_xbar__EVAL_91),
    ._EVAL_92(out_xbar__EVAL_92),
    ._EVAL_93(out_xbar__EVAL_93),
    ._EVAL_94(out_xbar__EVAL_94),
    ._EVAL_95(out_xbar__EVAL_95),
    ._EVAL_96(out_xbar__EVAL_96),
    ._EVAL_97(out_xbar__EVAL_97),
    ._EVAL_98(out_xbar__EVAL_98),
    ._EVAL_99(out_xbar__EVAL_99),
    ._EVAL_100(out_xbar__EVAL_100),
    ._EVAL_101(out_xbar__EVAL_101),
    ._EVAL_102(out_xbar__EVAL_102),
    ._EVAL_103(out_xbar__EVAL_103),
    ._EVAL_104(out_xbar__EVAL_104),
    ._EVAL_105(out_xbar__EVAL_105),
    ._EVAL_106(out_xbar__EVAL_106),
    ._EVAL_107(out_xbar__EVAL_107),
    ._EVAL_108(out_xbar__EVAL_108),
    ._EVAL_109(out_xbar__EVAL_109),
    ._EVAL_110(out_xbar__EVAL_110),
    ._EVAL_111(out_xbar__EVAL_111),
    ._EVAL_112(out_xbar__EVAL_112),
    ._EVAL_113(out_xbar__EVAL_113),
    ._EVAL_114(out_xbar__EVAL_114),
    ._EVAL_115(out_xbar__EVAL_115),
    ._EVAL_116(out_xbar__EVAL_116),
    ._EVAL_117(out_xbar__EVAL_117),
    ._EVAL_118(out_xbar__EVAL_118),
    ._EVAL_119(out_xbar__EVAL_119),
    ._EVAL_120(out_xbar__EVAL_120),
    ._EVAL_121(out_xbar__EVAL_121),
    ._EVAL_122(out_xbar__EVAL_122),
    ._EVAL_123(out_xbar__EVAL_123),
    ._EVAL_124(out_xbar__EVAL_124),
    ._EVAL_125(out_xbar__EVAL_125),
    ._EVAL_126(out_xbar__EVAL_126),
    ._EVAL_127(out_xbar__EVAL_127),
    ._EVAL_128(out_xbar__EVAL_128),
    ._EVAL_129(out_xbar__EVAL_129),
    ._EVAL_130(out_xbar__EVAL_130),
    ._EVAL_131(out_xbar__EVAL_131),
    ._EVAL_132(out_xbar__EVAL_132),
    ._EVAL_133(out_xbar__EVAL_133),
    ._EVAL_134(out_xbar__EVAL_134),
    ._EVAL_135(out_xbar__EVAL_135),
    ._EVAL_136(out_xbar__EVAL_136),
    ._EVAL_137(out_xbar__EVAL_137),
    ._EVAL_138(out_xbar__EVAL_138),
    ._EVAL_139(out_xbar__EVAL_139),
    ._EVAL_140(out_xbar__EVAL_140),
    ._EVAL_141(out_xbar__EVAL_141),
    ._EVAL_142(out_xbar__EVAL_142),
    ._EVAL_143(out_xbar__EVAL_143),
    ._EVAL_144(out_xbar__EVAL_144),
    ._EVAL_145(out_xbar__EVAL_145),
    ._EVAL_146(out_xbar__EVAL_146)
  );
  _EVAL_71 coupler_to_debug (
    ._EVAL(coupler_to_debug__EVAL),
    ._EVAL_0(coupler_to_debug__EVAL_0),
    ._EVAL_1(coupler_to_debug__EVAL_1),
    ._EVAL_2(coupler_to_debug__EVAL_2),
    ._EVAL_3(coupler_to_debug__EVAL_3),
    ._EVAL_4(coupler_to_debug__EVAL_4),
    ._EVAL_5(coupler_to_debug__EVAL_5),
    ._EVAL_6(coupler_to_debug__EVAL_6),
    ._EVAL_7(coupler_to_debug__EVAL_7),
    ._EVAL_8(coupler_to_debug__EVAL_8),
    ._EVAL_9(coupler_to_debug__EVAL_9),
    ._EVAL_10(coupler_to_debug__EVAL_10),
    ._EVAL_11(coupler_to_debug__EVAL_11),
    ._EVAL_12(coupler_to_debug__EVAL_12),
    ._EVAL_13(coupler_to_debug__EVAL_13),
    ._EVAL_14(coupler_to_debug__EVAL_14),
    ._EVAL_15(coupler_to_debug__EVAL_15),
    ._EVAL_16(coupler_to_debug__EVAL_16),
    ._EVAL_17(coupler_to_debug__EVAL_17),
    ._EVAL_18(coupler_to_debug__EVAL_18),
    ._EVAL_19(coupler_to_debug__EVAL_19),
    ._EVAL_20(coupler_to_debug__EVAL_20),
    ._EVAL_21(coupler_to_debug__EVAL_21),
    ._EVAL_22(coupler_to_debug__EVAL_22),
    ._EVAL_23(coupler_to_debug__EVAL_23),
    ._EVAL_24(coupler_to_debug__EVAL_24),
    ._EVAL_25(coupler_to_debug__EVAL_25),
    ._EVAL_26(coupler_to_debug__EVAL_26),
    ._EVAL_27(coupler_to_debug__EVAL_27),
    ._EVAL_28(coupler_to_debug__EVAL_28),
    ._EVAL_29(coupler_to_debug__EVAL_29),
    ._EVAL_30(coupler_to_debug__EVAL_30),
    ._EVAL_31(coupler_to_debug__EVAL_31),
    ._EVAL_32(coupler_to_debug__EVAL_32)
  );
  _EVAL_42 fixedClockNode (
    ._EVAL(fixedClockNode__EVAL),
    ._EVAL_0(fixedClockNode__EVAL_0),
    ._EVAL_1(fixedClockNode__EVAL_1),
    ._EVAL_2(fixedClockNode__EVAL_2),
    ._EVAL_3(fixedClockNode__EVAL_3),
    ._EVAL_4(fixedClockNode__EVAL_4),
    ._EVAL_5(fixedClockNode__EVAL_5),
    ._EVAL_6(fixedClockNode__EVAL_6)
  );
  _EVAL_89 coupler_to_port_named_ahb_periph_port (
    ._EVAL(coupler_to_port_named_ahb_periph_port__EVAL),
    ._EVAL_0(coupler_to_port_named_ahb_periph_port__EVAL_0),
    ._EVAL_1(coupler_to_port_named_ahb_periph_port__EVAL_1),
    ._EVAL_2(coupler_to_port_named_ahb_periph_port__EVAL_2),
    ._EVAL_3(coupler_to_port_named_ahb_periph_port__EVAL_3),
    ._EVAL_4(coupler_to_port_named_ahb_periph_port__EVAL_4),
    ._EVAL_5(coupler_to_port_named_ahb_periph_port__EVAL_5),
    ._EVAL_6(coupler_to_port_named_ahb_periph_port__EVAL_6),
    ._EVAL_7(coupler_to_port_named_ahb_periph_port__EVAL_7),
    ._EVAL_8(coupler_to_port_named_ahb_periph_port__EVAL_8),
    ._EVAL_9(coupler_to_port_named_ahb_periph_port__EVAL_9),
    ._EVAL_10(coupler_to_port_named_ahb_periph_port__EVAL_10),
    ._EVAL_11(coupler_to_port_named_ahb_periph_port__EVAL_11),
    ._EVAL_12(coupler_to_port_named_ahb_periph_port__EVAL_12),
    ._EVAL_13(coupler_to_port_named_ahb_periph_port__EVAL_13),
    ._EVAL_14(coupler_to_port_named_ahb_periph_port__EVAL_14),
    ._EVAL_15(coupler_to_port_named_ahb_periph_port__EVAL_15),
    ._EVAL_16(coupler_to_port_named_ahb_periph_port__EVAL_16),
    ._EVAL_17(coupler_to_port_named_ahb_periph_port__EVAL_17),
    ._EVAL_18(coupler_to_port_named_ahb_periph_port__EVAL_18),
    ._EVAL_19(coupler_to_port_named_ahb_periph_port__EVAL_19),
    ._EVAL_20(coupler_to_port_named_ahb_periph_port__EVAL_20),
    ._EVAL_21(coupler_to_port_named_ahb_periph_port__EVAL_21),
    ._EVAL_22(coupler_to_port_named_ahb_periph_port__EVAL_22),
    ._EVAL_23(coupler_to_port_named_ahb_periph_port__EVAL_23),
    ._EVAL_24(coupler_to_port_named_ahb_periph_port__EVAL_24),
    ._EVAL_25(coupler_to_port_named_ahb_periph_port__EVAL_25),
    ._EVAL_26(coupler_to_port_named_ahb_periph_port__EVAL_26),
    ._EVAL_27(coupler_to_port_named_ahb_periph_port__EVAL_27),
    ._EVAL_28(coupler_to_port_named_ahb_periph_port__EVAL_28),
    ._EVAL_29(coupler_to_port_named_ahb_periph_port__EVAL_29),
    ._EVAL_30(coupler_to_port_named_ahb_periph_port__EVAL_30),
    ._EVAL_31(coupler_to_port_named_ahb_periph_port__EVAL_31),
    ._EVAL_32(coupler_to_port_named_ahb_periph_port__EVAL_32),
    ._EVAL_33(coupler_to_port_named_ahb_periph_port__EVAL_33)
  );
  _EVAL_44 fixer (
    ._EVAL(fixer__EVAL),
    ._EVAL_0(fixer__EVAL_0),
    ._EVAL_1(fixer__EVAL_1),
    ._EVAL_2(fixer__EVAL_2),
    ._EVAL_3(fixer__EVAL_3),
    ._EVAL_4(fixer__EVAL_4),
    ._EVAL_5(fixer__EVAL_5),
    ._EVAL_6(fixer__EVAL_6),
    ._EVAL_7(fixer__EVAL_7),
    ._EVAL_8(fixer__EVAL_8),
    ._EVAL_9(fixer__EVAL_9),
    ._EVAL_10(fixer__EVAL_10),
    ._EVAL_11(fixer__EVAL_11),
    ._EVAL_12(fixer__EVAL_12),
    ._EVAL_13(fixer__EVAL_13),
    ._EVAL_14(fixer__EVAL_14),
    ._EVAL_15(fixer__EVAL_15),
    ._EVAL_16(fixer__EVAL_16),
    ._EVAL_17(fixer__EVAL_17),
    ._EVAL_18(fixer__EVAL_18),
    ._EVAL_19(fixer__EVAL_19),
    ._EVAL_20(fixer__EVAL_20),
    ._EVAL_21(fixer__EVAL_21),
    ._EVAL_22(fixer__EVAL_22),
    ._EVAL_23(fixer__EVAL_23),
    ._EVAL_24(fixer__EVAL_24),
    ._EVAL_25(fixer__EVAL_25),
    ._EVAL_26(fixer__EVAL_26),
    ._EVAL_27(fixer__EVAL_27),
    ._EVAL_28(fixer__EVAL_28),
    ._EVAL_29(fixer__EVAL_29),
    ._EVAL_30(fixer__EVAL_30),
    ._EVAL_31(fixer__EVAL_31),
    ._EVAL_32(fixer__EVAL_32),
    ._EVAL_33(fixer__EVAL_33),
    ._EVAL_34(fixer__EVAL_34),
    ._EVAL_35(fixer__EVAL_35),
    ._EVAL_36(fixer__EVAL_36),
    ._EVAL_37(fixer__EVAL_37),
    ._EVAL_38(fixer__EVAL_38),
    ._EVAL_39(fixer__EVAL_39),
    ._EVAL_40(fixer__EVAL_40),
    ._EVAL_41(fixer__EVAL_41),
    ._EVAL_42(fixer__EVAL_42),
    ._EVAL_43(fixer__EVAL_43),
    ._EVAL_44(fixer__EVAL_44),
    ._EVAL_45(fixer__EVAL_45),
    ._EVAL_46(fixer__EVAL_46),
    ._EVAL_47(fixer__EVAL_47),
    ._EVAL_48(fixer__EVAL_48)
  );
  _EVAL_93 coupler_to_testIndicator (
    ._EVAL(coupler_to_testIndicator__EVAL),
    ._EVAL_0(coupler_to_testIndicator__EVAL_0),
    ._EVAL_1(coupler_to_testIndicator__EVAL_1),
    ._EVAL_2(coupler_to_testIndicator__EVAL_2),
    ._EVAL_3(coupler_to_testIndicator__EVAL_3),
    ._EVAL_4(coupler_to_testIndicator__EVAL_4),
    ._EVAL_5(coupler_to_testIndicator__EVAL_5),
    ._EVAL_6(coupler_to_testIndicator__EVAL_6),
    ._EVAL_7(coupler_to_testIndicator__EVAL_7),
    ._EVAL_8(coupler_to_testIndicator__EVAL_8),
    ._EVAL_9(coupler_to_testIndicator__EVAL_9),
    ._EVAL_10(coupler_to_testIndicator__EVAL_10),
    ._EVAL_11(coupler_to_testIndicator__EVAL_11),
    ._EVAL_12(coupler_to_testIndicator__EVAL_12),
    ._EVAL_13(coupler_to_testIndicator__EVAL_13),
    ._EVAL_14(coupler_to_testIndicator__EVAL_14),
    ._EVAL_15(coupler_to_testIndicator__EVAL_15),
    ._EVAL_16(coupler_to_testIndicator__EVAL_16),
    ._EVAL_17(coupler_to_testIndicator__EVAL_17),
    ._EVAL_18(coupler_to_testIndicator__EVAL_18),
    ._EVAL_19(coupler_to_testIndicator__EVAL_19),
    ._EVAL_20(coupler_to_testIndicator__EVAL_20),
    ._EVAL_21(coupler_to_testIndicator__EVAL_21),
    ._EVAL_22(coupler_to_testIndicator__EVAL_22),
    ._EVAL_23(coupler_to_testIndicator__EVAL_23),
    ._EVAL_24(coupler_to_testIndicator__EVAL_24),
    ._EVAL_25(coupler_to_testIndicator__EVAL_25),
    ._EVAL_26(coupler_to_testIndicator__EVAL_26),
    ._EVAL_27(coupler_to_testIndicator__EVAL_27),
    ._EVAL_28(coupler_to_testIndicator__EVAL_28),
    ._EVAL_29(coupler_to_testIndicator__EVAL_29),
    ._EVAL_30(coupler_to_testIndicator__EVAL_30),
    ._EVAL_31(coupler_to_testIndicator__EVAL_31),
    ._EVAL_32(coupler_to_testIndicator__EVAL_32)
  );
  _EVAL_63 coupler_to_plic (
    ._EVAL(coupler_to_plic__EVAL),
    ._EVAL_0(coupler_to_plic__EVAL_0),
    ._EVAL_1(coupler_to_plic__EVAL_1),
    ._EVAL_2(coupler_to_plic__EVAL_2),
    ._EVAL_3(coupler_to_plic__EVAL_3),
    ._EVAL_4(coupler_to_plic__EVAL_4),
    ._EVAL_5(coupler_to_plic__EVAL_5),
    ._EVAL_6(coupler_to_plic__EVAL_6),
    ._EVAL_7(coupler_to_plic__EVAL_7),
    ._EVAL_8(coupler_to_plic__EVAL_8),
    ._EVAL_9(coupler_to_plic__EVAL_9),
    ._EVAL_10(coupler_to_plic__EVAL_10),
    ._EVAL_11(coupler_to_plic__EVAL_11),
    ._EVAL_12(coupler_to_plic__EVAL_12),
    ._EVAL_13(coupler_to_plic__EVAL_13),
    ._EVAL_14(coupler_to_plic__EVAL_14),
    ._EVAL_15(coupler_to_plic__EVAL_15),
    ._EVAL_16(coupler_to_plic__EVAL_16),
    ._EVAL_17(coupler_to_plic__EVAL_17),
    ._EVAL_18(coupler_to_plic__EVAL_18),
    ._EVAL_19(coupler_to_plic__EVAL_19),
    ._EVAL_20(coupler_to_plic__EVAL_20),
    ._EVAL_21(coupler_to_plic__EVAL_21),
    ._EVAL_22(coupler_to_plic__EVAL_22),
    ._EVAL_23(coupler_to_plic__EVAL_23),
    ._EVAL_24(coupler_to_plic__EVAL_24),
    ._EVAL_25(coupler_to_plic__EVAL_25),
    ._EVAL_26(coupler_to_plic__EVAL_26),
    ._EVAL_27(coupler_to_plic__EVAL_27),
    ._EVAL_28(coupler_to_plic__EVAL_28),
    ._EVAL_29(coupler_to_plic__EVAL_29),
    ._EVAL_30(coupler_to_plic__EVAL_30),
    ._EVAL_31(coupler_to_plic__EVAL_31),
    ._EVAL_32(coupler_to_plic__EVAL_32)
  );
  assign _EVAL_147 = _EVAL_61;
  assign atomics__EVAL_40 = buffer__EVAL_23;
  assign _EVAL_163 = _EVAL_225;
  assign buffer__EVAL_5 = atomics__EVAL_29;
  assign _EVAL_88 = coupler_to_plic__EVAL_5;
  assign buffer__EVAL_26 = fixedClockNode__EVAL;
  assign coupler_to_port_named_ahb_periph_port__EVAL_25 = fixedClockNode__EVAL;
  assign coupler_to_tile__EVAL_34 = _EVAL_107;
  assign _EVAL_86 = coupler_to_plic__EVAL_32;
  assign coupler_to_debug__EVAL_21 = out_xbar__EVAL_119;
  assign out_xbar__EVAL_104 = coupler_to_debug__EVAL_14;
  assign coupler_to_debug__EVAL_28 = out_xbar__EVAL_51;
  assign _EVAL_200 = _EVAL_212;
  assign _EVAL_21 = coupler_to_testIndicator__EVAL_17;
  assign _EVAL_190 = _EVAL_50;
  assign coupler_to_port_named_ahb_periph_port__EVAL_5 = out_xbar__EVAL_103;
  assign coupler_to_clint__EVAL_5 = _EVAL_11;
  assign _EVAL_48 = coupler_to_tile__EVAL_30;
  assign out_xbar__EVAL_14 = fixer__EVAL_17;
  assign _EVAL_25 = coupler_to_debug__EVAL_16;
  assign coupler_to_port_named_ahb_periph_port__EVAL_17 = out_xbar__EVAL_87;
  assign fixer__EVAL_9 = out_xbar__EVAL_2;
  assign _EVAL_29 = coupler_to_port_named_ahb_periph_port__EVAL_14;
  assign _EVAL_97 = coupler_to_tile__EVAL_15;
  assign atomics__EVAL_48 = _EVAL_146;
  assign atomics__EVAL_11 = buffer__EVAL_12;
  assign coupler_to_testIndicator__EVAL_20 = out_xbar__EVAL_11;
  assign out_xbar__EVAL_130 = wrapped_error_device__EVAL_3;
  assign _EVAL_130 = coupler_to_tile__EVAL_42;
  assign out_xbar__EVAL_17 = coupler_to_tile__EVAL_28;
  assign out_xbar__EVAL_113 = fixer__EVAL_33;
  assign coupler_to_tile__EVAL_41 = _EVAL_98;
  assign _EVAL_8 = coupler_to_debug__EVAL_20;
  assign coupler_to_debug__EVAL_9 = out_xbar__EVAL_140;
  assign out_xbar__EVAL_77 = coupler_to_clint__EVAL_14;
  assign coupler_to_debug__EVAL_12 = _EVAL_128;
  assign buffer__EVAL_25 = atomics__EVAL_42;
  assign coupler_to_tile__EVAL_21 = fixedClockNode__EVAL;
  assign out_xbar__EVAL_22 = fixedClockNode__EVAL;
  assign coupler_to_port_named_ahb_periph_port__EVAL_27 = _EVAL_15;
  assign _EVAL_132 = fixedClockNode__EVAL_4;
  assign _EVAL_222 = _EVAL_229;
  assign _EVAL_182 = _EVAL_140;
  assign atomics__EVAL_6 = buffer__EVAL_42;
  assign coupler_to_tile__EVAL_3 = _EVAL_5;
  assign _EVAL_127 = coupler_to_port_named_ahb_periph_port__EVAL_3;
  assign coupler_to_tile__EVAL_26 = _EVAL_27;
  assign _EVAL_207 = _EVAL_152;
  assign coupler_to_port_named_ahb_periph_port__EVAL_12 = _EVAL_68;
  assign coupler_to_port_named_ahb_periph_port__EVAL_9 = out_xbar__EVAL_109;
  assign out_xbar__EVAL_19 = fixer__EVAL_43;
  assign wrapped_error_device__EVAL_1 = out_xbar__EVAL_126;
  assign _EVAL_227 = _EVAL_237;
  assign _EVAL_169 = _EVAL_150;
  assign out_xbar__EVAL_141 = coupler_to_tile__EVAL_10;
  assign _EVAL_183 = _EVAL_177;
  assign _EVAL_87 = coupler_to_tile__EVAL_39;
  assign coupler_to_tile__EVAL_45 = _EVAL_63;
  assign atomics__EVAL_45 = _EVAL_231;
  assign fixer__EVAL_21 = out_xbar__EVAL_144;
  assign _EVAL_92 = coupler_to_clint__EVAL_16;
  assign _EVAL_72 = _EVAL_235;
  assign atomics__EVAL_25 = buffer__EVAL_33;
  assign _EVAL = coupler_to_debug__EVAL_10;
  assign out_xbar__EVAL_146 = coupler_to_port_named_ahb_periph_port__EVAL_26;
  assign _EVAL_179 = _EVAL_227;
  assign _EVAL_194 = _EVAL_224;
  assign coupler_to_debug__EVAL_0 = _EVAL_67;
  assign _EVAL_129 = coupler_to_clint__EVAL_9;
  assign _EVAL_140 = _EVAL_169;
  assign coupler_to_tile__EVAL_5 = _EVAL_94;
  assign _EVAL_148 = _EVAL_223;
  assign _EVAL_196 = _EVAL_183;
  assign _EVAL_198 = atomics__EVAL_43;
  assign atomics__EVAL_31 = buffer__EVAL_16;
  assign _EVAL_22 = coupler_to_clint__EVAL_27;
  assign _EVAL_79 = coupler_to_tile__EVAL_25;
  assign _EVAL_154 = _EVAL_142;
  assign coupler_to_tile__EVAL_18 = out_xbar__EVAL_34;
  assign fixer__EVAL_25 = out_xbar__EVAL_0;
  assign coupler_to_port_named_ahb_periph_port__EVAL_8 = out_xbar__EVAL_47;
  assign _EVAL_230 = _EVAL_181;
  assign out_xbar__EVAL_23 = fixer__EVAL_41;
  assign buffer__EVAL_15 = fixer__EVAL_14;
  assign out_xbar__EVAL = wrapped_error_device__EVAL_13;
  assign buffer__EVAL_0 = atomics__EVAL_17;
  assign fixer__EVAL_29 = buffer__EVAL;
  assign out_xbar__EVAL_125 = coupler_to_debug__EVAL_4;
  assign _EVAL_121 = coupler_to_tile__EVAL_22;
  assign _EVAL_112 = coupler_to_testIndicator__EVAL_32;
  assign atomics__EVAL_2 = _EVAL_217;
  assign out_xbar__EVAL_33 = fixer__EVAL_22;
  assign _EVAL_167 = atomics__EVAL_39;
  assign out_xbar__EVAL_29 = coupler_to_clint__EVAL_15;
  assign _EVAL_2 = coupler_to_tile__EVAL_7;
  assign out_xbar__EVAL_37 = coupler_to_tile__EVAL_17;
  assign fixer__EVAL_48 = out_xbar__EVAL_54;
  assign fixer__EVAL_16 = buffer__EVAL_21;
  assign _EVAL_170 = _EVAL_173;
  assign _EVAL_236 = _EVAL_233;
  assign _EVAL_125 = coupler_to_plic__EVAL_2;
  assign coupler_to_port_named_ahb_periph_port__EVAL_30 = out_xbar__EVAL_85;
  assign coupler_to_debug__EVAL_15 = fixedClockNode__EVAL;
  assign _EVAL_152 = _EVAL_168;
  assign _EVAL_157 = _EVAL_164;
  assign _EVAL_141 = _EVAL_195;
  assign _EVAL_39 = coupler_to_debug__EVAL_5;
  assign coupler_to_clint__EVAL_24 = _EVAL_62;
  assign out_xbar__EVAL_128 = wrapped_error_device__EVAL_12;
  assign coupler_to_port_named_ahb_periph_port__EVAL = out_xbar__EVAL_31;
  assign wrapped_error_device__EVAL_19 = fixedClockNode__EVAL_6;
  assign coupler_to_plic__EVAL_9 = out_xbar__EVAL_62;
  assign fixer__EVAL_38 = out_xbar__EVAL_28;
  assign fixer__EVAL_36 = buffer__EVAL_31;
  assign fixer__EVAL_27 = out_xbar__EVAL_110;
  assign _EVAL_138 = _EVAL_141;
  assign _EVAL_136 = _EVAL_207;
  assign _EVAL_199 = _EVAL_197;
  assign atomics__EVAL_8 = fixedClockNode__EVAL;
  assign coupler_to_testIndicator__EVAL_6 = fixedClockNode__EVAL;
  assign _EVAL_31 = coupler_to_tile__EVAL_29;
  assign fixedClockNode__EVAL_3 = _EVAL_215;
  assign fixer__EVAL_35 = buffer__EVAL_35;
  assign coupler_to_testIndicator__EVAL_19 = out_xbar__EVAL_6;
  assign _EVAL_171 = _EVAL_176;
  assign _EVAL_1 = coupler_to_tile__EVAL_27;
  assign _EVAL_150 = _EVAL_42;
  assign coupler_to_clint__EVAL_18 = out_xbar__EVAL_117;
  assign _EVAL_166 = _EVAL_153;
  assign coupler_to_testIndicator__EVAL_18 = out_xbar__EVAL_122;
  assign wrapped_error_device__EVAL_10 = out_xbar__EVAL_95;
  assign out_xbar__EVAL_107 = coupler_to_clint__EVAL;
  assign atomics__EVAL_35 = buffer__EVAL_1;
  assign _EVAL_137 = _EVAL_219;
  assign out_xbar__EVAL_78 = coupler_to_debug__EVAL_11;
  assign _EVAL_93 = coupler_to_debug__EVAL_19;
  assign _EVAL_57 = coupler_to_tile__EVAL_14;
  assign _EVAL_7 = coupler_to_plic__EVAL_12;
  assign buffer__EVAL_32 = atomics__EVAL_15;
  assign fixer__EVAL_12 = fixedClockNode__EVAL;
  assign coupler_to_tile__EVAL = _EVAL_83;
  assign _EVAL_185 = _EVAL_144;
  assign out_xbar__EVAL_53 = fixer__EVAL_24;
  assign _EVAL_193 = _EVAL_184;
  assign coupler_to_tile__EVAL_9 = out_xbar__EVAL_50;
  assign _EVAL_233 = _EVAL_193;
  assign _EVAL_158 = _EVAL_170;
  assign coupler_to_port_named_ahb_periph_port__EVAL_20 = fixedClockNode__EVAL_6;
  assign out_xbar__EVAL_74 = coupler_to_testIndicator__EVAL_10;
  assign coupler_to_clint__EVAL_20 = out_xbar__EVAL_90;
  assign coupler_to_plic__EVAL_0 = _EVAL_123;
  assign coupler_to_plic__EVAL_16 = _EVAL_70;
  assign atomics__EVAL_33 = _EVAL_149;
  assign out_xbar__EVAL_82 = wrapped_error_device__EVAL_5;
  assign coupler_to_clint__EVAL_11 = out_xbar__EVAL_57;
  assign out_xbar__EVAL_65 = coupler_to_plic__EVAL_19;
  assign coupler_to_testIndicator__EVAL_21 = out_xbar__EVAL_92;
  assign _EVAL_232 = _EVAL_199;
  assign out_xbar__EVAL_118 = coupler_to_debug__EVAL_2;
  assign coupler_to_tile__EVAL_12 = _EVAL_28;
  assign out_xbar__EVAL_36 = wrapped_error_device__EVAL_8;
  assign _EVAL_174 = _EVAL_155;
  assign _EVAL_224 = _EVAL_216;
  assign fixer__EVAL_15 = buffer__EVAL_9;
  assign out_xbar__EVAL_127 = coupler_to_testIndicator__EVAL_13;
  assign coupler_to_debug__EVAL_22 = out_xbar__EVAL_120;
  assign coupler_to_plic__EVAL = out_xbar__EVAL_3;
  assign buffer__EVAL_18 = atomics__EVAL_19;
  assign coupler_to_port_named_ahb_periph_port__EVAL_19 = out_xbar__EVAL_67;
  assign atomics__EVAL_16 = _EVAL_221;
  assign out_xbar__EVAL_143 = coupler_to_plic__EVAL_29;
  assign out_xbar__EVAL_16 = coupler_to_port_named_ahb_periph_port__EVAL_13;
  assign fixer__EVAL_19 = buffer__EVAL_8;
  assign _EVAL_115 = _EVAL_172;
  assign coupler_to_clint__EVAL_26 = out_xbar__EVAL_18;
  assign _EVAL_204 = _EVAL_122;
  assign coupler_to_tile__EVAL_13 = out_xbar__EVAL_137;
  assign coupler_to_port_named_ahb_periph_port__EVAL_22 = out_xbar__EVAL_114;
  assign coupler_to_clint__EVAL_13 = _EVAL_16;
  assign _EVAL_153 = _EVAL_230;
  assign buffer__EVAL_46 = fixer__EVAL_31;
  assign _EVAL_109 = _EVAL_191;
  assign atomics__EVAL_44 = fixedClockNode__EVAL_6;
  assign buffer__EVAL_36 = fixer__EVAL_28;
  assign coupler_to_clint__EVAL_10 = fixedClockNode__EVAL;
  assign coupler_to_testIndicator__EVAL_4 = out_xbar__EVAL_58;
  assign atomics__EVAL_12 = _EVAL_182;
  assign atomics__EVAL_9 = _EVAL_166;
  assign buffer__EVAL_22 = fixedClockNode__EVAL_6;
  assign wrapped_error_device__EVAL_11 = out_xbar__EVAL_25;
  assign _EVAL_181 = _EVAL_36;
  assign _EVAL_210 = _EVAL_185;
  assign _EVAL_221 = _EVAL_175;
  assign buffer__EVAL_11 = fixer__EVAL_32;
  assign coupler_to_port_named_ahb_periph_port__EVAL_7 = out_xbar__EVAL_66;
  assign coupler_to_plic__EVAL_24 = out_xbar__EVAL_55;
  assign coupler_to_testIndicator__EVAL_28 = _EVAL_114;
  assign out_xbar__EVAL_9 = coupler_to_clint__EVAL_25;
  assign _EVAL_12 = coupler_to_testIndicator__EVAL_22;
  assign _EVAL_176 = _EVAL_160;
  assign out_xbar__EVAL_44 = fixer__EVAL_39;
  assign fixer__EVAL_3 = out_xbar__EVAL_70;
  assign coupler_to_plic__EVAL_8 = _EVAL_32;
  assign _EVAL_64 = coupler_to_testIndicator__EVAL;
  assign out_xbar__EVAL_97 = coupler_to_plic__EVAL_21;
  assign _EVAL_6 = coupler_to_debug__EVAL_3;
  assign out_xbar__EVAL_35 = coupler_to_clint__EVAL_21;
  assign coupler_to_tile__EVAL_20 = out_xbar__EVAL_139;
  assign out_xbar__EVAL_24 = coupler_to_debug__EVAL_26;
  assign _EVAL_225 = atomics__EVAL_23;
  assign fixer__EVAL_20 = buffer__EVAL_7;
  assign out_xbar__EVAL_84 = fixer__EVAL_34;
  assign buffer__EVAL_6 = fixer__EVAL_5;
  assign coupler_to_tile__EVAL_38 = out_xbar__EVAL_136;
  assign coupler_to_clint__EVAL_19 = _EVAL_126;
  assign _EVAL_144 = _EVAL_76;
  assign _EVAL_33 = coupler_to_debug__EVAL_6;
  assign coupler_to_testIndicator__EVAL_0 = out_xbar__EVAL_134;
  assign fixer__EVAL_1 = out_xbar__EVAL_1;
  assign out_xbar__EVAL_111 = coupler_to_tile__EVAL_6;
  assign coupler_to_plic__EVAL_15 = out_xbar__EVAL_115;
  assign _EVAL_223 = _EVAL_26;
  assign _EVAL_195 = atomics__EVAL_20;
  assign coupler_to_debug__EVAL_25 = out_xbar__EVAL_21;
  assign _EVAL_124 = coupler_to_clint__EVAL_6;
  assign coupler_to_port_named_ahb_periph_port__EVAL_18 = out_xbar__EVAL_26;
  assign _EVAL_162 = _EVAL_158;
  assign out_xbar__EVAL_38 = coupler_to_port_named_ahb_periph_port__EVAL_29;
  assign _EVAL_187 = _EVAL_192;
  assign coupler_to_tile__EVAL_4 = _EVAL_24;
  assign coupler_to_port_named_ahb_periph_port__EVAL_32 = out_xbar__EVAL_121;
  assign coupler_to_testIndicator__EVAL_24 = out_xbar__EVAL_145;
  assign _EVAL_117 = coupler_to_plic__EVAL_11;
  assign coupler_to_debug__EVAL_29 = _EVAL_19;
  assign coupler_to_testIndicator__EVAL_23 = _EVAL_120;
  assign _EVAL_202 = atomics__EVAL_37;
  assign atomics__EVAL_4 = _EVAL_179;
  assign coupler_to_debug__EVAL_32 = _EVAL_118;
  assign _EVAL_237 = _EVAL_211;
  assign coupler_to_port_named_ahb_periph_port__EVAL_4 = out_xbar__EVAL_142;
  assign _EVAL_108 = coupler_to_tile__EVAL_40;
  assign coupler_to_plic__EVAL_23 = out_xbar__EVAL_60;
  assign coupler_to_tile__EVAL_31 = out_xbar__EVAL_80;
  assign _EVAL_215 = _EVAL_194;
  assign buffer__EVAL_30 = atomics__EVAL_10;
  assign buffer__EVAL_28 = fixer__EVAL_46;
  assign _EVAL_226 = _EVAL_174;
  assign _EVAL_20 = coupler_to_clint__EVAL_22;
  assign _EVAL_131 = coupler_to_testIndicator__EVAL_26;
  assign out_xbar__EVAL_75 = coupler_to_testIndicator__EVAL_11;
  assign coupler_to_plic__EVAL_30 = out_xbar__EVAL_124;
  assign out_xbar__EVAL_102 = coupler_to_plic__EVAL_13;
  assign atomics__EVAL_28 = buffer__EVAL_14;
  assign _EVAL_155 = _EVAL_188;
  assign _EVAL_84 = _EVAL_226;
  assign _EVAL_191 = _EVAL_214;
  assign _EVAL_160 = _EVAL_165;
  assign coupler_to_plic__EVAL_7 = out_xbar__EVAL_101;
  assign _EVAL_228 = _EVAL_198;
  assign fixer__EVAL_40 = out_xbar__EVAL_52;
  assign _EVAL_159 = _EVAL_75;
  assign _EVAL_65 = _EVAL_205;
  assign buffer__EVAL_4 = atomics__EVAL_1;
  assign _EVAL_145 = _EVAL_190;
  assign _EVAL_89 = _EVAL_171;
  assign out_xbar__EVAL_105 = wrapped_error_device__EVAL_6;
  assign fixer__EVAL_44 = buffer__EVAL_43;
  assign out_xbar__EVAL_81 = coupler_to_testIndicator__EVAL_14;
  assign _EVAL_103 = coupler_to_plic__EVAL_3;
  assign coupler_to_port_named_ahb_periph_port__EVAL_11 = out_xbar__EVAL_30;
  assign wrapped_error_device__EVAL_7 = out_xbar__EVAL_93;
  assign _EVAL_205 = _EVAL_208;
  assign _EVAL_186 = _EVAL_138;
  assign coupler_to_clint__EVAL_31 = out_xbar__EVAL_42;
  assign out_xbar__EVAL_76 = coupler_to_port_named_ahb_periph_port__EVAL_33;
  assign _EVAL_69 = coupler_to_tile__EVAL_44;
  assign _EVAL_111 = coupler_to_testIndicator__EVAL_30;
  assign _EVAL_161 = _EVAL_209;
  assign buffer__EVAL_48 = fixer__EVAL_2;
  assign _EVAL_91 = coupler_to_plic__EVAL_1;
  assign _EVAL_208 = _EVAL_228;
  assign _EVAL_77 = coupler_to_clint__EVAL_30;
  assign wrapped_error_device__EVAL_4 = out_xbar__EVAL_63;
  assign coupler_to_tile__EVAL_33 = out_xbar__EVAL_59;
  assign _EVAL_105 = coupler_to_port_named_ahb_periph_port__EVAL_2;
  assign atomics__EVAL_18 = buffer__EVAL_34;
  assign _EVAL_231 = _EVAL_206;
  assign fixer__EVAL_8 = buffer__EVAL_29;
  assign coupler_to_clint__EVAL_4 = out_xbar__EVAL_116;
  assign coupler_to_testIndicator__EVAL_16 = out_xbar__EVAL_40;
  assign _EVAL_173 = _EVAL_35;
  assign coupler_to_debug__EVAL_7 = _EVAL_40;
  assign out_xbar__EVAL_10 = wrapped_error_device__EVAL_15;
  assign _EVAL_201 = _EVAL_55;
  assign _EVAL_73 = coupler_to_tile__EVAL_1;
  assign _EVAL_53 = coupler_to_plic__EVAL_10;
  assign buffer__EVAL_27 = atomics__EVAL_22;
  assign _EVAL_203 = _EVAL_200;
  assign _EVAL_229 = _EVAL_189;
  assign _EVAL_45 = coupler_to_testIndicator__EVAL_12;
  assign coupler_to_clint__EVAL_28 = fixedClockNode__EVAL_6;
  assign _EVAL_218 = _EVAL_145;
  assign atomics__EVAL_27 = _EVAL_180;
  assign coupler_to_tile__EVAL_19 = _EVAL_34;
  assign out_xbar__EVAL_72 = coupler_to_plic__EVAL_25;
  assign _EVAL_135 = _EVAL_85;
  assign buffer__EVAL_47 = atomics__EVAL_41;
  assign buffer__EVAL_45 = atomics__EVAL_30;
  assign _EVAL_178 = _EVAL_159;
  assign _EVAL_156 = _EVAL_202;
  assign coupler_to_tile__EVAL_23 = out_xbar__EVAL_138;
  assign _EVAL_38 = _EVAL_154;
  assign coupler_to_port_named_ahb_periph_port__EVAL_21 = out_xbar__EVAL_129;
  assign coupler_to_port_named_ahb_periph_port__EVAL_23 = _EVAL_82;
  assign out_xbar__EVAL_45 = coupler_to_debug__EVAL_1;
  assign _EVAL_209 = _EVAL_135;
  assign out_xbar__EVAL_112 = fixer__EVAL_18;
  assign _EVAL_146 = _EVAL_210;
  assign _EVAL_110 = coupler_to_tile__EVAL_37;
  assign _EVAL_43 = _EVAL_186;
  assign out_xbar__EVAL_132 = wrapped_error_device__EVAL;
  assign _EVAL_3 = _EVAL_236;
  assign atomics__EVAL_0 = _EVAL_157;
  assign atomics__EVAL_5 = buffer__EVAL_17;
  assign atomics__EVAL_24 = buffer__EVAL_2;
  assign out_xbar__EVAL_135 = fixer__EVAL_42;
  assign coupler_to_testIndicator__EVAL_1 = out_xbar__EVAL_64;
  assign coupler_to_clint__EVAL_29 = _EVAL_74;
  assign _EVAL_189 = _EVAL_113;
  assign fixer__EVAL_10 = buffer__EVAL_20;
  assign coupler_to_debug__EVAL_30 = out_xbar__EVAL_49;
  assign coupler_to_testIndicator__EVAL_15 = out_xbar__EVAL_13;
  assign fixer__EVAL_13 = buffer__EVAL_39;
  assign wrapped_error_device__EVAL_14 = fixedClockNode__EVAL;
  assign coupler_to_tile__EVAL_2 = _EVAL_96;
  assign out_xbar__EVAL_15 = coupler_to_port_named_ahb_periph_port__EVAL_15;
  assign _EVAL_37 = coupler_to_tile__EVAL_8;
  assign _EVAL_142 = _EVAL_213;
  assign _EVAL_234 = _EVAL_167;
  assign coupler_to_clint__EVAL_1 = out_xbar__EVAL_8;
  assign out_xbar__EVAL_5 = coupler_to_clint__EVAL_17;
  assign _EVAL_214 = _EVAL_234;
  assign coupler_to_tile__EVAL_35 = fixedClockNode__EVAL_6;
  assign _EVAL_52 = coupler_to_tile__EVAL_11;
  assign _EVAL_17 = fixedClockNode__EVAL_6;
  assign _EVAL_180 = _EVAL_187;
  assign _EVAL_95 = fixedClockNode__EVAL_5;
  assign coupler_to_clint__EVAL_23 = _EVAL_4;
  assign coupler_to_plic__EVAL_22 = _EVAL_9;
  assign _EVAL_46 = fixedClockNode__EVAL_0;
  assign _EVAL_100 = coupler_to_tile__EVAL_0;
  assign coupler_to_plic__EVAL_26 = out_xbar__EVAL_73;
  assign coupler_to_debug__EVAL_17 = out_xbar__EVAL_61;
  assign coupler_to_tile__EVAL_43 = _EVAL_23;
  assign _EVAL_81 = coupler_to_plic__EVAL_6;
  assign coupler_to_clint__EVAL_12 = out_xbar__EVAL_91;
  assign _EVAL_175 = _EVAL_178;
  assign wrapped_error_device__EVAL_9 = out_xbar__EVAL_94;
  assign _EVAL_164 = _EVAL_139;
  assign atomics__EVAL_34 = _EVAL_162;
  assign _EVAL_168 = _EVAL_80;
  assign _EVAL_54 = coupler_to_plic__EVAL_14;
  assign coupler_to_debug__EVAL_8 = _EVAL_104;
  assign coupler_to_plic__EVAL_17 = _EVAL_30;
  assign _EVAL_101 = coupler_to_tile__EVAL_32;
  assign _EVAL_172 = _EVAL_220;
  assign out_xbar__EVAL_71 = coupler_to_port_named_ahb_periph_port__EVAL_1;
  assign out_xbar__EVAL_68 = fixedClockNode__EVAL_6;
  assign buffer__EVAL_41 = atomics__EVAL_38;
  assign wrapped_error_device__EVAL_18 = out_xbar__EVAL_98;
  assign _EVAL_188 = atomics__EVAL_32;
  assign atomics__EVAL_26 = _EVAL_136;
  assign coupler_to_plic__EVAL_31 = fixedClockNode__EVAL_6;
  assign _EVAL_0 = coupler_to_testIndicator__EVAL_3;
  assign buffer__EVAL_37 = fixer__EVAL_6;
  assign coupler_to_debug__EVAL_27 = out_xbar__EVAL_4;
  assign out_xbar__EVAL_32 = coupler_to_port_named_ahb_periph_port__EVAL_16;
  assign _EVAL_134 = _EVAL_196;
  assign _EVAL_177 = _EVAL_49;
  assign buffer__EVAL_19 = atomics__EVAL;
  assign fixer__EVAL_37 = buffer__EVAL_44;
  assign coupler_to_tile__EVAL_24 = out_xbar__EVAL_43;
  assign fixer__EVAL_4 = fixedClockNode__EVAL_6;
  assign out_xbar__EVAL_86 = coupler_to_testIndicator__EVAL_8;
  assign _EVAL_14 = coupler_to_port_named_ahb_periph_port__EVAL_31;
  assign _EVAL_10 = coupler_to_testIndicator__EVAL_2;
  assign out_xbar__EVAL_123 = wrapped_error_device__EVAL_2;
  assign _EVAL_47 = coupler_to_testIndicator__EVAL_9;
  assign _EVAL_149 = _EVAL_222;
  assign atomics__EVAL_46 = _EVAL_232;
  assign _EVAL_151 = atomics__EVAL_13;
  assign _EVAL_44 = _EVAL_137;
  assign _EVAL_211 = _EVAL_56;
  assign _EVAL_41 = coupler_to_clint__EVAL_2;
  assign wrapped_error_device__EVAL_17 = out_xbar__EVAL_7;
  assign out_xbar__EVAL_48 = fixer__EVAL_45;
  assign coupler_to_testIndicator__EVAL_25 = _EVAL_51;
  assign _EVAL_184 = atomics__EVAL_21;
  assign _EVAL_58 = coupler_to_port_named_ahb_periph_port__EVAL_28;
  assign out_xbar__EVAL_100 = fixer__EVAL_7;
  assign _EVAL_99 = coupler_to_debug__EVAL_31;
  assign coupler_to_testIndicator__EVAL_29 = fixedClockNode__EVAL_6;
  assign _EVAL_197 = _EVAL_147;
  assign _EVAL_220 = _EVAL_163;
  assign atomics__EVAL_36 = _EVAL_134;
  assign _EVAL_212 = atomics__EVAL_3;
  assign coupler_to_testIndicator__EVAL_27 = _EVAL_119;
  assign out_xbar__EVAL_83 = fixer__EVAL_26;
  assign buffer__EVAL_3 = fixer__EVAL_23;
  assign out_xbar__EVAL_106 = coupler_to_testIndicator__EVAL_7;
  assign coupler_to_plic__EVAL_27 = _EVAL_59;
  assign out_xbar__EVAL_69 = coupler_to_port_named_ahb_periph_port__EVAL_0;
  assign fixer__EVAL_0 = buffer__EVAL_40;
  assign fixer__EVAL_47 = buffer__EVAL_38;
  assign fixedClockNode__EVAL_2 = _EVAL_143;
  assign coupler_to_plic__EVAL_20 = out_xbar__EVAL_12;
  assign coupler_to_debug__EVAL_24 = out_xbar__EVAL_39;
  assign _EVAL_13 = coupler_to_clint__EVAL_7;
  assign _EVAL_78 = coupler_to_debug__EVAL;
  assign coupler_to_plic__EVAL_4 = fixedClockNode__EVAL;
  assign _EVAL_71 = coupler_to_clint__EVAL_32;
  assign _EVAL_216 = _EVAL_133;
  assign coupler_to_clint__EVAL_3 = out_xbar__EVAL_133;
  assign fixer__EVAL_11 = out_xbar__EVAL_88;
  assign out_xbar__EVAL_89 = coupler_to_tile__EVAL_36;
  assign out_xbar__EVAL_96 = coupler_to_plic__EVAL_18;
  assign coupler_to_clint__EVAL_8 = out_xbar__EVAL_46;
  assign _EVAL_66 = fixedClockNode__EVAL_1;
  assign coupler_to_debug__EVAL_23 = fixedClockNode__EVAL_6;
  assign out_xbar__EVAL_41 = coupler_to_port_named_ahb_periph_port__EVAL_10;
  assign out_xbar__EVAL_20 = coupler_to_tile__EVAL_16;
  assign _EVAL_139 = _EVAL_204;
  assign out_xbar__EVAL_99 = coupler_to_port_named_ahb_periph_port__EVAL_6;
  assign coupler_to_plic__EVAL_28 = out_xbar__EVAL_27;
  assign coupler_to_testIndicator__EVAL_5 = _EVAL_18;
  assign buffer__EVAL_10 = fixer__EVAL;
  assign _EVAL_165 = atomics__EVAL_7;
  assign wrapped_error_device__EVAL_0 = out_xbar__EVAL_108;
  assign coupler_to_testIndicator__EVAL_31 = _EVAL_60;
  assign _EVAL_235 = _EVAL_203;
  assign _EVAL_106 = coupler_to_port_named_ahb_periph_port__EVAL_24;
  assign _EVAL_192 = _EVAL_201;
  assign _EVAL_213 = _EVAL_151;
  assign buffer__EVAL_24 = atomics__EVAL_47;
  assign _EVAL_206 = _EVAL_148;
  assign _EVAL_90 = coupler_to_clint__EVAL_0;
  assign out_xbar__EVAL_79 = fixer__EVAL_30;
  assign _EVAL_143 = _EVAL_218;
  assign coupler_to_debug__EVAL_18 = out_xbar__EVAL_56;
  assign _EVAL_116 = coupler_to_debug__EVAL_13;
  assign out_xbar__EVAL_131 = wrapped_error_device__EVAL_16;
  assign buffer__EVAL_13 = atomics__EVAL_14;
  assign _EVAL_219 = _EVAL_156;
  assign _EVAL_217 = _EVAL_161;
  assign _EVAL_102 = fixedClockNode__EVAL;
endmodule
