//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_147(
  input   _EVAL,
  output  _EVAL_0,
  input   _EVAL_1,
  input   _EVAL_2,
  input   _EVAL_3,
  output  _EVAL_4,
  output  _EVAL_5,
  output  _EVAL_6,
  input   _EVAL_7,
  output  _EVAL_8,
  output  _EVAL_9,
  input   _EVAL_10,
  output  _EVAL_11,
  input   _EVAL_12,
  output  _EVAL_13,
  input   _EVAL_14,
  input   _EVAL_15,
  input   _EVAL_16,
  output  _EVAL_17,
  output  _EVAL_18,
  output  _EVAL_19,
  output  _EVAL_20,
  input   _EVAL_21,
  input   _EVAL_22,
  input   _EVAL_23,
  input   _EVAL_24,
  output  _EVAL_25,
  output  _EVAL_26,
  input   _EVAL_27,
  output  _EVAL_28,
  input   _EVAL_29,
  output  _EVAL_30
);
  assign _EVAL_17 = _EVAL_21;
  assign _EVAL_0 = _EVAL;
  assign _EVAL_28 = _EVAL_12;
  assign _EVAL_9 = _EVAL_10;
  assign _EVAL_25 = _EVAL_1;
  assign _EVAL_19 = _EVAL_16;
  assign _EVAL_18 = _EVAL_22;
  assign _EVAL_13 = _EVAL_24;
  assign _EVAL_26 = _EVAL_23;
  assign _EVAL_11 = _EVAL_14;
  assign _EVAL_30 = _EVAL_29;
  assign _EVAL_6 = _EVAL_2;
  assign _EVAL_4 = _EVAL_7;
  assign _EVAL_5 = _EVAL_15;
  assign _EVAL_8 = _EVAL_3;
  assign _EVAL_20 = _EVAL_27;
endmodule
