//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_105_assert(
  input        _EVAL_2,
  input        _EVAL_3,
  input        _EVAL_4,
  input        _EVAL_6,
  input  [1:0] _EVAL_7,
  input        _EVAL_8,
  input  [1:0] _EVAL_10,
  input  [1:0] _EVAL_11,
  input  [1:0] _EVAL_12,
  input        _EVAL_13,
  input        _EVAL_14,
  input        _EVAL_15,
  input  [1:0] _EVAL_16,
  input        _EVAL_17,
  input        _EVAL_18,
  input        _EVAL_19,
  input        _EVAL_21,
  input        _EVAL_22,
  input        _EVAL_23,
  input        _EVAL_25,
  input        _EVAL_26,
  input        _EVAL_30,
  input  [1:0] _EVAL_31,
  input  [1:0] _EVAL_32,
  input        _EVAL_35,
  input        _EVAL_36,
  input        _EVAL_37,
  input  [1:0] _EVAL_40,
  input        _EVAL_43,
  input        _EVAL_44,
  input        _EVAL_48,
  input        _EVAL_49,
  input        _EVAL_50,
  input        _EVAL_51,
  input        _EVAL_52,
  input        _EVAL_55,
  input        _EVAL_56,
  input        _EVAL_57,
  input        _EVAL_58,
  input        _EVAL_59,
  input        _EVAL_60,
  input        _EVAL_61,
  input        _EVAL_84,
  input        _EVAL_113,
  input        _EVAL_119,
  input        _EVAL_125,
  input        _EVAL_159,
  input        _EVAL_173,
  input        _EVAL_181,
  input        _EVAL_204,
  input        _EVAL_248,
  input        _EVAL_254,
  input        _EVAL_285,
  input        _EVAL_308,
  input        _EVAL_328,
  input        _EVAL_332,
  input        _EVAL_378,
  input        _EVAL_396
);
  wire [2:0] _EVAL_62;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_69;
  wire  _EVAL_71;
  wire  _EVAL_73;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_87;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_101;
  wire [2:0] _EVAL_102;
  wire  _EVAL_104;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_112;
  wire  _EVAL_114;
  wire  _EVAL_118;
  wire  _EVAL_121;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_126;
  wire  _EVAL_129;
  wire  _EVAL_131;
  wire  _EVAL_133;
  wire  _EVAL_136;
  wire  _EVAL_138;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_149;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_170;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_178;
  wire  _EVAL_180;
  wire  _EVAL_184;
  wire  _EVAL_186;
  wire  _EVAL_194;
  wire [2:0] _EVAL_195;
  wire  _EVAL_197;
  wire [2:0] _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_206;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire [2:0] _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_222;
  wire [2:0] _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_232;
  wire [2:0] _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_243;
  wire  _EVAL_245;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_252;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_260;
  wire  _EVAL_262;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_273;
  wire  _EVAL_276;
  wire  _EVAL_278;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_284;
  wire  _EVAL_293;
  wire  _EVAL_295;
  wire  _EVAL_296;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_304;
  wire  _EVAL_307;
  wire  _EVAL_309;
  wire  _EVAL_310;
  wire  _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_326;
  wire  _EVAL_329;
  wire  _EVAL_333;
  wire  _EVAL_335;
  wire  _EVAL_337;
  wire  _EVAL_338;
  wire  _EVAL_339;
  wire  _EVAL_340;
  wire  _EVAL_341;
  wire  _EVAL_342;
  wire  _EVAL_343;
  wire  _EVAL_346;
  wire  _EVAL_347;
  wire  _EVAL_349;
  wire  _EVAL_350;
  wire  _EVAL_351;
  wire  _EVAL_352;
  wire  _EVAL_353;
  wire  _EVAL_355;
  wire  _EVAL_356;
  wire  _EVAL_358;
  wire  _EVAL_359;
  wire  _EVAL_360;
  wire [2:0] _EVAL_362;
  wire  _EVAL_363;
  wire  _EVAL_365;
  wire  _EVAL_368;
  wire  _EVAL_369;
  wire  _EVAL_371;
  wire  _EVAL_372;
  wire  _EVAL_373;
  wire  _EVAL_375;
  wire  _EVAL_380;
  wire  _EVAL_382;
  wire  _EVAL_383;
  wire  _EVAL_384;
  wire  _EVAL_385;
  wire  _EVAL_387;
  wire  _EVAL_388;
  wire  _EVAL_390;
  wire  _EVAL_391;
  wire  _EVAL_393;
  wire  _EVAL_394;
  wire  _EVAL_395;
  wire  _EVAL_398;
  wire  _EVAL_399;
  wire  _EVAL_402;
  assign _EVAL_402 = _EVAL_212 & _EVAL_95;
  assign _EVAL_81 = _EVAL_210 & _EVAL_311;
  assign _EVAL_342 = _EVAL_180 & _EVAL_109;
  assign _EVAL_238 = _EVAL_219 == 3'h4;
  assign _EVAL_71 = _EVAL_129 & _EVAL_351;
  assign _EVAL_309 = _EVAL_102 == 3'h1;
  assign _EVAL_382 = _EVAL_107 & _EVAL_313;
  assign _EVAL_149 = _EVAL_11 == 2'h3;
  assign _EVAL_206 = _EVAL_102 == 3'h4;
  assign _EVAL_92 = _EVAL_350 & _EVAL_174;
  assign _EVAL_213 = _EVAL_12 == 2'h3;
  assign _EVAL_359 = _EVAL_211 & _EVAL_394;
  assign _EVAL_312 = _EVAL_32 == 2'h3;
  assign _EVAL_262 = _EVAL_164 & _EVAL_371;
  assign _EVAL_398 = _EVAL_195 == 3'h7;
  assign _EVAL_101 = _EVAL_252 & _EVAL_175;
  assign _EVAL_310 = _EVAL_195 == 3'h4;
  assign _EVAL_346 = _EVAL_82 & _EVAL_75;
  assign _EVAL_375 = _EVAL_96 & _EVAL_213;
  assign _EVAL_250 = _EVAL_10 == 2'h3;
  assign _EVAL_102 = {_EVAL_8,_EVAL_44,_EVAL_3};
  assign _EVAL_82 = _EVAL_13 & _EVAL_181;
  assign _EVAL_339 = _EVAL_82 & _EVAL_149;
  assign _EVAL_164 = _EVAL_229 & _EVAL_254;
  assign _EVAL_216 = ~_EVAL_113;
  assign _EVAL_296 = _EVAL_107 & _EVAL_282;
  assign _EVAL_66 = _EVAL_164 & _EVAL_123;
  assign _EVAL_175 = _EVAL_7 == 2'h2;
  assign _EVAL_184 = _EVAL_362 == 3'h1;
  assign _EVAL_95 = _EVAL_12 == 2'h2;
  assign _EVAL_211 = _EVAL_220 & _EVAL_308;
  assign _EVAL_282 = _EVAL_31 == 2'h2;
  assign _EVAL_129 = _EVAL_319 & _EVAL_285;
  assign _EVAL_65 = _EVAL_199 == 3'h4;
  assign _EVAL_356 = _EVAL_258 & _EVAL_278;
  assign _EVAL_106 = _EVAL_131 & _EVAL_125;
  assign _EVAL_110 = _EVAL_195 == 3'h5;
  assign _EVAL_69 = _EVAL_82 & _EVAL_109;
  assign _EVAL_307 = _EVAL_62 == 3'h4;
  assign _EVAL_112 = _EVAL_129 & _EVAL_175;
  assign _EVAL_299 = ~_EVAL_159;
  assign _EVAL_383 = _EVAL_7 == 2'h0;
  assign _EVAL_107 = _EVAL_35 & _EVAL_125;
  assign _EVAL_243 = _EVAL_96 & _EVAL_315;
  assign _EVAL_104 = _EVAL_12 == 2'h0;
  assign _EVAL_114 = _EVAL_224 == 3'h4;
  assign _EVAL_225 = _EVAL_212 & _EVAL_315;
  assign _EVAL_351 = _EVAL_7 == 2'h3;
  assign _EVAL_252 = _EVAL_2 & _EVAL_285;
  assign _EVAL_142 = _EVAL_195 == 3'h1;
  assign _EVAL_385 = _EVAL_258 & _EVAL_221;
  assign _EVAL_338 = _EVAL_362 == 3'h0;
  assign _EVAL_197 = _EVAL_102 == 3'h7;
  assign _EVAL_249 = _EVAL_62 == 3'h7;
  assign _EVAL_349 = _EVAL_199 == 3'h1;
  assign _EVAL_126 = _EVAL_245 & _EVAL_278;
  assign _EVAL_270 = _EVAL_252 & _EVAL_154;
  assign _EVAL_281 = _EVAL_31 == 2'h3;
  assign _EVAL_230 = _EVAL_62 == 3'h5;
  assign _EVAL_194 = _EVAL_362 == 3'h4;
  assign _EVAL_273 = _EVAL_210 & _EVAL_337;
  assign _EVAL_257 = _EVAL_102 == 3'h5;
  assign _EVAL_93 = ~_EVAL_84;
  assign _EVAL_123 = _EVAL_40 == 2'h1;
  assign _EVAL_75 = _EVAL_11 == 2'h2;
  assign _EVAL_368 = _EVAL_199 == 3'h0;
  assign _EVAL_237 = {_EVAL_22,_EVAL_59,_EVAL_25};
  assign _EVAL_217 = _EVAL_102 == 3'h3;
  assign _EVAL_315 = _EVAL_12 == 2'h1;
  assign _EVAL_300 = _EVAL_237 == 3'h1;
  assign _EVAL_91 = _EVAL_219 == 3'h7;
  assign _EVAL_109 = _EVAL_11 == 2'h1;
  assign _EVAL_141 = _EVAL_224 == 3'h3;
  assign _EVAL_393 = _EVAL_180 & _EVAL_149;
  assign _EVAL_77 = _EVAL_10 == 2'h0;
  assign _EVAL_365 = _EVAL_362 == 3'h7;
  assign _EVAL_224 = {_EVAL_49,_EVAL_4,_EVAL_14};
  assign _EVAL_118 = _EVAL_106 & _EVAL_281;
  assign _EVAL_284 = _EVAL_96 & _EVAL_95;
  assign _EVAL_220 = ~_EVAL_332;
  assign _EVAL_341 = _EVAL_199 == 3'h5;
  assign _EVAL_76 = _EVAL_326 & _EVAL_311;
  assign _EVAL_136 = _EVAL_252 & _EVAL_351;
  assign _EVAL_362 = {_EVAL_55,_EVAL_17,_EVAL_56};
  assign _EVAL_384 = _EVAL_62 == 3'h1;
  assign _EVAL_352 = _EVAL_164 & _EVAL_174;
  assign _EVAL_124 = _EVAL_40 == 2'h0;
  assign _EVAL_295 = _EVAL_16 == 2'h0;
  assign _EVAL_360 = _EVAL_245 & _EVAL_250;
  assign _EVAL_316 = _EVAL_237 == 3'h5;
  assign _EVAL_180 = _EVAL_93 & _EVAL_181;
  assign _EVAL_276 = _EVAL_224 == 3'h0;
  assign _EVAL_131 = ~_EVAL_248;
  assign _EVAL_200 = _EVAL_6 & _EVAL_308;
  assign _EVAL_319 = ~_EVAL_378;
  assign _EVAL_210 = _EVAL_61 & _EVAL_396;
  assign _EVAL_154 = _EVAL_7 == 2'h1;
  assign _EVAL_333 = _EVAL_31 == 2'h0;
  assign _EVAL_335 = _EVAL_326 & _EVAL_312;
  assign _EVAL_371 = _EVAL_40 == 2'h2;
  assign _EVAL_278 = _EVAL_10 == 2'h1;
  assign _EVAL_133 = _EVAL_350 & _EVAL_371;
  assign _EVAL_353 = _EVAL_200 & _EVAL_394;
  assign _EVAL_199 = {_EVAL_18,_EVAL_50,_EVAL_26};
  assign _EVAL_174 = _EVAL_40 == 2'h3;
  assign _EVAL_153 = _EVAL_16 == 2'h1;
  assign _EVAL_121 = _EVAL_237 == 3'h4;
  assign _EVAL_390 = _EVAL_212 & _EVAL_213;
  assign _EVAL_97 = _EVAL_219 == 3'h3;
  assign _EVAL_313 = _EVAL_31 == 2'h1;
  assign _EVAL_372 = _EVAL_106 & _EVAL_313;
  assign _EVAL_355 = _EVAL_237 == 3'h0;
  assign _EVAL_298 = _EVAL_219 == 3'h5;
  assign _EVAL_108 = _EVAL_195 == 3'h3;
  assign _EVAL_391 = _EVAL_224 == 3'h5;
  assign _EVAL_195 = {_EVAL_21,_EVAL_57,_EVAL_48};
  assign _EVAL_258 = _EVAL_216 & _EVAL_204;
  assign _EVAL_176 = _EVAL_106 & _EVAL_282;
  assign _EVAL_395 = _EVAL_245 & _EVAL_221;
  assign _EVAL_388 = _EVAL_219 == 3'h0;
  assign _EVAL_212 = _EVAL_232 & _EVAL_119;
  assign _EVAL_394 = _EVAL_16 == 2'h3;
  assign _EVAL_311 = _EVAL_32 == 2'h2;
  assign _EVAL_380 = _EVAL_107 & _EVAL_281;
  assign _EVAL_350 = _EVAL_43 & _EVAL_254;
  assign _EVAL_340 = _EVAL_180 & _EVAL_75;
  assign _EVAL_343 = _EVAL_11 == 2'h0;
  assign _EVAL_293 = _EVAL_200 & _EVAL_153;
  assign _EVAL_201 = _EVAL_200 & _EVAL_170;
  assign _EVAL_219 = {_EVAL_23,_EVAL_60,_EVAL_36};
  assign _EVAL_229 = ~_EVAL_173;
  assign _EVAL_170 = _EVAL_16 == 2'h2;
  assign _EVAL_245 = _EVAL_19 & _EVAL_204;
  assign _EVAL_163 = _EVAL_102 == 3'h0;
  assign _EVAL_326 = _EVAL_299 & _EVAL_396;
  assign _EVAL_73 = _EVAL_237 == 3'h3;
  assign _EVAL_165 = _EVAL_219 == 3'h1;
  assign _EVAL_96 = _EVAL_51 & _EVAL_119;
  assign _EVAL_186 = _EVAL_211 & _EVAL_153;
  assign _EVAL_363 = _EVAL_195 == 3'h0;
  assign _EVAL_222 = _EVAL_224 == 3'h7;
  assign _EVAL_269 = _EVAL_199 == 3'h3;
  assign _EVAL_301 = _EVAL_237 == 3'h7;
  assign _EVAL_369 = _EVAL_326 & _EVAL_337;
  assign _EVAL_232 = ~_EVAL_328;
  assign _EVAL_358 = _EVAL_199 == 3'h7;
  assign _EVAL_98 = _EVAL_32 == 2'h0;
  assign _EVAL_178 = _EVAL_224 == 3'h1;
  assign _EVAL_62 = {_EVAL_58,_EVAL_15,_EVAL_52};
  assign _EVAL_87 = ~_EVAL_30;
  assign _EVAL_347 = _EVAL_362 == 3'h5;
  assign _EVAL_337 = _EVAL_32 == 2'h1;
  assign _EVAL_221 = _EVAL_10 == 2'h2;
  assign _EVAL_260 = _EVAL_62 == 3'h0;
  assign _EVAL_399 = _EVAL_362 == 3'h3;
  assign _EVAL_138 = _EVAL_350 & _EVAL_123;
  assign _EVAL_387 = _EVAL_210 & _EVAL_312;
  assign _EVAL_373 = _EVAL_62 == 3'h3;
  assign _EVAL_329 = _EVAL_211 & _EVAL_170;
  assign _EVAL_318 = _EVAL_129 & _EVAL_154;
  assign _EVAL_304 = _EVAL_258 & _EVAL_250;
  always @(posedge _EVAL_37) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_35 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab4a2067)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_385 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d9af433)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b41c097f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_316 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80c29208)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd0e2c90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_225 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96848f20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e7c1114)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_346 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c81655b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab4a2067)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_335 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23110130)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_372 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96848f20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab4a2067)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_81 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c81655b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_77 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77daa290)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_13 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab4a2067)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_399 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc7fe073)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_384 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd0e2c90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_278 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d295b97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_353 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7219d3a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c81655b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_340 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d9af433)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23110130)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d9af433)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_186 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96848f20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_149 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b69b937d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e7c1114)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70b51b49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c81655b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_249 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7237de2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_153 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d295b97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_329 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d9af433)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_342 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96848f20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_298 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80c29208)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_398 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7237de2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_201 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c81655b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e7c1114)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b69b937d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_351 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b69b937d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_371 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b41c097f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7237de2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc7fe073)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_101 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c81655b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_394 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b69b937d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d295b97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_260 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a044c85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab4a2067)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_368 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a044c85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_184 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd0e2c90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_91 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7237de2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_250 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b69b937d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc7fe073)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_373 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc7fe073)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_310 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e7c1114)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c81655b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_390 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23110130)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_375 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7219d3a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80c29208)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80c29208)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_109 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d295b97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_391 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80c29208)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d9af433)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b69b937d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_356 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96848f20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_395 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c81655b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_276 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a044c85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_124 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77daa290)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_380 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7219d3a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_293 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70b51b49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_307 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e7c1114)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_349 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd0e2c90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7237de2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_341 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80c29208)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_337 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d295b97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_304 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23110130)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_355 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a044c85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_393 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23110130)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd0e2c90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_170 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b41c097f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_363 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a044c85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_388 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a044c85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_97 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc7fe073)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_318 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96848f20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77daa290)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_75 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b41c097f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_95 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b41c097f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_118 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23110130)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7219d3a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7237de2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_360 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7219d3a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80c29208)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7219d3a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_141 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc7fe073)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_243 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70b51b49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd0e2c90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e7c1114)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b41c097f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_382 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70b51b49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab4a2067)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_295 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77daa290)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd0e2c90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_206 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e7c1114)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70b51b49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_165 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd0e2c90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc7fe073)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_343 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77daa290)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_51 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab4a2067)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_312 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b69b937d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_359 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23110130)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_402 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d9af433)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_383 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77daa290)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab4a2067)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc7fe073)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_333 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77daa290)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_387 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7219d3a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70b51b49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_315 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d295b97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a044c85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e7c1114)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80c29208)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_358 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7237de2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7237de2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b41c097f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d295b97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_313 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d295b97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_369 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96848f20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_71 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(23110130)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_92 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7219d3a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_175 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b41c097f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77daa290)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96848f20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_338 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a044c85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_174 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b69b937d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_112 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d9af433)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_176 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d9af433)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_273 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70b51b49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_126 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70b51b49)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
