//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_22(
  output [3:0]  _EVAL,
  input  [1:0]  _EVAL_0,
  output        _EVAL_1,
  output [1:0]  _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  output        _EVAL_5,
  input         _EVAL_6,
  input  [3:0]  _EVAL_7,
  input  [3:0]  _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  output [31:0] _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input  [31:0] _EVAL_14,
  input  [3:0]  _EVAL_15,
  output [30:0] _EVAL_16,
  output [1:0]  _EVAL_17,
  input  [31:0] _EVAL_18,
  input         _EVAL_19,
  output        _EVAL_20,
  output [2:0]  _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23,
  input         _EVAL_24,
  output [31:0] _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  output [3:0]  _EVAL_28,
  input  [2:0]  _EVAL_29,
  output        _EVAL_30,
  input         _EVAL_31,
  output [1:0]  _EVAL_32,
  output        _EVAL_33,
  output        _EVAL_34,
  output        _EVAL_35,
  output        _EVAL_36,
  input  [31:0] _EVAL_37,
  output [1:0]  _EVAL_38,
  output [31:0] _EVAL_39,
  output        _EVAL_40,
  output [2:0]  _EVAL_41,
  output        _EVAL_42,
  output        _EVAL_43,
  input         _EVAL_44,
  input         _EVAL_45,
  output [1:0]  _EVAL_46,
  input  [31:0] _EVAL_47,
  output        _EVAL_48,
  input  [31:0] _EVAL_49,
  output [2:0]  _EVAL_50,
  input  [2:0]  _EVAL_51,
  input         _EVAL_52,
  output        _EVAL_53,
  input         _EVAL_54,
  input  [1:0]  _EVAL_55,
  output        _EVAL_56,
  output        _EVAL_57,
  input  [1:0]  _EVAL_58,
  output [2:0]  _EVAL_59,
  input  [3:0]  _EVAL_60,
  input         _EVAL_61,
  output [3:0]  _EVAL_62,
  input         _EVAL_63,
  input         _EVAL_64,
  output [2:0]  _EVAL_65,
  input         _EVAL_66,
  output        _EVAL_67,
  input  [4:0]  _EVAL_68,
  input         _EVAL_69,
  input         _EVAL_70,
  output        _EVAL_71,
  output        _EVAL_72,
  input  [2:0]  _EVAL_73,
  output [3:0]  _EVAL_74,
  output        _EVAL_75,
  input         _EVAL_76,
  output [2:0]  _EVAL_77,
  input  [2:0]  _EVAL_78,
  input  [31:0] _EVAL_79,
  output        _EVAL_80,
  input  [31:0] _EVAL_81,
  input  [3:0]  _EVAL_82,
  output [1:0]  _EVAL_83,
  output        _EVAL_84,
  output        _EVAL_85,
  output [31:0] _EVAL_86,
  input         _EVAL_87,
  input  [3:0]  _EVAL_88,
  output        _EVAL_89,
  input  [31:0] _EVAL_90,
  input         _EVAL_91,
  input  [3:0]  _EVAL_92,
  input  [2:0]  _EVAL_93,
  output [3:0]  _EVAL_94,
  output        _EVAL_95,
  input         _EVAL_96,
  output [3:0]  _EVAL_97,
  input  [3:0]  _EVAL_98,
  output [31:0] _EVAL_99,
  output        _EVAL_100,
  input  [2:0]  _EVAL_101,
  input         _EVAL_102,
  input         _EVAL_103,
  input         _EVAL_104,
  output        _EVAL_105,
  output        _EVAL_106,
  input         _EVAL_107,
  input  [2:0]  _EVAL_108,
  input  [3:0]  _EVAL_109,
  output [2:0]  _EVAL_110,
  input         _EVAL_111,
  output [3:0]  _EVAL_112,
  input         _EVAL_113,
  output [3:0]  _EVAL_114,
  output [4:0]  _EVAL_115,
  input         _EVAL_116,
  output [31:0] _EVAL_117,
  output        _EVAL_118
);
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire [31:0] _EVAL_123;
  wire  _EVAL_124;
  wire [2:0] _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire [3:0] _EVAL_130;
  wire [3:0] _EVAL_131;
  wire  _EVAL_132;
  wire  fixedClockNode__EVAL;
  wire  fixedClockNode__EVAL_0;
  wire  fixedClockNode__EVAL_1;
  wire  fixedClockNode__EVAL_2;
  wire [4:0] _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire [31:0] _EVAL_136;
  wire  _EVAL_137;
  wire [3:0] _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire [31:0] _EVAL_143;
  wire [3:0] _EVAL_144;
  wire [31:0] _EVAL_145;
  wire [2:0] _EVAL_146;
  wire  _EVAL_147;
  wire [2:0] _EVAL_148;
  wire  _EVAL_149;
  wire [1:0] _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire [31:0] coupler_from_tile__EVAL;
  wire  coupler_from_tile__EVAL_0;
  wire  coupler_from_tile__EVAL_1;
  wire [31:0] coupler_from_tile__EVAL_2;
  wire [3:0] coupler_from_tile__EVAL_3;
  wire [3:0] coupler_from_tile__EVAL_4;
  wire [31:0] coupler_from_tile__EVAL_5;
  wire [2:0] coupler_from_tile__EVAL_6;
  wire  coupler_from_tile__EVAL_7;
  wire  coupler_from_tile__EVAL_8;
  wire [31:0] coupler_from_tile__EVAL_9;
  wire [3:0] coupler_from_tile__EVAL_10;
  wire  coupler_from_tile__EVAL_11;
  wire [3:0] coupler_from_tile__EVAL_12;
  wire [2:0] coupler_from_tile__EVAL_13;
  wire  coupler_from_tile__EVAL_14;
  wire [31:0] coupler_from_tile__EVAL_15;
  wire [3:0] coupler_from_tile__EVAL_16;
  wire [2:0] coupler_from_tile__EVAL_17;
  wire  coupler_from_tile__EVAL_18;
  wire  coupler_from_tile__EVAL_19;
  wire [3:0] coupler_from_tile__EVAL_20;
  wire  coupler_from_tile__EVAL_21;
  wire [2:0] coupler_from_tile__EVAL_22;
  wire [3:0] coupler_from_tile__EVAL_23;
  wire [3:0] coupler_from_tile__EVAL_24;
  wire [2:0] coupler_from_tile__EVAL_25;
  wire  coupler_from_tile__EVAL_26;
  wire  coupler_from_tile__EVAL_27;
  wire [3:0] coupler_from_tile__EVAL_28;
  wire  coupler_from_tile__EVAL_29;
  wire  coupler_from_tile__EVAL_30;
  wire  coupler_from_tile__EVAL_31;
  wire [3:0] coupler_from_tile__EVAL_32;
  wire  coupler_from_tile__EVAL_33;
  wire [1:0] coupler_from_tile__EVAL_34;
  wire  coupler_from_tile__EVAL_35;
  wire [1:0] coupler_from_tile__EVAL_36;
  wire  coupler_from_tile__EVAL_37;
  wire [3:0] coupler_from_tile__EVAL_38;
  wire [1:0] coupler_from_tile__EVAL_39;
  wire [2:0] coupler_from_tile__EVAL_40;
  wire  coupler_from_tile__EVAL_41;
  wire  coupler_from_tile__EVAL_42;
  wire  coupler_from_tile__EVAL_43;
  wire [1:0] coupler_from_tile__EVAL_44;
  wire [31:0] coupler_from_tile__EVAL_45;
  wire  coupler_from_tile__EVAL_46;
  wire [2:0] coupler_from_tile__EVAL_47;
  wire  coupler_from_tile__EVAL_48;
  wire [2:0] coupler_from_tile__EVAL_49;
  wire [3:0] coupler_from_tile__EVAL_50;
  wire  coupler_from_tile__EVAL_51;
  wire [3:0] coupler_from_tile__EVAL_52;
  wire  coupler_from_tile__EVAL_53;
  wire  coupler_from_tile__EVAL_54;
  wire [1:0] coupler_from_tile__EVAL_55;
  wire [3:0] coupler_from_tile__EVAL_56;
  wire  coupler_from_tile__EVAL_57;
  wire  coupler_from_tile__EVAL_58;
  wire  coupler_from_tile__EVAL_59;
  wire [2:0] coupler_from_tile__EVAL_60;
  wire [31:0] coupler_from_tile__EVAL_61;
  wire [1:0] coupler_from_tile__EVAL_62;
  wire  coupler_from_tile__EVAL_63;
  wire  coupler_from_tile__EVAL_64;
  wire  coupler_from_tile__EVAL_65;
  wire  coupler_from_tile__EVAL_66;
  wire [31:0] coupler_from_tile__EVAL_67;
  wire [3:0] coupler_from_tile__EVAL_68;
  wire [31:0] coupler_from_tile__EVAL_69;
  wire [1:0] coupler_from_tile__EVAL_70;
  wire  coupler_from_tile__EVAL_71;
  wire  coupler_from_tile__EVAL_72;
  wire [3:0] _EVAL_155;
  wire  _EVAL_156;
  wire [31:0] _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire [31:0] _EVAL_163;
  wire [31:0] _EVAL_164;
  wire [3:0] _EVAL_165;
  wire [2:0] _EVAL_166;
  wire [4:0] _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire [4:0] _EVAL_170;
  wire [2:0] _EVAL_171;
  wire  _EVAL_172;
  wire [4:0] _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire [2:0] _EVAL_176;
  wire [1:0] _EVAL_177;
  wire [3:0] _EVAL_178;
  wire [3:0] _EVAL_179;
  wire [31:0] _EVAL_180;
  wire [3:0] _EVAL_181;
  wire [31:0] _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire [31:0] _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire [3:0] _EVAL_192;
  wire  _EVAL_193;
  wire [1:0] _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire [31:0] _EVAL_198;
  wire  system_bus_xbar__EVAL;
  wire  system_bus_xbar__EVAL_0;
  wire  system_bus_xbar__EVAL_1;
  wire [3:0] system_bus_xbar__EVAL_2;
  wire  system_bus_xbar__EVAL_3;
  wire [3:0] system_bus_xbar__EVAL_4;
  wire [3:0] system_bus_xbar__EVAL_5;
  wire [3:0] system_bus_xbar__EVAL_6;
  wire  system_bus_xbar__EVAL_7;
  wire [31:0] system_bus_xbar__EVAL_8;
  wire [2:0] system_bus_xbar__EVAL_9;
  wire  system_bus_xbar__EVAL_10;
  wire [2:0] system_bus_xbar__EVAL_11;
  wire  system_bus_xbar__EVAL_12;
  wire  system_bus_xbar__EVAL_13;
  wire  system_bus_xbar__EVAL_14;
  wire [2:0] system_bus_xbar__EVAL_15;
  wire [31:0] system_bus_xbar__EVAL_16;
  wire [31:0] system_bus_xbar__EVAL_17;
  wire [31:0] system_bus_xbar__EVAL_18;
  wire [2:0] system_bus_xbar__EVAL_19;
  wire [2:0] system_bus_xbar__EVAL_20;
  wire [1:0] system_bus_xbar__EVAL_21;
  wire  system_bus_xbar__EVAL_22;
  wire [31:0] system_bus_xbar__EVAL_23;
  wire  system_bus_xbar__EVAL_24;
  wire [31:0] system_bus_xbar__EVAL_25;
  wire  system_bus_xbar__EVAL_26;
  wire  system_bus_xbar__EVAL_27;
  wire  system_bus_xbar__EVAL_28;
  wire [3:0] system_bus_xbar__EVAL_29;
  wire  system_bus_xbar__EVAL_30;
  wire [1:0] system_bus_xbar__EVAL_31;
  wire  system_bus_xbar__EVAL_32;
  wire  system_bus_xbar__EVAL_33;
  wire  system_bus_xbar__EVAL_34;
  wire  system_bus_xbar__EVAL_35;
  wire  system_bus_xbar__EVAL_36;
  wire  system_bus_xbar__EVAL_37;
  wire [4:0] system_bus_xbar__EVAL_38;
  wire  system_bus_xbar__EVAL_39;
  wire [2:0] system_bus_xbar__EVAL_40;
  wire  system_bus_xbar__EVAL_41;
  wire  system_bus_xbar__EVAL_42;
  wire  system_bus_xbar__EVAL_43;
  wire  system_bus_xbar__EVAL_44;
  wire  system_bus_xbar__EVAL_45;
  wire  system_bus_xbar__EVAL_46;
  wire [30:0] system_bus_xbar__EVAL_47;
  wire  system_bus_xbar__EVAL_48;
  wire  system_bus_xbar__EVAL_49;
  wire [4:0] system_bus_xbar__EVAL_50;
  wire [2:0] system_bus_xbar__EVAL_51;
  wire [4:0] system_bus_xbar__EVAL_52;
  wire [31:0] system_bus_xbar__EVAL_53;
  wire [2:0] system_bus_xbar__EVAL_54;
  wire  system_bus_xbar__EVAL_55;
  wire [2:0] system_bus_xbar__EVAL_56;
  wire  system_bus_xbar__EVAL_57;
  wire [2:0] system_bus_xbar__EVAL_58;
  wire  system_bus_xbar__EVAL_59;
  wire [3:0] system_bus_xbar__EVAL_60;
  wire  system_bus_xbar__EVAL_61;
  wire  system_bus_xbar__EVAL_62;
  wire  system_bus_xbar__EVAL_63;
  wire  system_bus_xbar__EVAL_64;
  wire  system_bus_xbar__EVAL_65;
  wire [2:0] system_bus_xbar__EVAL_66;
  wire  system_bus_xbar__EVAL_67;
  wire  system_bus_xbar__EVAL_68;
  wire  system_bus_xbar__EVAL_69;
  wire [3:0] system_bus_xbar__EVAL_70;
  wire  system_bus_xbar__EVAL_71;
  wire  system_bus_xbar__EVAL_72;
  wire [1:0] system_bus_xbar__EVAL_73;
  wire  system_bus_xbar__EVAL_74;
  wire  system_bus_xbar__EVAL_75;
  wire [3:0] system_bus_xbar__EVAL_76;
  wire  system_bus_xbar__EVAL_77;
  wire [2:0] system_bus_xbar__EVAL_78;
  wire [31:0] system_bus_xbar__EVAL_79;
  wire [3:0] system_bus_xbar__EVAL_80;
  wire [2:0] system_bus_xbar__EVAL_81;
  wire [31:0] system_bus_xbar__EVAL_82;
  wire  system_bus_xbar__EVAL_83;
  wire [2:0] system_bus_xbar__EVAL_84;
  wire [3:0] system_bus_xbar__EVAL_85;
  wire  system_bus_xbar__EVAL_86;
  wire  system_bus_xbar__EVAL_87;
  wire [4:0] system_bus_xbar__EVAL_88;
  wire  system_bus_xbar__EVAL_89;
  wire  system_bus_xbar__EVAL_90;
  wire [3:0] system_bus_xbar__EVAL_91;
  wire [1:0] system_bus_xbar__EVAL_92;
  wire  system_bus_xbar__EVAL_93;
  wire [31:0] system_bus_xbar__EVAL_94;
  wire [3:0] system_bus_xbar__EVAL_95;
  wire [31:0] system_bus_xbar__EVAL_96;
  wire [2:0] _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire [31:0] _EVAL_203;
  wire [3:0] _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire [3:0] _EVAL_208;
  wire [2:0] _EVAL_209;
  wire [3:0] _EVAL_210;
  wire [31:0] fixer__EVAL;
  wire [2:0] fixer__EVAL_0;
  wire  fixer__EVAL_1;
  wire [31:0] fixer__EVAL_2;
  wire [3:0] fixer__EVAL_3;
  wire [2:0] fixer__EVAL_4;
  wire  fixer__EVAL_5;
  wire  fixer__EVAL_6;
  wire [1:0] fixer__EVAL_7;
  wire  fixer__EVAL_8;
  wire [3:0] fixer__EVAL_9;
  wire [1:0] fixer__EVAL_10;
  wire  fixer__EVAL_11;
  wire  fixer__EVAL_12;
  wire [3:0] fixer__EVAL_13;
  wire  fixer__EVAL_14;
  wire  fixer__EVAL_15;
  wire [2:0] fixer__EVAL_16;
  wire [31:0] fixer__EVAL_17;
  wire  fixer__EVAL_18;
  wire  fixer__EVAL_19;
  wire [3:0] fixer__EVAL_20;
  wire  fixer__EVAL_21;
  wire  fixer__EVAL_22;
  wire [31:0] fixer__EVAL_23;
  wire  fixer__EVAL_24;
  wire [2:0] fixer__EVAL_25;
  wire  fixer__EVAL_26;
  wire  fixer__EVAL_27;
  wire [2:0] fixer__EVAL_28;
  wire [3:0] fixer__EVAL_29;
  wire  fixer__EVAL_30;
  wire  fixer__EVAL_31;
  wire  fixer__EVAL_32;
  wire  fixer__EVAL_33;
  wire  fixer__EVAL_34;
  wire [31:0] fixer__EVAL_35;
  wire  fixer__EVAL_36;
  wire  fixer__EVAL_37;
  wire  fixer__EVAL_38;
  wire [3:0] fixer__EVAL_39;
  wire  fixer__EVAL_40;
  wire [3:0] fixer__EVAL_41;
  wire  fixer__EVAL_42;
  wire  fixer__EVAL_43;
  wire [3:0] fixer__EVAL_44;
  wire  fixer__EVAL_45;
  wire [31:0] fixer__EVAL_46;
  wire  fixer__EVAL_47;
  wire [31:0] fixer__EVAL_48;
  wire [3:0] fixer__EVAL_49;
  wire [3:0] fixer__EVAL_50;
  wire  fixer__EVAL_51;
  wire [31:0] fixer__EVAL_52;
  wire [1:0] fixer__EVAL_53;
  wire [2:0] fixer__EVAL_54;
  wire  fixer__EVAL_55;
  wire [2:0] fixer__EVAL_56;
  wire  fixer__EVAL_57;
  wire [2:0] fixer__EVAL_58;
  wire  fixer__EVAL_59;
  wire  fixer__EVAL_60;
  wire  fixer__EVAL_61;
  wire [2:0] fixer__EVAL_62;
  wire  fixer__EVAL_63;
  wire  fixer__EVAL_64;
  wire  fixer__EVAL_65;
  wire [1:0] fixer__EVAL_66;
  wire [3:0] fixer__EVAL_67;
  wire [3:0] fixer__EVAL_68;
  wire  fixer__EVAL_69;
  wire  fixer__EVAL_70;
  wire  fixer__EVAL_71;
  wire  fixer__EVAL_72;
  wire  fixer__EVAL_73;
  wire  fixer__EVAL_74;
  wire  fixer__EVAL_75;
  wire [2:0] fixer__EVAL_76;
  wire  fixer__EVAL_77;
  wire  fixer__EVAL_78;
  wire [31:0] fixer__EVAL_79;
  wire  fixer__EVAL_80;
  wire  fixer__EVAL_81;
  wire [2:0] fixer__EVAL_82;
  wire  fixer__EVAL_83;
  wire [3:0] fixer__EVAL_84;
  wire  fixer__EVAL_85;
  wire  fixer__EVAL_86;
  wire [3:0] fixer__EVAL_87;
  wire [31:0] fixer__EVAL_88;
  wire [31:0] fixer__EVAL_89;
  wire [3:0] fixer__EVAL_90;
  wire [3:0] fixer__EVAL_91;
  wire  fixer__EVAL_92;
  wire  fixer__EVAL_93;
  wire [2:0] fixer__EVAL_94;
  wire [31:0] fixer__EVAL_95;
  wire  fixer__EVAL_96;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire [2:0] _EVAL_213;
  wire  _EVAL_214;
  wire [3:0] _EVAL_215;
  wire [1:0] _EVAL_216;
  wire [2:0] _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire [4:0] _EVAL_220;
  wire [31:0] _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire [2:0] _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire [2:0] _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire [2:0] _EVAL_234;
  wire [2:0] _EVAL_235;
  wire [4:0] _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire [2:0] _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire [1:0] _EVAL_246;
  wire  _EVAL_247;
  wire [31:0] _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire [4:0] _EVAL_254;
  wire [2:0] _EVAL_255;
  wire [31:0] _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire [2:0] _EVAL_259;
  wire [1:0] _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire [2:0] _EVAL_267;
  wire [31:0] _EVAL_268;
  wire [31:0] _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire [3:0] _EVAL_272;
  wire  _EVAL_273;
  wire [3:0] _EVAL_274;
  wire  _EVAL_275;
  wire  coupler_to_port_named_ahb_sys_port__EVAL;
  wire [4:0] coupler_to_port_named_ahb_sys_port__EVAL_0;
  wire [31:0] coupler_to_port_named_ahb_sys_port__EVAL_1;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_2;
  wire [30:0] coupler_to_port_named_ahb_sys_port__EVAL_3;
  wire [2:0] coupler_to_port_named_ahb_sys_port__EVAL_4;
  wire [2:0] coupler_to_port_named_ahb_sys_port__EVAL_5;
  wire [31:0] coupler_to_port_named_ahb_sys_port__EVAL_6;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_7;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_8;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_9;
  wire [30:0] coupler_to_port_named_ahb_sys_port__EVAL_10;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_11;
  wire [2:0] coupler_to_port_named_ahb_sys_port__EVAL_12;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_13;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_14;
  wire [2:0] coupler_to_port_named_ahb_sys_port__EVAL_15;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_16;
  wire [4:0] coupler_to_port_named_ahb_sys_port__EVAL_17;
  wire [1:0] coupler_to_port_named_ahb_sys_port__EVAL_18;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_19;
  wire [2:0] coupler_to_port_named_ahb_sys_port__EVAL_20;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_21;
  wire [3:0] coupler_to_port_named_ahb_sys_port__EVAL_22;
  wire [1:0] coupler_to_port_named_ahb_sys_port__EVAL_23;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_24;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_25;
  wire [3:0] coupler_to_port_named_ahb_sys_port__EVAL_26;
  wire [31:0] coupler_to_port_named_ahb_sys_port__EVAL_27;
  wire [2:0] coupler_to_port_named_ahb_sys_port__EVAL_28;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_29;
  wire [2:0] coupler_to_port_named_ahb_sys_port__EVAL_30;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_31;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_32;
  wire [31:0] coupler_to_port_named_ahb_sys_port__EVAL_33;
  wire  coupler_to_port_named_ahb_sys_port__EVAL_34;
  wire [31:0] _EVAL_276;
  wire [31:0] _EVAL_277;
  wire [2:0] _EVAL_278;
  wire [2:0] _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire [3:0] _EVAL_286;
  wire [31:0] _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire [4:0] _EVAL_290;
  wire  _EVAL_291;
  wire [2:0] _EVAL_292;
  wire  _EVAL_293;
  wire [2:0] _EVAL_294;
  wire  _EVAL_295;
  wire  _EVAL_296;
  wire  _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire [31:0] _EVAL_307;
  wire  _EVAL_308;
  wire  _EVAL_309;
  wire  _EVAL_310;
  wire  _EVAL_311;
  wire [2:0] _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_314;
  wire [31:0] _EVAL_315;
  wire [3:0] _EVAL_316;
  wire [3:0] _EVAL_317;
  wire [3:0] _EVAL_318;
  wire  _EVAL_319;
  wire [3:0] _EVAL_320;
  wire [3:0] _EVAL_321;
  wire  _EVAL_322;
  wire  _EVAL_323;
  wire [31:0] _EVAL_324;
  wire  _EVAL_325;
  wire [1:0] _EVAL_326;
  wire  _EVAL_327;
  wire [2:0] _EVAL_328;
  wire  _EVAL_329;
  wire [1:0] _EVAL_330;
  wire [3:0] _EVAL_331;
  wire  _EVAL_332;
  wire [31:0] _EVAL_333;
  wire [3:0] _EVAL_334;
  _EVAL_0 fixedClockNode (
    ._EVAL(fixedClockNode__EVAL),
    ._EVAL_0(fixedClockNode__EVAL_0),
    ._EVAL_1(fixedClockNode__EVAL_1),
    ._EVAL_2(fixedClockNode__EVAL_2)
  );
  _EVAL_12 coupler_from_tile (
    ._EVAL(coupler_from_tile__EVAL),
    ._EVAL_0(coupler_from_tile__EVAL_0),
    ._EVAL_1(coupler_from_tile__EVAL_1),
    ._EVAL_2(coupler_from_tile__EVAL_2),
    ._EVAL_3(coupler_from_tile__EVAL_3),
    ._EVAL_4(coupler_from_tile__EVAL_4),
    ._EVAL_5(coupler_from_tile__EVAL_5),
    ._EVAL_6(coupler_from_tile__EVAL_6),
    ._EVAL_7(coupler_from_tile__EVAL_7),
    ._EVAL_8(coupler_from_tile__EVAL_8),
    ._EVAL_9(coupler_from_tile__EVAL_9),
    ._EVAL_10(coupler_from_tile__EVAL_10),
    ._EVAL_11(coupler_from_tile__EVAL_11),
    ._EVAL_12(coupler_from_tile__EVAL_12),
    ._EVAL_13(coupler_from_tile__EVAL_13),
    ._EVAL_14(coupler_from_tile__EVAL_14),
    ._EVAL_15(coupler_from_tile__EVAL_15),
    ._EVAL_16(coupler_from_tile__EVAL_16),
    ._EVAL_17(coupler_from_tile__EVAL_17),
    ._EVAL_18(coupler_from_tile__EVAL_18),
    ._EVAL_19(coupler_from_tile__EVAL_19),
    ._EVAL_20(coupler_from_tile__EVAL_20),
    ._EVAL_21(coupler_from_tile__EVAL_21),
    ._EVAL_22(coupler_from_tile__EVAL_22),
    ._EVAL_23(coupler_from_tile__EVAL_23),
    ._EVAL_24(coupler_from_tile__EVAL_24),
    ._EVAL_25(coupler_from_tile__EVAL_25),
    ._EVAL_26(coupler_from_tile__EVAL_26),
    ._EVAL_27(coupler_from_tile__EVAL_27),
    ._EVAL_28(coupler_from_tile__EVAL_28),
    ._EVAL_29(coupler_from_tile__EVAL_29),
    ._EVAL_30(coupler_from_tile__EVAL_30),
    ._EVAL_31(coupler_from_tile__EVAL_31),
    ._EVAL_32(coupler_from_tile__EVAL_32),
    ._EVAL_33(coupler_from_tile__EVAL_33),
    ._EVAL_34(coupler_from_tile__EVAL_34),
    ._EVAL_35(coupler_from_tile__EVAL_35),
    ._EVAL_36(coupler_from_tile__EVAL_36),
    ._EVAL_37(coupler_from_tile__EVAL_37),
    ._EVAL_38(coupler_from_tile__EVAL_38),
    ._EVAL_39(coupler_from_tile__EVAL_39),
    ._EVAL_40(coupler_from_tile__EVAL_40),
    ._EVAL_41(coupler_from_tile__EVAL_41),
    ._EVAL_42(coupler_from_tile__EVAL_42),
    ._EVAL_43(coupler_from_tile__EVAL_43),
    ._EVAL_44(coupler_from_tile__EVAL_44),
    ._EVAL_45(coupler_from_tile__EVAL_45),
    ._EVAL_46(coupler_from_tile__EVAL_46),
    ._EVAL_47(coupler_from_tile__EVAL_47),
    ._EVAL_48(coupler_from_tile__EVAL_48),
    ._EVAL_49(coupler_from_tile__EVAL_49),
    ._EVAL_50(coupler_from_tile__EVAL_50),
    ._EVAL_51(coupler_from_tile__EVAL_51),
    ._EVAL_52(coupler_from_tile__EVAL_52),
    ._EVAL_53(coupler_from_tile__EVAL_53),
    ._EVAL_54(coupler_from_tile__EVAL_54),
    ._EVAL_55(coupler_from_tile__EVAL_55),
    ._EVAL_56(coupler_from_tile__EVAL_56),
    ._EVAL_57(coupler_from_tile__EVAL_57),
    ._EVAL_58(coupler_from_tile__EVAL_58),
    ._EVAL_59(coupler_from_tile__EVAL_59),
    ._EVAL_60(coupler_from_tile__EVAL_60),
    ._EVAL_61(coupler_from_tile__EVAL_61),
    ._EVAL_62(coupler_from_tile__EVAL_62),
    ._EVAL_63(coupler_from_tile__EVAL_63),
    ._EVAL_64(coupler_from_tile__EVAL_64),
    ._EVAL_65(coupler_from_tile__EVAL_65),
    ._EVAL_66(coupler_from_tile__EVAL_66),
    ._EVAL_67(coupler_from_tile__EVAL_67),
    ._EVAL_68(coupler_from_tile__EVAL_68),
    ._EVAL_69(coupler_from_tile__EVAL_69),
    ._EVAL_70(coupler_from_tile__EVAL_70),
    ._EVAL_71(coupler_from_tile__EVAL_71),
    ._EVAL_72(coupler_from_tile__EVAL_72)
  );
  _EVAL_3 system_bus_xbar (
    ._EVAL(system_bus_xbar__EVAL),
    ._EVAL_0(system_bus_xbar__EVAL_0),
    ._EVAL_1(system_bus_xbar__EVAL_1),
    ._EVAL_2(system_bus_xbar__EVAL_2),
    ._EVAL_3(system_bus_xbar__EVAL_3),
    ._EVAL_4(system_bus_xbar__EVAL_4),
    ._EVAL_5(system_bus_xbar__EVAL_5),
    ._EVAL_6(system_bus_xbar__EVAL_6),
    ._EVAL_7(system_bus_xbar__EVAL_7),
    ._EVAL_8(system_bus_xbar__EVAL_8),
    ._EVAL_9(system_bus_xbar__EVAL_9),
    ._EVAL_10(system_bus_xbar__EVAL_10),
    ._EVAL_11(system_bus_xbar__EVAL_11),
    ._EVAL_12(system_bus_xbar__EVAL_12),
    ._EVAL_13(system_bus_xbar__EVAL_13),
    ._EVAL_14(system_bus_xbar__EVAL_14),
    ._EVAL_15(system_bus_xbar__EVAL_15),
    ._EVAL_16(system_bus_xbar__EVAL_16),
    ._EVAL_17(system_bus_xbar__EVAL_17),
    ._EVAL_18(system_bus_xbar__EVAL_18),
    ._EVAL_19(system_bus_xbar__EVAL_19),
    ._EVAL_20(system_bus_xbar__EVAL_20),
    ._EVAL_21(system_bus_xbar__EVAL_21),
    ._EVAL_22(system_bus_xbar__EVAL_22),
    ._EVAL_23(system_bus_xbar__EVAL_23),
    ._EVAL_24(system_bus_xbar__EVAL_24),
    ._EVAL_25(system_bus_xbar__EVAL_25),
    ._EVAL_26(system_bus_xbar__EVAL_26),
    ._EVAL_27(system_bus_xbar__EVAL_27),
    ._EVAL_28(system_bus_xbar__EVAL_28),
    ._EVAL_29(system_bus_xbar__EVAL_29),
    ._EVAL_30(system_bus_xbar__EVAL_30),
    ._EVAL_31(system_bus_xbar__EVAL_31),
    ._EVAL_32(system_bus_xbar__EVAL_32),
    ._EVAL_33(system_bus_xbar__EVAL_33),
    ._EVAL_34(system_bus_xbar__EVAL_34),
    ._EVAL_35(system_bus_xbar__EVAL_35),
    ._EVAL_36(system_bus_xbar__EVAL_36),
    ._EVAL_37(system_bus_xbar__EVAL_37),
    ._EVAL_38(system_bus_xbar__EVAL_38),
    ._EVAL_39(system_bus_xbar__EVAL_39),
    ._EVAL_40(system_bus_xbar__EVAL_40),
    ._EVAL_41(system_bus_xbar__EVAL_41),
    ._EVAL_42(system_bus_xbar__EVAL_42),
    ._EVAL_43(system_bus_xbar__EVAL_43),
    ._EVAL_44(system_bus_xbar__EVAL_44),
    ._EVAL_45(system_bus_xbar__EVAL_45),
    ._EVAL_46(system_bus_xbar__EVAL_46),
    ._EVAL_47(system_bus_xbar__EVAL_47),
    ._EVAL_48(system_bus_xbar__EVAL_48),
    ._EVAL_49(system_bus_xbar__EVAL_49),
    ._EVAL_50(system_bus_xbar__EVAL_50),
    ._EVAL_51(system_bus_xbar__EVAL_51),
    ._EVAL_52(system_bus_xbar__EVAL_52),
    ._EVAL_53(system_bus_xbar__EVAL_53),
    ._EVAL_54(system_bus_xbar__EVAL_54),
    ._EVAL_55(system_bus_xbar__EVAL_55),
    ._EVAL_56(system_bus_xbar__EVAL_56),
    ._EVAL_57(system_bus_xbar__EVAL_57),
    ._EVAL_58(system_bus_xbar__EVAL_58),
    ._EVAL_59(system_bus_xbar__EVAL_59),
    ._EVAL_60(system_bus_xbar__EVAL_60),
    ._EVAL_61(system_bus_xbar__EVAL_61),
    ._EVAL_62(system_bus_xbar__EVAL_62),
    ._EVAL_63(system_bus_xbar__EVAL_63),
    ._EVAL_64(system_bus_xbar__EVAL_64),
    ._EVAL_65(system_bus_xbar__EVAL_65),
    ._EVAL_66(system_bus_xbar__EVAL_66),
    ._EVAL_67(system_bus_xbar__EVAL_67),
    ._EVAL_68(system_bus_xbar__EVAL_68),
    ._EVAL_69(system_bus_xbar__EVAL_69),
    ._EVAL_70(system_bus_xbar__EVAL_70),
    ._EVAL_71(system_bus_xbar__EVAL_71),
    ._EVAL_72(system_bus_xbar__EVAL_72),
    ._EVAL_73(system_bus_xbar__EVAL_73),
    ._EVAL_74(system_bus_xbar__EVAL_74),
    ._EVAL_75(system_bus_xbar__EVAL_75),
    ._EVAL_76(system_bus_xbar__EVAL_76),
    ._EVAL_77(system_bus_xbar__EVAL_77),
    ._EVAL_78(system_bus_xbar__EVAL_78),
    ._EVAL_79(system_bus_xbar__EVAL_79),
    ._EVAL_80(system_bus_xbar__EVAL_80),
    ._EVAL_81(system_bus_xbar__EVAL_81),
    ._EVAL_82(system_bus_xbar__EVAL_82),
    ._EVAL_83(system_bus_xbar__EVAL_83),
    ._EVAL_84(system_bus_xbar__EVAL_84),
    ._EVAL_85(system_bus_xbar__EVAL_85),
    ._EVAL_86(system_bus_xbar__EVAL_86),
    ._EVAL_87(system_bus_xbar__EVAL_87),
    ._EVAL_88(system_bus_xbar__EVAL_88),
    ._EVAL_89(system_bus_xbar__EVAL_89),
    ._EVAL_90(system_bus_xbar__EVAL_90),
    ._EVAL_91(system_bus_xbar__EVAL_91),
    ._EVAL_92(system_bus_xbar__EVAL_92),
    ._EVAL_93(system_bus_xbar__EVAL_93),
    ._EVAL_94(system_bus_xbar__EVAL_94),
    ._EVAL_95(system_bus_xbar__EVAL_95),
    ._EVAL_96(system_bus_xbar__EVAL_96)
  );
  _EVAL_6 fixer (
    ._EVAL(fixer__EVAL),
    ._EVAL_0(fixer__EVAL_0),
    ._EVAL_1(fixer__EVAL_1),
    ._EVAL_2(fixer__EVAL_2),
    ._EVAL_3(fixer__EVAL_3),
    ._EVAL_4(fixer__EVAL_4),
    ._EVAL_5(fixer__EVAL_5),
    ._EVAL_6(fixer__EVAL_6),
    ._EVAL_7(fixer__EVAL_7),
    ._EVAL_8(fixer__EVAL_8),
    ._EVAL_9(fixer__EVAL_9),
    ._EVAL_10(fixer__EVAL_10),
    ._EVAL_11(fixer__EVAL_11),
    ._EVAL_12(fixer__EVAL_12),
    ._EVAL_13(fixer__EVAL_13),
    ._EVAL_14(fixer__EVAL_14),
    ._EVAL_15(fixer__EVAL_15),
    ._EVAL_16(fixer__EVAL_16),
    ._EVAL_17(fixer__EVAL_17),
    ._EVAL_18(fixer__EVAL_18),
    ._EVAL_19(fixer__EVAL_19),
    ._EVAL_20(fixer__EVAL_20),
    ._EVAL_21(fixer__EVAL_21),
    ._EVAL_22(fixer__EVAL_22),
    ._EVAL_23(fixer__EVAL_23),
    ._EVAL_24(fixer__EVAL_24),
    ._EVAL_25(fixer__EVAL_25),
    ._EVAL_26(fixer__EVAL_26),
    ._EVAL_27(fixer__EVAL_27),
    ._EVAL_28(fixer__EVAL_28),
    ._EVAL_29(fixer__EVAL_29),
    ._EVAL_30(fixer__EVAL_30),
    ._EVAL_31(fixer__EVAL_31),
    ._EVAL_32(fixer__EVAL_32),
    ._EVAL_33(fixer__EVAL_33),
    ._EVAL_34(fixer__EVAL_34),
    ._EVAL_35(fixer__EVAL_35),
    ._EVAL_36(fixer__EVAL_36),
    ._EVAL_37(fixer__EVAL_37),
    ._EVAL_38(fixer__EVAL_38),
    ._EVAL_39(fixer__EVAL_39),
    ._EVAL_40(fixer__EVAL_40),
    ._EVAL_41(fixer__EVAL_41),
    ._EVAL_42(fixer__EVAL_42),
    ._EVAL_43(fixer__EVAL_43),
    ._EVAL_44(fixer__EVAL_44),
    ._EVAL_45(fixer__EVAL_45),
    ._EVAL_46(fixer__EVAL_46),
    ._EVAL_47(fixer__EVAL_47),
    ._EVAL_48(fixer__EVAL_48),
    ._EVAL_49(fixer__EVAL_49),
    ._EVAL_50(fixer__EVAL_50),
    ._EVAL_51(fixer__EVAL_51),
    ._EVAL_52(fixer__EVAL_52),
    ._EVAL_53(fixer__EVAL_53),
    ._EVAL_54(fixer__EVAL_54),
    ._EVAL_55(fixer__EVAL_55),
    ._EVAL_56(fixer__EVAL_56),
    ._EVAL_57(fixer__EVAL_57),
    ._EVAL_58(fixer__EVAL_58),
    ._EVAL_59(fixer__EVAL_59),
    ._EVAL_60(fixer__EVAL_60),
    ._EVAL_61(fixer__EVAL_61),
    ._EVAL_62(fixer__EVAL_62),
    ._EVAL_63(fixer__EVAL_63),
    ._EVAL_64(fixer__EVAL_64),
    ._EVAL_65(fixer__EVAL_65),
    ._EVAL_66(fixer__EVAL_66),
    ._EVAL_67(fixer__EVAL_67),
    ._EVAL_68(fixer__EVAL_68),
    ._EVAL_69(fixer__EVAL_69),
    ._EVAL_70(fixer__EVAL_70),
    ._EVAL_71(fixer__EVAL_71),
    ._EVAL_72(fixer__EVAL_72),
    ._EVAL_73(fixer__EVAL_73),
    ._EVAL_74(fixer__EVAL_74),
    ._EVAL_75(fixer__EVAL_75),
    ._EVAL_76(fixer__EVAL_76),
    ._EVAL_77(fixer__EVAL_77),
    ._EVAL_78(fixer__EVAL_78),
    ._EVAL_79(fixer__EVAL_79),
    ._EVAL_80(fixer__EVAL_80),
    ._EVAL_81(fixer__EVAL_81),
    ._EVAL_82(fixer__EVAL_82),
    ._EVAL_83(fixer__EVAL_83),
    ._EVAL_84(fixer__EVAL_84),
    ._EVAL_85(fixer__EVAL_85),
    ._EVAL_86(fixer__EVAL_86),
    ._EVAL_87(fixer__EVAL_87),
    ._EVAL_88(fixer__EVAL_88),
    ._EVAL_89(fixer__EVAL_89),
    ._EVAL_90(fixer__EVAL_90),
    ._EVAL_91(fixer__EVAL_91),
    ._EVAL_92(fixer__EVAL_92),
    ._EVAL_93(fixer__EVAL_93),
    ._EVAL_94(fixer__EVAL_94),
    ._EVAL_95(fixer__EVAL_95),
    ._EVAL_96(fixer__EVAL_96)
  );
  _EVAL_21 coupler_to_port_named_ahb_sys_port (
    ._EVAL(coupler_to_port_named_ahb_sys_port__EVAL),
    ._EVAL_0(coupler_to_port_named_ahb_sys_port__EVAL_0),
    ._EVAL_1(coupler_to_port_named_ahb_sys_port__EVAL_1),
    ._EVAL_2(coupler_to_port_named_ahb_sys_port__EVAL_2),
    ._EVAL_3(coupler_to_port_named_ahb_sys_port__EVAL_3),
    ._EVAL_4(coupler_to_port_named_ahb_sys_port__EVAL_4),
    ._EVAL_5(coupler_to_port_named_ahb_sys_port__EVAL_5),
    ._EVAL_6(coupler_to_port_named_ahb_sys_port__EVAL_6),
    ._EVAL_7(coupler_to_port_named_ahb_sys_port__EVAL_7),
    ._EVAL_8(coupler_to_port_named_ahb_sys_port__EVAL_8),
    ._EVAL_9(coupler_to_port_named_ahb_sys_port__EVAL_9),
    ._EVAL_10(coupler_to_port_named_ahb_sys_port__EVAL_10),
    ._EVAL_11(coupler_to_port_named_ahb_sys_port__EVAL_11),
    ._EVAL_12(coupler_to_port_named_ahb_sys_port__EVAL_12),
    ._EVAL_13(coupler_to_port_named_ahb_sys_port__EVAL_13),
    ._EVAL_14(coupler_to_port_named_ahb_sys_port__EVAL_14),
    ._EVAL_15(coupler_to_port_named_ahb_sys_port__EVAL_15),
    ._EVAL_16(coupler_to_port_named_ahb_sys_port__EVAL_16),
    ._EVAL_17(coupler_to_port_named_ahb_sys_port__EVAL_17),
    ._EVAL_18(coupler_to_port_named_ahb_sys_port__EVAL_18),
    ._EVAL_19(coupler_to_port_named_ahb_sys_port__EVAL_19),
    ._EVAL_20(coupler_to_port_named_ahb_sys_port__EVAL_20),
    ._EVAL_21(coupler_to_port_named_ahb_sys_port__EVAL_21),
    ._EVAL_22(coupler_to_port_named_ahb_sys_port__EVAL_22),
    ._EVAL_23(coupler_to_port_named_ahb_sys_port__EVAL_23),
    ._EVAL_24(coupler_to_port_named_ahb_sys_port__EVAL_24),
    ._EVAL_25(coupler_to_port_named_ahb_sys_port__EVAL_25),
    ._EVAL_26(coupler_to_port_named_ahb_sys_port__EVAL_26),
    ._EVAL_27(coupler_to_port_named_ahb_sys_port__EVAL_27),
    ._EVAL_28(coupler_to_port_named_ahb_sys_port__EVAL_28),
    ._EVAL_29(coupler_to_port_named_ahb_sys_port__EVAL_29),
    ._EVAL_30(coupler_to_port_named_ahb_sys_port__EVAL_30),
    ._EVAL_31(coupler_to_port_named_ahb_sys_port__EVAL_31),
    ._EVAL_32(coupler_to_port_named_ahb_sys_port__EVAL_32),
    ._EVAL_33(coupler_to_port_named_ahb_sys_port__EVAL_33),
    ._EVAL_34(coupler_to_port_named_ahb_sys_port__EVAL_34)
  );
  assign _EVAL_182 = _EVAL_315;
  assign _EVAL_261 = _EVAL_134;
  assign _EVAL_156 = system_bus_xbar__EVAL_45;
  assign coupler_to_port_named_ahb_sys_port__EVAL_2 = system_bus_xbar__EVAL_93;
  assign _EVAL_192 = system_bus_xbar__EVAL_2;
  assign fixer__EVAL_1 = _EVAL_232;
  assign _EVAL_84 = _EVAL_314;
  assign coupler_from_tile__EVAL_26 = _EVAL_44;
  assign fixer__EVAL_69 = system_bus_xbar__EVAL_46;
  assign _EVAL_249 = _EVAL_285;
  assign system_bus_xbar__EVAL_68 = coupler_to_port_named_ahb_sys_port__EVAL_29;
  assign coupler_from_tile__EVAL_63 = _EVAL_66;
  assign _EVAL_304 = _EVAL_76;
  assign _EVAL_323 = _EVAL_142;
  assign _EVAL_48 = coupler_from_tile__EVAL_53;
  assign _EVAL_97 = coupler_from_tile__EVAL_20;
  assign system_bus_xbar__EVAL_56 = coupler_to_port_named_ahb_sys_port__EVAL_4;
  assign coupler_to_port_named_ahb_sys_port__EVAL_15 = system_bus_xbar__EVAL_51;
  assign _EVAL_1 = coupler_from_tile__EVAL_41;
  assign fixer__EVAL_41 = system_bus_xbar__EVAL_85;
  assign _EVAL_316 = fixer__EVAL_13;
  assign _EVAL_30 = _EVAL_249;
  assign _EVAL_306 = _EVAL_156;
  assign _EVAL_267 = _EVAL_217;
  assign fixer__EVAL_18 = coupler_from_tile__EVAL_29;
  assign _EVAL_170 = _EVAL_290;
  assign _EVAL_138 = _EVAL_204;
  assign _EVAL_324 = _EVAL_164;
  assign _EVAL_143 = _EVAL_188;
  assign _EVAL_127 = system_bus_xbar__EVAL_86;
  assign _EVAL_256 = _EVAL_123;
  assign system_bus_xbar__EVAL_11 = fixer__EVAL_0;
  assign _EVAL_199 = _EVAL_146;
  assign coupler_to_port_named_ahb_sys_port__EVAL_13 = system_bus_xbar__EVAL_44;
  assign _EVAL_290 = _EVAL_167;
  assign system_bus_xbar__EVAL_6 = fixer__EVAL_67;
  assign fixer__EVAL_56 = coupler_from_tile__EVAL_17;
  assign _EVAL_302 = _EVAL_135;
  assign fixer__EVAL_90 = coupler_from_tile__EVAL_38;
  assign _EVAL_235 = _EVAL_199;
  assign _EVAL_150 = _EVAL_177;
  assign _EVAL_334 = _EVAL_131;
  assign _EVAL_154 = _EVAL_306;
  assign _EVAL_244 = _EVAL_253;
  assign _EVAL_260 = _EVAL_330;
  assign system_bus_xbar__EVAL_74 = fixer__EVAL_6;
  assign _EVAL_189 = _EVAL_251;
  assign _EVAL_231 = _EVAL_166;
  assign _EVAL_59 = coupler_to_port_named_ahb_sys_port__EVAL_30;
  assign _EVAL_320 = _EVAL_272;
  assign system_bus_xbar__EVAL_16 = fixer__EVAL_95;
  assign _EVAL_225 = _EVAL_231;
  assign _EVAL_110 = coupler_from_tile__EVAL_25;
  assign _EVAL_292 = _EVAL_255;
  assign _EVAL_99 = _EVAL_145;
  assign _EVAL_20 = _EVAL_263;
  assign _EVAL_224 = _EVAL_280;
  assign coupler_from_tile__EVAL_46 = fixer__EVAL_40;
  assign _EVAL_137 = _EVAL_308;
  assign system_bus_xbar__EVAL_5 = fixer__EVAL_87;
  assign system_bus_xbar__EVAL_36 = fixer__EVAL_32;
  assign _EVAL_2 = coupler_from_tile__EVAL_34;
  assign _EVAL_147 = _EVAL_201;
  assign _EVAL_181 = _EVAL_286;
  assign fixer__EVAL_91 = system_bus_xbar__EVAL_60;
  assign _EVAL_126 = _EVAL_154;
  assign fixer__EVAL_16 = system_bus_xbar__EVAL_15;
  assign _EVAL_180 = _EVAL_276;
  assign fixer__EVAL_31 = coupler_from_tile__EVAL_59;
  assign _EVAL_221 = _EVAL_287;
  assign fixer__EVAL_47 = coupler_from_tile__EVAL_42;
  assign _EVAL_28 = coupler_to_port_named_ahb_sys_port__EVAL_26;
  assign fixer__EVAL_81 = coupler_from_tile__EVAL_7;
  assign fixer__EVAL_70 = fixedClockNode__EVAL;
  assign _EVAL_294 = _EVAL_239;
  assign _EVAL_140 = _EVAL_288;
  assign _EVAL_117 = coupler_from_tile__EVAL_9;
  assign _EVAL_161 = _EVAL_111;
  assign _EVAL_133 = _EVAL_68;
  assign _EVAL_206 = _EVAL_189;
  assign _EVAL_187 = _EVAL_172;
  assign coupler_from_tile__EVAL_57 = _EVAL_23;
  assign system_bus_xbar__EVAL_75 = fixer__EVAL_86;
  assign _EVAL_227 = _EVAL_311;
  assign _EVAL_136 = _EVAL_268;
  assign _EVAL_169 = _EVAL_128;
  assign _EVAL_74 = coupler_from_tile__EVAL_28;
  assign _EVAL_195 = fixer__EVAL_36;
  assign fixedClockNode__EVAL_2 = _EVAL_183;
  assign system_bus_xbar__EVAL_20 = coupler_to_port_named_ahb_sys_port__EVAL_28;
  assign _EVAL_175 = _EVAL_26;
  assign coupler_from_tile__EVAL_61 = _EVAL_49;
  assign _EVAL_258 = _EVAL_91;
  assign _EVAL_146 = fixer__EVAL_25;
  assign system_bus_xbar__EVAL_21 = coupler_to_port_named_ahb_sys_port__EVAL_18;
  assign _EVAL_308 = system_bus_xbar__EVAL_35;
  assign _EVAL_46 = _EVAL_260;
  assign _EVAL_135 = _EVAL_233;
  assign _EVAL_270 = system_bus_xbar__EVAL_90;
  assign system_bus_xbar__EVAL_96 = _EVAL_180;
  assign coupler_to_port_named_ahb_sys_port__EVAL_10 = system_bus_xbar__EVAL_47;
  assign coupler_from_tile__EVAL_58 = _EVAL_6;
  assign _EVAL_25 = _EVAL_221;
  assign _EVAL_286 = _EVAL_321;
  assign coupler_from_tile__EVAL_2 = fixer__EVAL_23;
  assign _EVAL_149 = _EVAL_160;
  assign fixer__EVAL_38 = system_bus_xbar__EVAL_24;
  assign _EVAL_247 = _EVAL_211;
  assign _EVAL_220 = _EVAL_254;
  assign _EVAL_144 = _EVAL_318;
  assign _EVAL_153 = _EVAL_122;
  assign _EVAL_159 = _EVAL_206;
  assign _EVAL_212 = _EVAL_283;
  assign coupler_from_tile__EVAL_27 = _EVAL_31;
  assign _EVAL_278 = system_bus_xbar__EVAL_66;
  assign _EVAL_124 = _EVAL_197;
  assign _EVAL_72 = _EVAL_310;
  assign _EVAL_114 = _EVAL_317;
  assign coupler_from_tile__EVAL_21 = _EVAL_64;
  assign _EVAL_311 = _EVAL_195;
  assign system_bus_xbar__EVAL_30 = fixer__EVAL_74;
  assign _EVAL_276 = _EVAL_324;
  assign system_bus_xbar__EVAL_64 = fixer__EVAL_34;
  assign _EVAL_312 = _EVAL_101;
  assign _EVAL_300 = fixer__EVAL_55;
  assign _EVAL_157 = _EVAL_307;
  assign _EVAL_313 = _EVAL_4;
  assign coupler_from_tile__EVAL_64 = _EVAL_69;
  assign _EVAL_250 = fixer__EVAL_83;
  assign system_bus_xbar__EVAL_94 = fixer__EVAL_35;
  assign fixer__EVAL_63 = system_bus_xbar__EVAL_3;
  assign _EVAL_315 = _EVAL_157;
  assign system_bus_xbar__EVAL_57 = _EVAL_262;
  assign coupler_from_tile__EVAL_22 = _EVAL_29;
  assign _EVAL_165 = _EVAL_208;
  assign _EVAL_115 = _EVAL_170;
  assign fixer__EVAL_45 = system_bus_xbar__EVAL_83;
  assign _EVAL_166 = _EVAL_148;
  assign _EVAL_265 = _EVAL_257;
  assign _EVAL_163 = system_bus_xbar__EVAL_17;
  assign coupler_from_tile__EVAL_60 = _EVAL_108;
  assign _EVAL_128 = _EVAL_305;
  assign _EVAL_85 = _EVAL_126;
  assign fixer__EVAL_17 = system_bus_xbar__EVAL_25;
  assign _EVAL_234 = _EVAL_209;
  assign fixer__EVAL_58 = _EVAL_267;
  assign _EVAL_272 = _EVAL_8;
  assign coupler_to_port_named_ahb_sys_port__EVAL_19 = _EVAL_113;
  assign system_bus_xbar__EVAL_54 = fixer__EVAL_82;
  assign _EVAL_203 = fixer__EVAL_88;
  assign coupler_to_port_named_ahb_sys_port__EVAL_0 = system_bus_xbar__EVAL_88;
  assign _EVAL_39 = _EVAL_248;
  assign fixer__EVAL_93 = system_bus_xbar__EVAL_59;
  assign _EVAL_232 = _EVAL_265;
  assign _EVAL_288 = _EVAL_120;
  assign _EVAL_240 = _EVAL_299;
  assign _EVAL_319 = _EVAL_186;
  assign fixer__EVAL_61 = _EVAL_243;
  assign _EVAL_213 = _EVAL_312;
  assign fixer__EVAL = _EVAL_256;
  assign fixer__EVAL_49 = coupler_from_tile__EVAL_10;
  assign _EVAL_139 = _EVAL_223;
  assign _EVAL_236 = _EVAL_133;
  assign system_bus_xbar__EVAL_58 = fixer__EVAL_54;
  assign _EVAL_201 = system_bus_xbar__EVAL_28;
  assign _EVAL_280 = fixer__EVAL_80;
  assign _EVAL_120 = _EVAL_27;
  assign _EVAL_222 = _EVAL_313;
  assign _EVAL_215 = _EVAL_130;
  assign _EVAL_179 = _EVAL_210;
  assign _EVAL_298 = _EVAL_152;
  assign _EVAL_214 = _EVAL_185;
  assign system_bus_xbar__EVAL_42 = coupler_to_port_named_ahb_sys_port__EVAL_8;
  assign system_bus_xbar__EVAL_31 = _EVAL_150;
  assign fixedClockNode__EVAL_1 = _EVAL_319;
  assign _EVAL_36 = coupler_from_tile__EVAL_71;
  assign fixer__EVAL_42 = system_bus_xbar__EVAL_13;
  assign _EVAL_141 = _EVAL_61;
  assign coupler_from_tile__EVAL_50 = fixer__EVAL_84;
  assign system_bus_xbar__EVAL_18 = fixer__EVAL_46;
  assign _EVAL_310 = _EVAL_329;
  assign _EVAL_327 = _EVAL_137;
  assign _EVAL_259 = _EVAL_294;
  assign _EVAL_11 = coupler_from_tile__EVAL_67;
  assign coupler_to_port_named_ahb_sys_port__EVAL_21 = system_bus_xbar__EVAL_67;
  assign coupler_from_tile__EVAL_43 = _EVAL_19;
  assign _EVAL_229 = _EVAL_191;
  assign _EVAL_148 = system_bus_xbar__EVAL_19;
  assign _EVAL_257 = _EVAL_304;
  assign _EVAL_207 = _EVAL_309;
  assign _EVAL_242 = _EVAL_3;
  assign fixer__EVAL_9 = system_bus_xbar__EVAL_76;
  assign _EVAL_228 = _EVAL_13;
  assign fixer__EVAL_15 = _EVAL_200;
  assign _EVAL_317 = _EVAL_215;
  assign _EVAL_325 = _EVAL_241;
  assign fixer__EVAL_11 = coupler_from_tile__EVAL_8;
  assign _EVAL_197 = _EVAL_247;
  assign _EVAL_16 = coupler_to_port_named_ahb_sys_port__EVAL_3;
  assign fixer__EVAL_92 = system_bus_xbar__EVAL_41;
  assign fixer__EVAL_39 = _EVAL_138;
  assign _EVAL_34 = _EVAL_119;
  assign _EVAL_177 = _EVAL_326;
  assign fixer__EVAL_14 = _EVAL_296;
  assign coupler_from_tile__EVAL_44 = _EVAL_55;
  assign _EVAL_217 = _EVAL_234;
  assign _EVAL_185 = _EVAL_238;
  assign coupler_to_port_named_ahb_sys_port__EVAL_11 = fixedClockNode__EVAL_0;
  assign _EVAL_204 = _EVAL_179;
  assign _EVAL_86 = coupler_to_port_named_ahb_sys_port__EVAL_33;
  assign _EVAL_134 = _EVAL_147;
  assign fixer__EVAL_89 = coupler_from_tile__EVAL_15;
  assign fixer__EVAL_2 = coupler_from_tile__EVAL_5;
  assign _EVAL_167 = _EVAL_173;
  assign _EVAL_121 = _EVAL_264;
  assign fixer__EVAL_4 = coupler_from_tile__EVAL_40;
  assign coupler_from_tile__EVAL_13 = _EVAL_78;
  assign _EVAL_190 = _EVAL_332;
  assign system_bus_xbar__EVAL_0 = fixer__EVAL_19;
  assign _EVAL_174 = _EVAL_139;
  assign fixer__EVAL_5 = _EVAL_281;
  assign _EVAL_299 = _EVAL_275;
  assign _EVAL_118 = _EVAL_190;
  assign system_bus_xbar__EVAL = fixedClockNode__EVAL_0;
  assign coupler_from_tile__EVAL_69 = _EVAL_79;
  assign _EVAL_282 = fixer__EVAL_72;
  assign system_bus_xbar__EVAL_48 = _EVAL_124;
  assign _EVAL_284 = _EVAL_228;
  assign _EVAL_287 = _EVAL_269;
  assign _EVAL_184 = _EVAL_271;
  assign _EVAL_122 = _EVAL_24;
  assign _EVAL_38 = coupler_to_port_named_ahb_sys_port__EVAL_23;
  assign _EVAL_330 = _EVAL_246;
  assign _EVAL_307 = _EVAL_47;
  assign system_bus_xbar__EVAL_71 = coupler_to_port_named_ahb_sys_port__EVAL_7;
  assign _EVAL_331 = _EVAL_165;
  assign _EVAL_248 = _EVAL_143;
  assign system_bus_xbar__EVAL_70 = fixer__EVAL_20;
  assign _EVAL_239 = _EVAL_73;
  assign system_bus_xbar__EVAL_10 = fixedClockNode__EVAL;
  assign _EVAL_241 = _EVAL_116;
  assign coupler_to_port_named_ahb_sys_port__EVAL_12 = system_bus_xbar__EVAL_40;
  assign coupler_from_tile__EVAL_16 = _EVAL_15;
  assign _EVAL_321 = _EVAL_178;
  assign _EVAL_252 = _EVAL_322;
  assign _EVAL_132 = _EVAL_218;
  assign _EVAL_129 = _EVAL_121;
  assign coupler_from_tile__EVAL_45 = _EVAL_90;
  assign _EVAL_216 = fixer__EVAL_7;
  assign coupler_to_port_named_ahb_sys_port__EVAL_14 = system_bus_xbar__EVAL_12;
  assign fixer__EVAL_76 = system_bus_xbar__EVAL_84;
  assign coupler_to_port_named_ahb_sys_port__EVAL_6 = system_bus_xbar__EVAL_8;
  assign fixer__EVAL_78 = coupler_from_tile__EVAL_54;
  assign _EVAL_211 = _EVAL_10;
  assign _EVAL_208 = _EVAL_192;
  assign _EVAL_243 = _EVAL_196;
  assign _EVAL_155 = _EVAL_274;
  assign _EVAL_273 = _EVAL_300;
  assign _EVAL_130 = _EVAL_316;
  assign _EVAL_21 = _EVAL_225;
  assign _EVAL_295 = _EVAL_162;
  assign coupler_from_tile__EVAL_24 = fixer__EVAL_29;
  assign _EVAL_266 = _EVAL_327;
  assign fixer__EVAL_22 = _EVAL_303;
  assign _EVAL_297 = _EVAL_107;
  assign _EVAL_309 = _EVAL_54;
  assign _EVAL_318 = _EVAL_155;
  assign _EVAL_164 = _EVAL_18;
  assign _EVAL_160 = _EVAL_70;
  assign _EVAL_95 = _EVAL_298;
  assign coupler_from_tile__EVAL = _EVAL_81;
  assign coupler_from_tile__EVAL_4 = _EVAL_60;
  assign _EVAL_226 = _EVAL_12;
  assign system_bus_xbar__EVAL_89 = fixer__EVAL_51;
  assign system_bus_xbar__EVAL_61 = fixer__EVAL_96;
  assign _EVAL_205 = _EVAL_270;
  assign _EVAL_218 = _EVAL_141;
  assign _EVAL_237 = _EVAL_175;
  assign _EVAL_43 = _EVAL_159;
  assign _EVAL_183 = _EVAL_169;
  assign _EVAL_314 = _EVAL_202;
  assign system_bus_xbar__EVAL_78 = _EVAL_176;
  assign _EVAL_57 = coupler_to_port_named_ahb_sys_port__EVAL;
  assign system_bus_xbar__EVAL_32 = fixer__EVAL_60;
  assign system_bus_xbar__EVAL_77 = fixer__EVAL_26;
  assign coupler_from_tile__EVAL_68 = _EVAL_82;
  assign _EVAL_158 = _EVAL_302;
  assign system_bus_xbar__EVAL_14 = fixer__EVAL_77;
  assign coupler_from_tile__EVAL_49 = fixer__EVAL_62;
  assign _EVAL_219 = _EVAL_205;
  assign coupler_from_tile__EVAL_14 = _EVAL_63;
  assign fixer__EVAL_79 = system_bus_xbar__EVAL_23;
  assign fixer__EVAL_8 = coupler_from_tile__EVAL_31;
  assign system_bus_xbar__EVAL_91 = fixer__EVAL_68;
  assign _EVAL_35 = _EVAL_245;
  assign _EVAL_106 = _EVAL_240;
  assign _EVAL_303 = _EVAL_140;
  assign fixer__EVAL_27 = _EVAL_214;
  assign _EVAL_186 = _EVAL_325;
  assign _EVAL_210 = _EVAL_88;
  assign _EVAL_200 = _EVAL_252;
  assign _EVAL_281 = _EVAL_151;
  assign system_bus_xbar__EVAL_39 = fixer__EVAL_85;
  assign _EVAL_83 = coupler_from_tile__EVAL_70;
  assign _EVAL_328 = _EVAL_235;
  assign _EVAL_176 = _EVAL_171;
  assign coupler_to_port_named_ahb_sys_port__EVAL_32 = fixedClockNode__EVAL;
  assign _EVAL_71 = _EVAL_261;
  assign _EVAL_67 = coupler_from_tile__EVAL_11;
  assign _EVAL_80 = _EVAL_187;
  assign _EVAL_145 = _EVAL_333;
  assign _EVAL_50 = _EVAL_292;
  assign _EVAL_125 = _EVAL_259;
  assign fixer__EVAL_94 = _EVAL_125;
  assign system_bus_xbar__EVAL_69 = fixer__EVAL_73;
  assign _EVAL_194 = _EVAL_0;
  assign _EVAL_178 = system_bus_xbar__EVAL_95;
  assign _EVAL_209 = _EVAL_93;
  assign _EVAL_301 = _EVAL_297;
  assign fixer__EVAL_52 = _EVAL_182;
  assign _EVAL_251 = _EVAL_45;
  assign coupler_from_tile__EVAL_0 = fixer__EVAL_37;
  assign _EVAL_253 = fixer__EVAL_65;
  assign fixer__EVAL_44 = _EVAL_334;
  assign system_bus_xbar__EVAL_27 = coupler_to_port_named_ahb_sys_port__EVAL_9;
  assign _EVAL_5 = _EVAL_266;
  assign coupler_from_tile__EVAL_62 = fixer__EVAL_66;
  assign _EVAL_41 = coupler_to_port_named_ahb_sys_port__EVAL_20;
  assign _EVAL_238 = _EVAL_161;
  assign _EVAL_255 = _EVAL_279;
  assign _EVAL_285 = _EVAL_224;
  assign _EVAL_262 = _EVAL_132;
  assign coupler_from_tile__EVAL_36 = _EVAL_58;
  assign _EVAL_193 = _EVAL_227;
  assign system_bus_xbar__EVAL_1 = fixer__EVAL_64;
  assign _EVAL_89 = _EVAL_153;
  assign _EVAL_230 = system_bus_xbar__EVAL_55;
  assign coupler_from_tile__EVAL_30 = _EVAL_102;
  assign coupler_from_tile__EVAL_33 = fixedClockNode__EVAL_0;
  assign coupler_from_tile__EVAL_51 = fixer__EVAL_12;
  assign _EVAL_264 = _EVAL_242;
  assign _EVAL_94 = coupler_from_tile__EVAL_52;
  assign coupler_to_port_named_ahb_sys_port__EVAL_34 = _EVAL_103;
  assign _EVAL_162 = _EVAL_207;
  assign coupler_from_tile__EVAL_66 = fixer__EVAL_59;
  assign _EVAL_105 = coupler_from_tile__EVAL_65;
  assign coupler_from_tile__EVAL_56 = _EVAL_98;
  assign _EVAL_268 = _EVAL_14;
  assign coupler_to_port_named_ahb_sys_port__EVAL_16 = system_bus_xbar__EVAL_62;
  assign _EVAL_322 = _EVAL_226;
  assign _EVAL_171 = _EVAL_213;
  assign _EVAL_173 = system_bus_xbar__EVAL_38;
  assign _EVAL_293 = _EVAL_282;
  assign _EVAL_332 = _EVAL_244;
  assign _EVAL_245 = _EVAL_219;
  assign _EVAL_33 = coupler_from_tile__EVAL_1;
  assign coupler_from_tile__EVAL_48 = _EVAL_104;
  assign _EVAL_223 = system_bus_xbar__EVAL_22;
  assign _EVAL_168 = _EVAL_229;
  assign _EVAL_269 = _EVAL_198;
  assign _EVAL_65 = _EVAL_328;
  assign coupler_to_port_named_ahb_sys_port__EVAL_5 = system_bus_xbar__EVAL_81;
  assign coupler_to_port_named_ahb_sys_port__EVAL_25 = system_bus_xbar__EVAL_7;
  assign coupler_from_tile__EVAL_47 = _EVAL_51;
  assign _EVAL_283 = _EVAL_87;
  assign _EVAL_62 = _EVAL_181;
  assign fixer__EVAL_57 = system_bus_xbar__EVAL_33;
  assign _EVAL_53 = _EVAL_193;
  assign _EVAL_279 = _EVAL_278;
  assign _EVAL_152 = _EVAL_293;
  assign system_bus_xbar__EVAL_29 = fixer__EVAL_3;
  assign system_bus_xbar__EVAL_82 = fixer__EVAL_48;
  assign system_bus_xbar__EVAL_52 = _EVAL_220;
  assign _EVAL_246 = _EVAL_216;
  assign system_bus_xbar__EVAL_50 = coupler_to_port_named_ahb_sys_port__EVAL_17;
  assign _EVAL_40 = coupler_from_tile__EVAL_35;
  assign system_bus_xbar__EVAL_43 = fixer__EVAL_30;
  assign _EVAL_75 = _EVAL_301;
  assign _EVAL_131 = _EVAL_320;
  assign _EVAL_326 = _EVAL_194;
  assign _EVAL_42 = coupler_from_tile__EVAL_72;
  assign _EVAL_112 = _EVAL_331;
  assign _EVAL_296 = _EVAL_289;
  assign fixer__EVAL_50 = coupler_from_tile__EVAL_23;
  assign _EVAL_56 = _EVAL_168;
  assign fixer__EVAL_71 = system_bus_xbar__EVAL_65;
  assign _EVAL_202 = _EVAL_22;
  assign coupler_from_tile__EVAL_19 = _EVAL_52;
  assign _EVAL_142 = _EVAL_230;
  assign _EVAL_254 = _EVAL_236;
  assign system_bus_xbar__EVAL_87 = _EVAL_158;
  assign _EVAL_271 = _EVAL_212;
  assign _EVAL_289 = _EVAL_149;
  assign _EVAL_100 = _EVAL_291;
  assign system_bus_xbar__EVAL_80 = _EVAL_144;
  assign system_bus_xbar__EVAL_9 = fixer__EVAL_28;
  assign system_bus_xbar__EVAL_72 = _EVAL_184;
  assign _EVAL_333 = _EVAL_277;
  assign _EVAL_263 = _EVAL_258;
  assign _EVAL_275 = _EVAL_250;
  assign coupler_to_port_named_ahb_sys_port__EVAL_22 = system_bus_xbar__EVAL_4;
  assign _EVAL_277 = _EVAL_163;
  assign _EVAL_305 = _EVAL_96;
  assign _EVAL_188 = _EVAL_203;
  assign coupler_from_tile__EVAL_12 = _EVAL_7;
  assign _EVAL_123 = _EVAL_136;
  assign _EVAL_172 = _EVAL_284;
  assign system_bus_xbar__EVAL_34 = coupler_to_port_named_ahb_sys_port__EVAL_31;
  assign system_bus_xbar__EVAL_26 = _EVAL_295;
  assign system_bus_xbar__EVAL_53 = coupler_to_port_named_ahb_sys_port__EVAL_27;
  assign _EVAL_196 = _EVAL_222;
  assign _EVAL = coupler_from_tile__EVAL_32;
  assign _EVAL_233 = _EVAL_9;
  assign fixer__EVAL_10 = system_bus_xbar__EVAL_92;
  assign coupler_from_tile__EVAL_18 = fixedClockNode__EVAL;
  assign _EVAL_198 = system_bus_xbar__EVAL_79;
  assign _EVAL_191 = _EVAL_127;
  assign coupler_to_port_named_ahb_sys_port__EVAL_1 = _EVAL_37;
  assign coupler_from_tile__EVAL_3 = _EVAL_109;
  assign fixer__EVAL_24 = _EVAL_129;
  assign fixer__EVAL_75 = fixedClockNode__EVAL_0;
  assign fixer__EVAL_21 = system_bus_xbar__EVAL_49;
  assign _EVAL_274 = _EVAL_92;
  assign coupler_from_tile__EVAL_37 = fixer__EVAL_33;
  assign _EVAL_77 = coupler_from_tile__EVAL_6;
  assign fixer__EVAL_43 = system_bus_xbar__EVAL_37;
  assign _EVAL_151 = _EVAL_237;
  assign fixer__EVAL_53 = system_bus_xbar__EVAL_73;
  assign _EVAL_329 = _EVAL_273;
  assign _EVAL_32 = coupler_from_tile__EVAL_39;
  assign coupler_to_port_named_ahb_sys_port__EVAL_24 = system_bus_xbar__EVAL_63;
  assign _EVAL_291 = _EVAL_323;
  assign _EVAL_119 = _EVAL_174;
  assign _EVAL_17 = coupler_from_tile__EVAL_55;
endmodule
