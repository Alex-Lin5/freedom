//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_47_assert(
  input         _EVAL,
  input  [3:0]  _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input  [1:0]  _EVAL_4,
  input  [3:0]  _EVAL_5,
  input  [4:0]  _EVAL_6,
  input  [2:0]  _EVAL_7,
  input         _EVAL_8,
  input  [4:0]  _EVAL_9,
  input  [3:0]  _EVAL_10,
  input  [2:0]  _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input  [2:0]  _EVAL_16,
  input         _EVAL_17,
  input  [31:0] _EVAL_18
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  reg [5:0] _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire [31:0] _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire [1:0] _EVAL_37;
  wire  _EVAL_38;
  wire [5:0] _EVAL_39;
  wire  _EVAL_40;
  wire [31:0] _EVAL_41;
  wire [32:0] _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire [3:0] _EVAL_54;
  wire [2:0] _EVAL_55;
  reg [2:0] _EVAL_56;
  wire  _EVAL_57;
  reg [1:0] _EVAL_58;
  wire [6:0] _EVAL_59;
  wire [32:0] _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire [32:0] _EVAL_68;
  wire [3:0] _EVAL_69;
  wire [32:0] _EVAL_70;
  wire [31:0] _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire [7:0] _EVAL_79;
  wire  _EVAL_81;
  wire [32:0] _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire [32:0] _EVAL_85;
  wire [31:0] _EVAL_86;
  wire  _EVAL_87;
  wire [32:0] _EVAL_88;
  wire  _EVAL_89;
  wire [5:0] _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire [31:0] _EVAL_96;
  wire [17:0] _EVAL_97;
  wire [32:0] _EVAL_98;
  wire [17:0] _EVAL_99;
  wire  _EVAL_100;
  wire [7:0] _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  reg [5:0] _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_108;
  wire [5:0] _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  reg [3:0] _EVAL_124;
  reg  _EVAL_125;
  wire [1:0] _EVAL_126;
  wire [32:0] _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire [32:0] _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_136;
  wire [32:0] _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire [31:0] _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire [6:0] _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  reg  _EVAL_168;
  wire [32:0] _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  reg [31:0] _EVAL_174;
  wire [32:0] _EVAL_175;
  wire [6:0] _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire [7:0] _EVAL_185;
  wire [31:0] _EVAL_186;
  wire [1:0] _EVAL_187;
  reg [3:0] _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire [32:0] _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire [3:0] _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  reg [2:0] _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire [22:0] _EVAL_209;
  wire [17:0] _EVAL_210;
  wire [22:0] _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_216;
  reg [4:0] _EVAL_217;
  wire  _EVAL_218;
  wire [31:0] _EVAL_219;
  wire [5:0] _EVAL_220;
  wire [31:0] _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire [31:0] _EVAL_226;
  wire [2:0] _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire [32:0] _EVAL_232;
  wire  _EVAL_233;
  wire [3:0] _EVAL_234;
  wire  _EVAL_235;
  reg [4:0] _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire [32:0] _EVAL_239;
  wire [17:0] _EVAL_240;
  reg [5:0] _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire [5:0] _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire [31:0] _EVAL_266;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire [32:0] _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire [5:0] _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire [17:0] _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire  _EVAL_293;
  reg [5:0] _EVAL_294;
  wire  _EVAL_295;
  wire [32:0] _EVAL_296;
  wire  _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire [7:0] _EVAL_301;
  wire  _EVAL_302;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_307;
  wire [32:0] _EVAL_308;
  wire [17:0] _EVAL_309;
  wire  _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_317;
  wire [32:0] _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_320;
  wire  _EVAL_321;
  wire  _EVAL_322;
  wire  _EVAL_323;
  wire  _EVAL_324;
  wire  _EVAL_325;
  wire  _EVAL_326;
  wire  _EVAL_327;
  wire  _EVAL_328;
  wire [31:0] _EVAL_329;
  wire [32:0] _EVAL_330;
  wire  _EVAL_331;
  wire  _EVAL_332;
  wire  _EVAL_333;
  wire [31:0] _EVAL_334;
  reg [17:0] _EVAL_335;
  wire  _EVAL_336;
  wire  _EVAL_337;
  wire  _EVAL_338;
  wire  _EVAL_339;
  wire  _EVAL_340;
  wire  _EVAL_341;
  wire  _EVAL_342;
  wire  _EVAL_343;
  wire  _EVAL_344;
  wire [6:0] _EVAL_345;
  wire  _EVAL_346;
  wire  _EVAL_347;
  wire  _EVAL_348;
  wire  _EVAL_349;
  wire  _EVAL_350;
  wire  _EVAL_351;
  wire  _EVAL_352;
  wire  _EVAL_353;
  wire [1:0] _EVAL_354;
  wire [32:0] _EVAL_355;
  wire  _EVAL_356;
  wire  _EVAL_357;
  wire  _EVAL_358;
  wire  _EVAL_359;
  wire [17:0] _EVAL_360;
  wire  _EVAL_361;
  wire  _EVAL_362;
  reg [2:0] _EVAL_363;
  wire  _EVAL_364;
  wire  _EVAL_365;
  wire  _EVAL_366;
  wire  _EVAL_367;
  wire  _EVAL_368;
  wire  _EVAL_369;
  wire [17:0] _EVAL_370;
  wire  _EVAL_371;
  reg [31:0] _EVAL_372;
  wire  _EVAL_373;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_35 = ~_EVAL_328;
  assign _EVAL_258 = ~_EVAL_208;
  assign _EVAL_76 = _EVAL_9 == _EVAL_217;
  assign _EVAL_162 = _EVAL_7 == 3'h6;
  assign _EVAL_71 = _EVAL_139 ? _EVAL_41 : 32'h0;
  assign _EVAL_40 = ~_EVAL_264;
  assign _EVAL_117 = _EVAL_360 != _EVAL_370;
  assign _EVAL_295 = _EVAL_263 & _EVAL_323;
  assign _EVAL_134 = _EVAL_253 | _EVAL_274;
  assign _EVAL_201 = ~_EVAL_69;
  assign _EVAL_284 = _EVAL_10 <= 4'h6;
  assign _EVAL_150 = ~_EVAL_3;
  assign _EVAL_166 = ~_EVAL_21;
  assign _EVAL_83 = _EVAL_349 | _EVAL_3;
  assign _EVAL_127 = _EVAL_131;
  assign _EVAL_28 = _EVAL_165 & _EVAL_81;
  assign _EVAL_193 = _EVAL_373 | _EVAL_3;
  assign _EVAL_119 = _EVAL_18 == _EVAL_174;
  assign _EVAL_242 = _EVAL_14 & _EVAL_328;
  assign _EVAL_229 = _EVAL_16 == 3'h2;
  assign _EVAL_31 = _EVAL_65 | _EVAL_3;
  assign _EVAL_63 = _EVAL_7 == 3'h1;
  assign _EVAL_208 = _EVAL_89 | _EVAL_3;
  assign _EVAL_367 = _EVAL_113 | _EVAL_279;
  assign _EVAL_186 = 32'h1 << _EVAL_9;
  assign _EVAL_308 = $signed(_EVAL_296) & -33'sh2000;
  assign _EVAL_120 = _EVAL_7 == 3'h3;
  assign _EVAL_200 = ~_EVAL_172;
  assign _EVAL_70 = _EVAL_330;
  assign _EVAL_271 = $signed(_EVAL_98) == 33'sh0;
  assign _EVAL_274 = _EVAL_263 & _EVAL_132;
  assign _EVAL_276 = _EVAL_312 | _EVAL_3;
  assign _EVAL_329 = _EVAL_355[31:0];
  assign _EVAL_87 = _EVAL_149 | _EVAL_3;
  assign _EVAL_197 = $signed(_EVAL_239) & -33'sh10000;
  assign _EVAL_354 = _EVAL_126 | 2'h1;
  assign _EVAL_43 = ~_EVAL_95;
  assign _EVAL_116 = _EVAL_112 | _EVAL_271;
  assign _EVAL_179 = _EVAL_141 | _EVAL_224;
  assign _EVAL_85 = {1'b0,$signed(_EVAL_86)};
  assign _EVAL_257 = _EVAL_11 == 3'h0;
  assign _EVAL_285 = _EVAL_228 | _EVAL_24;
  assign _EVAL_131 = $signed(_EVAL_137) & -33'sh400000;
  assign _EVAL_317 = _EVAL_44 | _EVAL_3;
  assign _EVAL_350 = _EVAL_245 | _EVAL_2;
  assign _EVAL_111 = _EVAL_0 == _EVAL_69;
  assign _EVAL_245 = ~_EVAL_13;
  assign _EVAL_336 = ~_EVAL_152;
  assign _EVAL_314 = ~_EVAL_290;
  assign _EVAL_53 = _EVAL_372 < plusarg_reader_out;
  assign _EVAL_61 = $signed(_EVAL_318) & -33'sh5000;
  assign _EVAL_145 = _EVAL_117 | _EVAL_314;
  assign _EVAL_289 = _EVAL_304 | _EVAL_3;
  assign _EVAL_280 = _EVAL_259 & _EVAL_272;
  assign _EVAL_187 = _EVAL_9[4:3];
  assign _EVAL_260 = _EVAL_183 | _EVAL_3;
  assign _EVAL_33 = _EVAL_248 | _EVAL_3;
  assign _EVAL_172 = _EVAL_265 | _EVAL_3;
  assign _EVAL_170 = _EVAL_362 & _EVAL_36;
  assign _EVAL_287 = _EVAL_231 | _EVAL_224;
  assign _EVAL_49 = _EVAL_230 | _EVAL_3;
  assign _EVAL_81 = _EVAL_9 == 5'h8;
  assign _EVAL_297 = _EVAL_294 == 6'h0;
  assign _EVAL_204 = _EVAL_173 & _EVAL_128;
  assign _EVAL_306 = ~_EVAL_147;
  assign _EVAL_270 = _EVAL_232;
  assign _EVAL_151 = _EVAL_7 == 3'h7;
  assign _EVAL_181 = ~_EVAL_31;
  assign _EVAL_338 = _EVAL_142 | _EVAL_3;
  assign _EVAL_332 = _EVAL_106 | _EVAL_3;
  assign _EVAL_348 = _EVAL_263 & _EVAL_32;
  assign _EVAL_356 = ~_EVAL_156;
  assign _EVAL_194 = ~_EVAL_268;
  assign _EVAL_298 = _EVAL_6 == 5'h10;
  assign _EVAL_263 = _EVAL_354[0];
  assign _EVAL_161 = _EVAL_11 <= 3'h4;
  assign _EVAL_207 = ~_EVAL_315;
  assign _EVAL_133 = _EVAL_6 == 5'h11;
  assign _EVAL_114 = _EVAL_259 | _EVAL_362;
  assign _EVAL_54 = _EVAL_0 & _EVAL_201;
  assign _EVAL_115 = _EVAL_234 == 4'h0;
  assign _EVAL_359 = ~_EVAL_282;
  assign _EVAL_315 = _EVAL_76 | _EVAL_3;
  assign _EVAL_357 = $signed(_EVAL_70) == 33'sh0;
  assign _EVAL_138 = _EVAL_6 == _EVAL_236;
  assign _EVAL_366 = ~_EVAL_278;
  assign _EVAL_159 = ~_EVAL_223;
  assign _EVAL_165 = 4'h6 == _EVAL_10;
  assign _EVAL_296 = {1'b0,$signed(_EVAL_334)};
  assign _EVAL_256 = _EVAL_115 | _EVAL_3;
  assign _EVAL_320 = ~_EVAL_347;
  assign _EVAL_153 = _EVAL_253 | _EVAL_108;
  assign _EVAL_246 = _EVAL_10[0];
  assign _EVAL_278 = _EVAL_257 | _EVAL_3;
  assign _EVAL_213 = _EVAL_17 & _EVAL_341;
  assign _EVAL_36 = _EVAL_29 == 6'h0;
  assign _EVAL_156 = _EVAL_350 | _EVAL_3;
  assign _EVAL_301 = ~_EVAL_185;
  assign _EVAL_288 = _EVAL_7 == 3'h4;
  assign _EVAL_152 = _EVAL_145 | _EVAL_3;
  assign _EVAL_72 = ~_EVAL_317;
  assign _EVAL_50 = _EVAL_14 & _EVAL_84;
  assign _EVAL_291 = _EVAL_17 & _EVAL_288;
  assign _EVAL_259 = _EVAL & _EVAL_17;
  assign _EVAL_371 = _EVAL_259 & _EVAL_297;
  assign _EVAL_91 = _EVAL_7 == 3'h5;
  assign _EVAL_34 = _EVAL_18 & _EVAL_266;
  assign _EVAL_344 = ~_EVAL_49;
  assign _EVAL_325 = ~_EVAL_346;
  assign _EVAL_24 = _EVAL_6 == 5'h8;
  assign _EVAL_94 = ~_EVAL_256;
  assign _EVAL_126 = 2'h1 << _EVAL_246;
  assign _EVAL_218 = ~_EVAL_171;
  assign _EVAL_290 = |_EVAL_360;
  assign _EVAL_243 = _EVAL_225 | _EVAL_3;
  assign _EVAL_48 = _EVAL_265 | _EVAL_343;
  assign _EVAL_292 = _EVAL_269 | _EVAL_3;
  assign _EVAL_78 = _EVAL_284 & _EVAL_238;
  assign _EVAL_106 = _EVAL_113 | _EVAL_337;
  assign _EVAL_328 = _EVAL_16 == 3'h6;
  assign _EVAL_305 = _EVAL_367 | _EVAL_3;
  assign _EVAL_97 = _EVAL_335 | _EVAL_360;
  assign _EVAL_349 = _EVAL_160 | _EVAL_28;
  assign _EVAL_74 = _EVAL_48 | _EVAL_348;
  assign _EVAL_198 = _EVAL_7 == 3'h2;
  assign _EVAL_203 = $signed(_EVAL_88) == 33'sh0;
  assign _EVAL_122 = ~_EVAL_243;
  assign _EVAL_324 = _EVAL_48 | _EVAL_295;
  assign _EVAL_307 = ~_EVAL_338;
  assign _EVAL_148 = ~_EVAL_100;
  assign _EVAL_22 = _EVAL_368 | _EVAL_167;
  assign _EVAL_219 = _EVAL_18 ^ 32'h1800000;
  assign _EVAL_211 = 23'hff << _EVAL_10;
  assign _EVAL_209 = 23'hff << _EVAL_5;
  assign _EVAL_265 = _EVAL_10 >= 4'h2;
  assign _EVAL_139 = _EVAL_170 & _EVAL_35;
  assign _EVAL_79 = ~_EVAL_101;
  assign _EVAL_237 = ~_EVAL_2;
  assign _EVAL_157 = _EVAL_299 | _EVAL_3;
  assign _EVAL_93 = _EVAL_4 != 2'h2;
  assign _EVAL_239 = {1'b0,$signed(_EVAL_143)};
  assign _EVAL_269 = _EVAL_13 == _EVAL_168;
  assign _EVAL_95 = _EVAL_119 | _EVAL_3;
  assign _EVAL_44 = _EVAL_10 == _EVAL_124;
  assign _EVAL_184 = ~_EVAL_189;
  assign _EVAL_137 = {1'b0,$signed(_EVAL_226)};
  assign _EVAL_309 = _EVAL_97 & _EVAL_99;
  assign _EVAL_96 = _EVAL_371 ? _EVAL_186 : 32'h0;
  assign _EVAL_123 = _EVAL_17 & _EVAL_63;
  assign _EVAL_226 = _EVAL_18 ^ 32'hc000000;
  assign _EVAL_46 = _EVAL_54 == 4'h0;
  assign _EVAL_129 = _EVAL_15 == _EVAL_125;
  assign _EVAL_346 = _EVAL_46 | _EVAL_3;
  assign _EVAL_154 = ~_EVAL_33;
  assign _EVAL_177 = _EVAL_75 | _EVAL_3;
  assign _EVAL_220 = _EVAL_301[7:2];
  assign _EVAL_130 = _EVAL_16 == 3'h4;
  assign _EVAL_345 = _EVAL_29 - 6'h1;
  assign _EVAL_244 = ~_EVAL_77;
  assign _EVAL_277 = ~_EVAL_365;
  assign _EVAL_191 = _EVAL_7[2];
  assign _EVAL_227 = _EVAL_6[2:0];
  assign _EVAL_169 = {1'b0,$signed(_EVAL_221)};
  assign _EVAL_68 = _EVAL_308;
  assign _EVAL_281 = _EVAL_182 & _EVAL_287;
  assign _EVAL_66 = _EVAL_326 & _EVAL_358;
  assign _EVAL_196 = _EVAL_195 | _EVAL_238;
  assign _EVAL_272 = _EVAL_104 == 6'h0;
  assign _EVAL_51 = _EVAL_241 == 6'h0;
  assign _EVAL_254 = _EVAL_17 & _EVAL_91;
  assign _EVAL_248 = _EVAL_7 == _EVAL_206;
  assign _EVAL_279 = _EVAL_284 & _EVAL_102;
  assign _EVAL_59 = _EVAL_104 - 6'h1;
  assign _EVAL_132 = _EVAL_247 & _EVAL_184;
  assign _EVAL_75 = _EVAL_113 | _EVAL_78;
  assign _EVAL_282 = _EVAL_111 | _EVAL_3;
  assign _EVAL_27 = ~_EVAL_19;
  assign _EVAL_110 = _EVAL_14 & _EVAL_361;
  assign _EVAL_266 = {{24'd0}, _EVAL_301};
  assign _EVAL_45 = $signed(_EVAL_270) == 33'sh0;
  assign _EVAL_176 = _EVAL_294 - 6'h1;
  assign _EVAL_146 = ~_EVAL_164;
  assign _EVAL_223 = _EVAL_364 | _EVAL_3;
  assign _EVAL_113 = _EVAL_327 & _EVAL_357;
  assign _EVAL_261 = _EVAL_17 & _EVAL_162;
  assign _EVAL_109 = _EVAL_176[5:0];
  assign _EVAL_163 = _EVAL_17 & _EVAL_120;
  assign _EVAL_128 = _EVAL_9 == 5'h10;
  assign _EVAL_142 = ~_EVAL_331;
  assign _EVAL_234 = ~_EVAL_0;
  assign _EVAL_318 = {1'b0,$signed(_EVAL_18)};
  assign _EVAL_339 = ~_EVAL_8;
  assign _EVAL_47 = _EVAL_14 & _EVAL_130;
  assign _EVAL_67 = _EVAL_4 == _EVAL_58;
  assign _EVAL_250 = _EVAL_362 & _EVAL_51;
  assign _EVAL_311 = _EVAL_16 == 3'h0;
  assign _EVAL_351 = ~_EVAL_276;
  assign _EVAL_102 = _EVAL_196 | _EVAL_45;
  assign _EVAL_321 = _EVAL_17 & _EVAL_151;
  assign _EVAL_369 = ~_EVAL_247;
  assign _EVAL_210 = _EVAL_335 >> _EVAL_9;
  assign _EVAL_147 = _EVAL_93 | _EVAL_3;
  assign _EVAL_57 = _EVAL_187 == 2'h0;
  assign _EVAL_327 = _EVAL_10 <= 4'h8;
  assign _EVAL_190 = ~_EVAL_191;
  assign _EVAL_20 = ~_EVAL_87;
  assign _EVAL_52 = _EVAL_262 | _EVAL_233;
  assign _EVAL_316 = _EVAL_354[1];
  assign _EVAL_240 = _EVAL_286 >> _EVAL_6;
  assign _EVAL_173 = _EVAL_10 <= 4'hb;
  assign _EVAL_105 = _EVAL_5 >= 4'h2;
  assign _EVAL_77 = _EVAL_138 | _EVAL_3;
  assign _EVAL_247 = _EVAL_18[1];
  assign _EVAL_362 = _EVAL_12 & _EVAL_14;
  assign _EVAL_141 = _EVAL_231 | _EVAL_128;
  assign _EVAL_185 = _EVAL_211[7:0];
  assign _EVAL_99 = ~_EVAL_370;
  assign _EVAL_253 = _EVAL_265 | _EVAL_313;
  assign _EVAL_180 = ~_EVAL_352;
  assign _EVAL_230 = _EVAL_5 == _EVAL_188;
  assign _EVAL_69 = {_EVAL_153,_EVAL_134,_EVAL_324,_EVAL_74};
  assign _EVAL_331 = _EVAL_210[0];
  assign _EVAL_360 = _EVAL_96[17:0];
  assign _EVAL_25 = _EVAL_199 & _EVAL_224;
  assign _EVAL_101 = _EVAL_209[7:0];
  assign _EVAL_238 = $signed(_EVAL_68) == 33'sh0;
  assign _EVAL_214 = ~_EVAL_305;
  assign _EVAL_268 = _EVAL_339 | _EVAL_3;
  assign _EVAL_182 = _EVAL_10 <= 4'h2;
  assign _EVAL_340 = _EVAL_11 <= 3'h1;
  assign _EVAL_160 = _EVAL_281 | _EVAL_204;
  assign _EVAL_65 = _EVAL_4 == 2'h0;
  assign _EVAL_149 = _EVAL_25 & _EVAL_22;
  assign _EVAL_313 = _EVAL_316 & _EVAL_247;
  assign _EVAL_38 = _EVAL_17 & _EVAL_198;
  assign _EVAL_19 = _EVAL_105 | _EVAL_3;
  assign _EVAL_283 = _EVAL_133 | _EVAL_298;
  assign _EVAL_221 = _EVAL_18 ^ 32'h80000000;
  assign _EVAL_361 = _EVAL_16 == 3'h1;
  assign _EVAL_264 = _EVAL_293 | _EVAL_3;
  assign _EVAL_255 = $signed(_EVAL_127) == 33'sh0;
  assign _EVAL_37 = _EVAL_6[4:3];
  assign _EVAL_262 = ~_EVAL_64;
  assign _EVAL_216 = ~_EVAL_157;
  assign _EVAL_30 = ~_EVAL_51;
  assign _EVAL_144 = _EVAL_11 <= 3'h2;
  assign _EVAL_171 = _EVAL_285 | _EVAL_3;
  assign _EVAL_373 = _EVAL_16 == _EVAL_363;
  assign _EVAL_337 = _EVAL_284 & _EVAL_92;
  assign _EVAL_326 = _EVAL_37 == 2'h0;
  assign _EVAL_175 = $signed(_EVAL_42) & -33'sh4000;
  assign _EVAL_232 = $signed(_EVAL_169) & -33'sh4000;
  assign _EVAL_167 = _EVAL_199 & _EVAL_45;
  assign _EVAL_158 = _EVAL_245 | _EVAL_3;
  assign _EVAL_222 = _EVAL_4 <= 2'h2;
  assign _EVAL_92 = _EVAL_195 | _EVAL_45;
  assign _EVAL_224 = _EVAL_57 & _EVAL_342;
  assign _EVAL_273 = _EVAL_237 | _EVAL_3;
  assign _EVAL_42 = {1'b0,$signed(_EVAL_219)};
  assign _EVAL_343 = _EVAL_316 & _EVAL_369;
  assign _EVAL_286 = _EVAL_360 | _EVAL_335;
  assign _EVAL_26 = ~_EVAL_260;
  assign _EVAL_88 = _EVAL_175;
  assign _EVAL_319 = _EVAL_160 & _EVAL_367;
  assign _EVAL_333 = ~_EVAL_193;
  assign _EVAL_205 = _EVAL_17 & _EVAL_23;
  assign _EVAL_32 = _EVAL_369 & _EVAL_184;
  assign _EVAL_293 = _EVAL_16 <= 3'h6;
  assign _EVAL_358 = _EVAL_227 <= 3'h6;
  assign _EVAL_312 = _EVAL_11 == _EVAL_56;
  assign _EVAL_235 = $signed(_EVAL_82) == 33'sh0;
  assign _EVAL_355 = _EVAL_372 + 32'h1;
  assign _EVAL_368 = _EVAL_182 & _EVAL_357;
  assign _EVAL_103 = _EVAL_247 & _EVAL_189;
  assign _EVAL_86 = _EVAL_18 ^ 32'h3000;
  assign _EVAL_136 = ~_EVAL_332;
  assign _EVAL_108 = _EVAL_263 & _EVAL_103;
  assign _EVAL_121 = _EVAL_14 & _EVAL_229;
  assign _EVAL_90 = _EVAL_79[7:2];
  assign _EVAL_189 = _EVAL_18[0];
  assign _EVAL_370 = _EVAL_71[17:0];
  assign _EVAL_334 = _EVAL_18 ^ 32'h20000000;
  assign _EVAL_89 = _EVAL_34 == 32'h0;
  assign _EVAL_23 = _EVAL_7 == 3'h0;
  assign _EVAL_252 = _EVAL_319 | _EVAL_3;
  assign _EVAL_300 = ~_EVAL_289;
  assign _EVAL_202 = _EVAL_16[0];
  assign _EVAL_164 = _EVAL_67 | _EVAL_3;
  assign _EVAL_55 = _EVAL_9[2:0];
  assign _EVAL_341 = ~_EVAL_272;
  assign _EVAL_275 = _EVAL_345[5:0];
  assign _EVAL_352 = _EVAL_161 | _EVAL_3;
  assign _EVAL_155 = _EVAL_241 - 6'h1;
  assign _EVAL_365 = _EVAL_144 | _EVAL_3;
  assign _EVAL_330 = $signed(_EVAL_85) & -33'sh1000;
  assign _EVAL_39 = _EVAL_59[5:0];
  assign _EVAL_231 = _EVAL_9 == 5'h11;
  assign _EVAL_249 = ~_EVAL_83;
  assign _EVAL_225 = _EVAL_240[0];
  assign _EVAL_251 = _EVAL_155[5:0];
  assign _EVAL_98 = _EVAL_197;
  assign _EVAL_64 = |_EVAL_335;
  assign _EVAL_84 = _EVAL_16 == 3'h5;
  assign _EVAL_199 = 4'h2 == _EVAL_10;
  assign _EVAL_62 = ~_EVAL_273;
  assign _EVAL_192 = ~_EVAL_158;
  assign _EVAL_183 = _EVAL_11 != 3'h0;
  assign _EVAL_178 = ~_EVAL_292;
  assign _EVAL_322 = ~_EVAL_252;
  assign _EVAL_302 = _EVAL_14 & _EVAL_30;
  assign _EVAL_353 = ~_EVAL_177;
  assign _EVAL_100 = _EVAL_129 | _EVAL_3;
  assign _EVAL_143 = _EVAL_18 ^ 32'h2000000;
  assign _EVAL_304 = _EVAL_52 | _EVAL_53;
  assign _EVAL_323 = _EVAL_369 & _EVAL_189;
  assign _EVAL_342 = _EVAL_55 <= 3'h6;
  assign _EVAL_41 = 32'h1 << _EVAL_6;
  assign _EVAL_364 = _EVAL_11 <= 3'h3;
  assign _EVAL_82 = _EVAL_61;
  assign _EVAL_212 = _EVAL_14 & _EVAL_311;
  assign _EVAL_112 = _EVAL_235 | _EVAL_203;
  assign _EVAL_21 = _EVAL_222 | _EVAL_3;
  assign _EVAL_299 = _EVAL_179 | _EVAL_81;
  assign _EVAL_228 = _EVAL_283 | _EVAL_66;
  assign _EVAL_233 = plusarg_reader_out == 32'h0;
  assign _EVAL_347 = _EVAL_340 | _EVAL_3;
  assign _EVAL_195 = _EVAL_116 | _EVAL_255;
  always @(posedge _EVAL_1) begin
    if (_EVAL_3) begin
      _EVAL_29 <= 6'h0;
    end else if (_EVAL_362) begin
      if (_EVAL_36) begin
        if (_EVAL_202) begin
          _EVAL_29 <= _EVAL_90;
        end else begin
          _EVAL_29 <= 6'h0;
        end
      end else begin
        _EVAL_29 <= _EVAL_275;
      end
    end
    if (_EVAL_280) begin
      _EVAL_56 <= _EVAL_11;
    end
    if (_EVAL_250) begin
      _EVAL_58 <= _EVAL_4;
    end
    if (_EVAL_3) begin
      _EVAL_104 <= 6'h0;
    end else if (_EVAL_259) begin
      if (_EVAL_272) begin
        if (_EVAL_190) begin
          _EVAL_104 <= _EVAL_220;
        end else begin
          _EVAL_104 <= 6'h0;
        end
      end else begin
        _EVAL_104 <= _EVAL_39;
      end
    end
    if (_EVAL_280) begin
      _EVAL_124 <= _EVAL_10;
    end
    if (_EVAL_250) begin
      _EVAL_125 <= _EVAL_15;
    end
    if (_EVAL_250) begin
      _EVAL_168 <= _EVAL_13;
    end
    if (_EVAL_280) begin
      _EVAL_174 <= _EVAL_18;
    end
    if (_EVAL_250) begin
      _EVAL_188 <= _EVAL_5;
    end
    if (_EVAL_280) begin
      _EVAL_206 <= _EVAL_7;
    end
    if (_EVAL_280) begin
      _EVAL_217 <= _EVAL_9;
    end
    if (_EVAL_250) begin
      _EVAL_236 <= _EVAL_6;
    end
    if (_EVAL_3) begin
      _EVAL_241 <= 6'h0;
    end else if (_EVAL_362) begin
      if (_EVAL_51) begin
        if (_EVAL_202) begin
          _EVAL_241 <= _EVAL_90;
        end else begin
          _EVAL_241 <= 6'h0;
        end
      end else begin
        _EVAL_241 <= _EVAL_251;
      end
    end
    if (_EVAL_3) begin
      _EVAL_294 <= 6'h0;
    end else if (_EVAL_259) begin
      if (_EVAL_297) begin
        if (_EVAL_190) begin
          _EVAL_294 <= _EVAL_220;
        end else begin
          _EVAL_294 <= 6'h0;
        end
      end else begin
        _EVAL_294 <= _EVAL_109;
      end
    end
    if (_EVAL_3) begin
      _EVAL_335 <= 18'h0;
    end else begin
      _EVAL_335 <= _EVAL_309;
    end
    if (_EVAL_250) begin
      _EVAL_363 <= _EVAL_16;
    end
    if (_EVAL_3) begin
      _EVAL_372 <= 32'h0;
    end else if (_EVAL_114) begin
      _EVAL_372 <= 32'h0;
    end else begin
      _EVAL_372 <= _EVAL_329;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46353ac4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32624eed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_322) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_371 & _EVAL_307) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(adebe008)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad837126)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f501b17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_366) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16f594af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(988a597f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1d7b640)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5dd203fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_356) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(680ce53d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_359) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_320) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_178) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4e995f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(922678c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c99bf1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f445a0d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_306) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e396478e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(224dbd32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_300) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(668dbb3d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30ece8c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_72) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_336) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc7dfa10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5188eac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_359) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77a5a25c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7117802f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6fb30f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(272879)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_366) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_325) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92d59f13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0d81f74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c14497c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ba6f7cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_351) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca7ee25f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_333) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_159) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75694818)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31b39aa7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea3dae63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_356) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_40) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3dd6630)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_366) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d20bbb87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(549e9f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_333) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f4c39ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c37d274a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_194) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_300) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_359) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94dd3707)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_249) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_366) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6caa6195)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_359) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60a052aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_122) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75560b1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(426e6ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17715120)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62e4a3db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_249) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce9f7766)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_181) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a40117d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_366) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cb36bb4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_344) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_366) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af08b89f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(861e703c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_359) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90930dfb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_258) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_344) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81201ba8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74de1520)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_178) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(109414ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aefde60e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d8380a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_359) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_136) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1308d567)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac0662c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_356) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd0293b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_14 & _EVAL_40) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cf770e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_306) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c064038c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af08b89f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_136) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_216) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(453aeb3d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e30cf63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_180) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_159) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f94919df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_306) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_322) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf709a17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ea84539)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_242 & _EVAL_181) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec7e6dec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8a94925)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_351) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_72) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(563a07eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_325) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98fd4b0d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9e64164)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5b2d4fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_302 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(786bdba8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_150) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_180) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4dd3305)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6240e7f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b457055b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_359) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b741c31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_122) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_216) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88c949c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_371 & _EVAL_307) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25014a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_150) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8fda73ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_110 & _EVAL_356) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5b66e48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_121 & _EVAL_218) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8cf403b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_163 & _EVAL_359) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e5dc540)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d06ea7f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(daf0a20a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_320) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eaae7d68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_336) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_258) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(63c6f3e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86121022)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_212 & _EVAL_218) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_359) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_359) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9670559e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_47 & _EVAL_306) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee7760bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_353) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0748023)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f46d359a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_254 & _EVAL_353) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_213 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eebb5832)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_321 & _EVAL_194) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28fb892c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_29 = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_56 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_58 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_104 = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_124 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_125 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_168 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_174 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_188 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_206 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_217 = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_236 = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_241 = _RAND_12[5:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_294 = _RAND_13[5:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_335 = _RAND_14[17:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_363 = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_372 = _RAND_16[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
