//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_60_assert(
  input  [4:0]  _EVAL,
  input         _EVAL_0,
  input  [2:0]  _EVAL_1,
  input         _EVAL_2,
  input  [27:0] _EVAL_3,
  input  [2:0]  _EVAL_4,
  input         _EVAL_5,
  input  [2:0]  _EVAL_6,
  input  [4:0]  _EVAL_7,
  input  [2:0]  _EVAL_8,
  input         _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input  [3:0]  _EVAL_13,
  input  [2:0]  _EVAL_14
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire [4:0] _EVAL_15;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire [31:0] _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  reg [2:0] _EVAL_25;
  wire  _EVAL_27;
  reg [2:0] _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  reg [27:0] _EVAL_35;
  wire [17:0] _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire [5:0] _EVAL_42;
  wire [1:0] _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire [17:0] _EVAL_48;
  wire [3:0] _EVAL_49;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire [12:0] _EVAL_56;
  wire [3:0] _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire [17:0] _EVAL_60;
  wire [32:0] _EVAL_61;
  wire [28:0] _EVAL_62;
  wire [2:0] _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire [3:0] _EVAL_67;
  wire [17:0] _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire [3:0] _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  reg [2:0] _EVAL_79;
  wire [3:0] _EVAL_80;
  wire  _EVAL_81;
  wire [27:0] _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire [1:0] _EVAL_88;
  wire [5:0] _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire [5:0] _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire [31:0] _EVAL_103;
  wire  _EVAL_104;
  wire [28:0] _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire [4:0] _EVAL_109;
  wire  _EVAL_110;
  wire [27:0] _EVAL_111;
  wire  _EVAL_112;
  wire [3:0] _EVAL_113;
  wire [31:0] _EVAL_114;
  wire  _EVAL_115;
  wire [27:0] _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire [17:0] _EVAL_119;
  wire [2:0] _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire [4:0] _EVAL_128;
  wire  _EVAL_129;
  wire [12:0] _EVAL_130;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  reg [2:0] _EVAL_145;
  wire  _EVAL_146;
  wire [3:0] _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire [4:0] _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire [3:0] _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire [17:0] _EVAL_171;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  reg [3:0] _EVAL_180;
  wire  _EVAL_181;
  reg [3:0] _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire [31:0] _EVAL_190;
  wire [5:0] _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire [1:0] _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  reg [4:0] _EVAL_208;
  wire  _EVAL_209;
  reg [4:0] _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire [31:0] _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  reg [3:0] _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire [1:0] _EVAL_238;
  wire  _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire [3:0] _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire [3:0] _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  reg [31:0] _EVAL_252;
  reg [2:0] _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire [17:0] _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire  _EVAL_261;
  reg [3:0] _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  reg [17:0] _EVAL_268;
  wire  _EVAL_269;
  wire [28:0] _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire [17:0] _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_177 = _EVAL_8 >= 3'h2;
  assign _EVAL_61 = _EVAL_252 + 32'h1;
  assign _EVAL_249 = _EVAL_1 == 3'h5;
  assign _EVAL_39 = ~_EVAL_276;
  assign _EVAL_272 = _EVAL_37 | _EVAL_85;
  assign _EVAL_276 = |_EVAL_268;
  assign _EVAL_188 = _EVAL_7 == 5'h10;
  assign _EVAL_103 = _EVAL_239 ? _EVAL_114 : 32'h0;
  assign _EVAL_57 = _EVAL_154[3:0];
  assign _EVAL_256 = _EVAL_143 | _EVAL_2;
  assign _EVAL_207 = _EVAL_10 & _EVAL_129;
  assign _EVAL_44 = _EVAL_10 & _EVAL_170;
  assign _EVAL_259 = _EVAL_13 == _EVAL_74;
  assign _EVAL_105 = _EVAL_62;
  assign _EVAL_282 = _EVAL_246 | _EVAL_99;
  assign _EVAL_178 = _EVAL_14[0];
  assign _EVAL_87 = _EVAL_139 & _EVAL_110;
  assign _EVAL_125 = _EVAL_225 == 4'h0;
  assign _EVAL_265 = _EVAL_3[1];
  assign _EVAL_227 = |_EVAL_36;
  assign _EVAL_222 = _EVAL_11 & _EVAL_149;
  assign _EVAL_245 = _EVAL_191[5:2];
  assign _EVAL_176 = _EVAL_228 & _EVAL_87;
  assign _EVAL_43 = 2'h1 << _EVAL_137;
  assign _EVAL_244 = _EVAL_4 == _EVAL_79;
  assign _EVAL_202 = _EVAL_182 == 4'h0;
  assign _EVAL_147 = _EVAL_92[5:2];
  assign _EVAL_206 = _EVAL_224 | _EVAL_140;
  assign _EVAL_120 = _EVAL_7[2:0];
  assign _EVAL_95 = _EVAL_262 == 4'h0;
  assign _EVAL_137 = _EVAL_4[0];
  assign _EVAL_144 = _EVAL_186 | _EVAL_2;
  assign _EVAL_254 = ~_EVAL_46;
  assign _EVAL_40 = _EVAL_201 & _EVAL_95;
  assign _EVAL_223 = _EVAL_10 & _EVAL_141;
  assign _EVAL_237 = ~_EVAL_211;
  assign _EVAL_31 = ~_EVAL_213;
  assign _EVAL_32 = _EVAL_121 | _EVAL_2;
  assign _EVAL_229 = _EVAL_219 | _EVAL_165;
  assign _EVAL_161 = _EVAL_6 <= 3'h2;
  assign _EVAL_195 = _EVAL_7 == 5'h11;
  assign _EVAL_109 = _EVAL_180 - 4'h1;
  assign _EVAL_193 = _EVAL_63 <= 3'h6;
  assign _EVAL_191 = ~_EVAL_42;
  assign _EVAL_146 = _EVAL_8 == _EVAL_25;
  assign _EVAL_37 = _EVAL_217 | _EVAL_281;
  assign _EVAL_127 = _EVAL_218 | _EVAL_2;
  assign _EVAL_218 = _EVAL_67 == 4'h0;
  assign _EVAL_126 = ~_EVAL_106;
  assign _EVAL_204 = _EVAL_1 == _EVAL_253;
  assign _EVAL_113 = _EVAL_109[3:0];
  assign _EVAL_119 = _EVAL_48 & _EVAL_273;
  assign _EVAL_250 = _EVAL_131 | _EVAL_2;
  assign _EVAL_139 = ~_EVAL_265;
  assign _EVAL_162 = _EVAL_1 == 3'h2;
  assign _EVAL_142 = ~_EVAL_77;
  assign _EVAL_98 = _EVAL_139 & _EVAL_45;
  assign _EVAL_102 = _EVAL_6 <= 3'h3;
  assign _EVAL_71 = _EVAL_14 == 3'h5;
  assign _EVAL_232 = _EVAL_194 | _EVAL_2;
  assign _EVAL_228 = _EVAL_238[0];
  assign _EVAL_117 = _EVAL_120 <= 3'h6;
  assign _EVAL_213 = _EVAL_264 | _EVAL_2;
  assign _EVAL_122 = _EVAL_14 == 3'h6;
  assign _EVAL_21 = _EVAL_40 ? _EVAL_190 : 32'h0;
  assign _EVAL_280 = ~_EVAL_65;
  assign _EVAL_269 = _EVAL_4 <= 3'h2;
  assign _EVAL_89 = _EVAL_56[5:0];
  assign _EVAL_136 = _EVAL == 5'h8;
  assign _EVAL_30 = _EVAL_3 == _EVAL_35;
  assign _EVAL_64 = _EVAL_6 <= 3'h1;
  assign _EVAL_99 = _EVAL_228 & _EVAL_23;
  assign _EVAL_114 = 32'h1 << _EVAL_7;
  assign _EVAL_74 = {_EVAL_240,_EVAL_282,_EVAL_53,_EVAL_138};
  assign _EVAL_80 = _EVAL_128[3:0];
  assign _EVAL_77 = _EVAL_164 | _EVAL_2;
  assign _EVAL_91 = _EVAL_4 <= 3'h6;
  assign _EVAL_75 = _EVAL_283 | _EVAL_2;
  assign _EVAL_134 = _EVAL_37 & _EVAL_216;
  assign _EVAL_16 = _EVAL_1 == 3'h0;
  assign _EVAL_216 = _EVAL_91 & _EVAL_151;
  assign _EVAL_101 = ~_EVAL_241;
  assign _EVAL_106 = _EVAL_214 | _EVAL_2;
  assign _EVAL_197 = _EVAL_7[4:3];
  assign _EVAL_278 = ~_EVAL_107;
  assign _EVAL_85 = _EVAL_169 & _EVAL_136;
  assign _EVAL_247 = _EVAL_229 | _EVAL_2;
  assign _EVAL_214 = _EVAL_6 != 3'h0;
  assign _EVAL_279 = ~_EVAL_261;
  assign _EVAL_56 = 13'h3f << _EVAL_4;
  assign _EVAL_219 = _EVAL_72 | _EVAL_184;
  assign _EVAL_107 = _EVAL_64 | _EVAL_2;
  assign _EVAL_15 = _EVAL_262 - 4'h1;
  assign _EVAL_261 = _EVAL_97 | _EVAL_2;
  assign _EVAL_94 = ~_EVAL_227;
  assign _EVAL_49 = ~_EVAL_74;
  assign _EVAL_264 = _EVAL == _EVAL_208;
  assign _EVAL_189 = _EVAL_197 == 2'h0;
  assign _EVAL_267 = _EVAL_7 == _EVAL_210;
  assign _EVAL_83 = ~_EVAL_55;
  assign _EVAL_184 = _EVAL_189 & _EVAL_117;
  assign _EVAL_168 = _EVAL_242 == 4'h0;
  assign _EVAL_185 = ~_EVAL_202;
  assign _EVAL_150 = _EVAL_274 & _EVAL_265;
  assign _EVAL_274 = _EVAL_238[1];
  assign _EVAL_248 = _EVAL_274 & _EVAL_139;
  assign _EVAL_233 = _EVAL_59 | _EVAL_2;
  assign _EVAL_88 = _EVAL[4:3];
  assign _EVAL_129 = _EVAL_14 == 3'h1;
  assign _EVAL_187 = ~_EVAL_32;
  assign _EVAL_73 = _EVAL_265 & _EVAL_45;
  assign _EVAL_217 = _EVAL_269 & _EVAL_206;
  assign _EVAL_246 = _EVAL_283 | _EVAL_150;
  assign _EVAL_255 = _EVAL_259 | _EVAL_2;
  assign _EVAL_121 = _EVAL_263 | _EVAL_199;
  assign _EVAL_63 = _EVAL[2:0];
  assign _EVAL_59 = ~_EVAL_9;
  assign _EVAL_108 = _EVAL_11 & _EVAL_152;
  assign _EVAL_221 = _EVAL_61[31:0];
  assign _EVAL_104 = _EVAL_148 | _EVAL_2;
  assign _EVAL_154 = _EVAL_225 - 4'h1;
  assign _EVAL_66 = _EVAL_201 & _EVAL_202;
  assign _EVAL_215 = _EVAL_180 == 4'h0;
  assign _EVAL_236 = _EVAL_11 & _EVAL_249;
  assign _EVAL_190 = 32'h1 << _EVAL;
  assign _EVAL_118 = _EVAL_5 & _EVAL_10;
  assign _EVAL_141 = _EVAL_14 == 3'h4;
  assign _EVAL_167 = _EVAL_36 != _EVAL_257;
  assign _EVAL_179 = ~_EVAL_212;
  assign _EVAL_65 = _EVAL_102 | _EVAL_2;
  assign _EVAL_23 = _EVAL_265 & _EVAL_110;
  assign _EVAL_152 = _EVAL_1 == 3'h4;
  assign _EVAL_93 = ~_EVAL_86;
  assign _EVAL_198 = _EVAL_96 | _EVAL_140;
  assign _EVAL_211 = _EVAL_30 | _EVAL_2;
  assign _EVAL_271 = ~_EVAL_255;
  assign _EVAL_148 = _EVAL_6 == _EVAL_145;
  assign _EVAL_58 = ~_EVAL_17;
  assign _EVAL_199 = _EVAL_252 < plusarg_reader_out;
  assign _EVAL_78 = _EVAL_11 & _EVAL_185;
  assign _EVAL_173 = ~_EVAL_250;
  assign _EVAL_67 = _EVAL_13 & _EVAL_49;
  assign _EVAL_156 = ~_EVAL_157;
  assign _EVAL_194 = _EVAL_167 | _EVAL_94;
  assign _EVAL_170 = ~_EVAL_125;
  assign _EVAL_239 = _EVAL_115 & _EVAL_54;
  assign _EVAL_135 = ~_EVAL_81;
  assign _EVAL_20 = ~_EVAL_256;
  assign _EVAL_166 = _EVAL_15[3:0];
  assign _EVAL_251 = _EVAL_177 | _EVAL_2;
  assign _EVAL_201 = _EVAL_0 & _EVAL_11;
  assign _EVAL_96 = _EVAL_224 | _EVAL_281;
  assign _EVAL_132 = _EVAL_10 & _EVAL_71;
  assign _EVAL_124 = _EVAL_201 | _EVAL_118;
  assign _EVAL_200 = ~_EVAL_144;
  assign _EVAL_155 = _EVAL_244 | _EVAL_2;
  assign _EVAL_60 = _EVAL_68 >> _EVAL_7;
  assign _EVAL_100 = ~_EVAL_275;
  assign _EVAL_275 = _EVAL_146 | _EVAL_2;
  assign _EVAL_46 = _EVAL_272 | _EVAL_2;
  assign _EVAL_116 = _EVAL_3 & _EVAL_82;
  assign _EVAL_263 = _EVAL_39 | _EVAL_196;
  assign _EVAL_19 = _EVAL_11 & _EVAL_16;
  assign _EVAL_277 = _EVAL_1 == 3'h1;
  assign _EVAL_157 = _EVAL_112 | _EVAL_2;
  assign _EVAL_160 = _EVAL_198 | _EVAL_136;
  assign _EVAL_111 = _EVAL_3 ^ 28'hc000000;
  assign _EVAL_92 = ~_EVAL_89;
  assign _EVAL_131 = ~_EVAL_234;
  assign _EVAL_51 = _EVAL_168 | _EVAL_2;
  assign _EVAL_72 = _EVAL_195 | _EVAL_188;
  assign _EVAL_33 = _EVAL_10 & _EVAL_122;
  assign _EVAL_283 = _EVAL_4 >= 3'h2;
  assign _EVAL_62 = $signed(_EVAL_270) & -29'sh400000;
  assign _EVAL_234 = _EVAL_171[0];
  assign _EVAL_90 = ~_EVAL_51;
  assign _EVAL_270 = {1'b0,$signed(_EVAL_111)};
  assign _EVAL_86 = _EVAL_134 | _EVAL_2;
  assign _EVAL_22 = _EVAL_11 & _EVAL_162;
  assign _EVAL_159 = _EVAL_228 & _EVAL_98;
  assign _EVAL_243 = _EVAL_1 == 3'h6;
  assign _EVAL_212 = _EVAL_204 | _EVAL_2;
  assign _EVAL_240 = _EVAL_246 | _EVAL_52;
  assign _EVAL_97 = _EVAL_116 == 28'h0;
  assign _EVAL_68 = _EVAL_36 | _EVAL_268;
  assign _EVAL_36 = _EVAL_21[17:0];
  assign _EVAL_260 = ~_EVAL_104;
  assign _EVAL_130 = 13'h3f << _EVAL_8;
  assign _EVAL_133 = ~_EVAL_75;
  assign _EVAL_163 = _EVAL_160 | _EVAL_2;
  assign _EVAL_258 = _EVAL_1 == 3'h7;
  assign _EVAL_149 = _EVAL_1 == 3'h3;
  assign _EVAL_205 = _EVAL_14 == 3'h2;
  assign _EVAL_241 = _EVAL_84 | _EVAL_2;
  assign _EVAL_55 = _EVAL_1[2];
  assign _EVAL_281 = _EVAL == 5'h10;
  assign _EVAL_140 = _EVAL_181 & _EVAL_193;
  assign _EVAL_27 = ~_EVAL_251;
  assign _EVAL_181 = _EVAL_88 == 2'h0;
  assign _EVAL_224 = _EVAL == 5'h11;
  assign _EVAL_128 = _EVAL_182 - 4'h1;
  assign _EVAL_24 = _EVAL_14 == 3'h0;
  assign _EVAL_123 = _EVAL_11 & _EVAL_277;
  assign _EVAL_171 = _EVAL_268 >> _EVAL;
  assign _EVAL_238 = _EVAL_43 | 2'h1;
  assign _EVAL_186 = _EVAL_14 <= 3'h6;
  assign _EVAL_76 = ~_EVAL_233;
  assign _EVAL_42 = _EVAL_130[5:0];
  assign _EVAL_151 = $signed(_EVAL_105) == 29'sh0;
  assign _EVAL_18 = _EVAL_11 & _EVAL_258;
  assign _EVAL_138 = _EVAL_183 | _EVAL_176;
  assign _EVAL_196 = plusarg_reader_out == 32'h0;
  assign _EVAL_165 = _EVAL_7 == 5'h8;
  assign _EVAL_17 = _EVAL_161 | _EVAL_2;
  assign _EVAL_53 = _EVAL_183 | _EVAL_159;
  assign _EVAL_174 = ~_EVAL_163;
  assign _EVAL_81 = _EVAL_267 | _EVAL_2;
  assign _EVAL_164 = _EVAL_60[0];
  assign _EVAL_69 = _EVAL_11 & _EVAL_243;
  assign _EVAL_242 = ~_EVAL_13;
  assign _EVAL_41 = ~_EVAL_34;
  assign _EVAL_235 = ~_EVAL_232;
  assign _EVAL_38 = ~_EVAL_247;
  assign _EVAL_169 = 3'h6 == _EVAL_4;
  assign _EVAL_29 = ~_EVAL_2;
  assign _EVAL_209 = _EVAL_10 & _EVAL_205;
  assign _EVAL_112 = _EVAL_6 <= 3'h4;
  assign _EVAL_82 = {{22'd0}, _EVAL_92};
  assign _EVAL_143 = _EVAL_14 == _EVAL_28;
  assign _EVAL_115 = _EVAL_118 & _EVAL_215;
  assign _EVAL_110 = ~_EVAL_45;
  assign _EVAL_84 = _EVAL_6 == 3'h0;
  assign _EVAL_48 = _EVAL_268 | _EVAL_36;
  assign _EVAL_192 = _EVAL_10 & _EVAL_24;
  assign _EVAL_273 = ~_EVAL_257;
  assign _EVAL_34 = _EVAL_216 | _EVAL_2;
  assign _EVAL_203 = ~_EVAL_127;
  assign _EVAL_52 = _EVAL_228 & _EVAL_73;
  assign _EVAL_183 = _EVAL_283 | _EVAL_248;
  assign _EVAL_257 = _EVAL_103[17:0];
  assign _EVAL_45 = _EVAL_3[0];
  assign _EVAL_54 = ~_EVAL_122;
  assign _EVAL_266 = _EVAL_118 & _EVAL_125;
  assign _EVAL_226 = ~_EVAL_155;
  always @(posedge _EVAL_12) begin
    if (_EVAL_266) begin
      _EVAL_25 <= _EVAL_8;
    end
    if (_EVAL_266) begin
      _EVAL_28 <= _EVAL_14;
    end
    if (_EVAL_66) begin
      _EVAL_35 <= _EVAL_3;
    end
    if (_EVAL_66) begin
      _EVAL_79 <= _EVAL_4;
    end
    if (_EVAL_66) begin
      _EVAL_145 <= _EVAL_6;
    end
    if (_EVAL_2) begin
      _EVAL_180 <= 4'h0;
    end else if (_EVAL_118) begin
      if (_EVAL_215) begin
        if (_EVAL_178) begin
          _EVAL_180 <= _EVAL_245;
        end else begin
          _EVAL_180 <= 4'h0;
        end
      end else begin
        _EVAL_180 <= _EVAL_113;
      end
    end
    if (_EVAL_2) begin
      _EVAL_182 <= 4'h0;
    end else if (_EVAL_201) begin
      if (_EVAL_202) begin
        if (_EVAL_83) begin
          _EVAL_182 <= _EVAL_147;
        end else begin
          _EVAL_182 <= 4'h0;
        end
      end else begin
        _EVAL_182 <= _EVAL_80;
      end
    end
    if (_EVAL_66) begin
      _EVAL_208 <= _EVAL;
    end
    if (_EVAL_266) begin
      _EVAL_210 <= _EVAL_7;
    end
    if (_EVAL_2) begin
      _EVAL_225 <= 4'h0;
    end else if (_EVAL_118) begin
      if (_EVAL_125) begin
        if (_EVAL_178) begin
          _EVAL_225 <= _EVAL_245;
        end else begin
          _EVAL_225 <= 4'h0;
        end
      end else begin
        _EVAL_225 <= _EVAL_57;
      end
    end
    if (_EVAL_2) begin
      _EVAL_252 <= 32'h0;
    end else if (_EVAL_124) begin
      _EVAL_252 <= 32'h0;
    end else begin
      _EVAL_252 <= _EVAL_221;
    end
    if (_EVAL_66) begin
      _EVAL_253 <= _EVAL_1;
    end
    if (_EVAL_2) begin
      _EVAL_262 <= 4'h0;
    end else if (_EVAL_201) begin
      if (_EVAL_95) begin
        if (_EVAL_83) begin
          _EVAL_262 <= _EVAL_147;
        end else begin
          _EVAL_262 <= 4'h0;
        end
      end else begin
        _EVAL_262 <= _EVAL_166;
      end
    end
    if (_EVAL_2) begin
      _EVAL_268 <= 18'h0;
    end else begin
      _EVAL_268 <= _EVAL_119;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_20) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd589b2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_280) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81f72501)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7740fd5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_254) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48d33483)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9fec35c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_226) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d4ecb9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_20) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_173) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(687f81d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d8a347b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3eda8050)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3aae2342)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_260) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11e088fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(502a6b16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1889c5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3076de1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8589475b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4495450e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62fb6356)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd840969)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(600f1c92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca8b2819)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_203) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d4c15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b81bc45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_203) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31bfe693)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_260) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74ee6189)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(489a3379)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_10 & _EVAL_200) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d26e49c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8e187c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_31) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(917ea7e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74b3e7f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(529a60dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9093eeb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d253493)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d098f65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_31) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78eca0b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91661c15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab244c55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8ddaf39)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0ac1149)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2f0d811)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d94e8648)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58385408)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e9ba579)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56c16c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee1d481a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c87fa1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d0748fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_209 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8d8ab0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0bd9344)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5fe06705)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(880ec6ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_174) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c7c2c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa39f125)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(598ec3cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9518a708)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(132659e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f79e4174)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_40 & _EVAL_173) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_280) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9ed87fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8d8ab0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c06285f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_44 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f03f35f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ff3fcad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_279) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3df604b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9db00002)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22e7fa2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_132 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_237) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b0e199f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cae6bc3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_174) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_226) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9df2b631)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7db72dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_38) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81cc08a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54e5f540)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6852f032)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_207 & _EVAL_38) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f53aad1e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_237) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_108 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_18 & _EVAL_279) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_78 & _EVAL_179) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4ea521c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_10 & _EVAL_200) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb95c4b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_278) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d17facc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f9d5a98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_25 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_28 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_35 = _RAND_2[27:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_79 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_145 = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_180 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_182 = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_208 = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_210 = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_225 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_252 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_253 = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_262 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_268 = _RAND_13[17:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
