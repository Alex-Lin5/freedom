//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_175_assert(
  input  [2:0]  _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input  [9:0]  _EVAL_2,
  input  [1:0]  _EVAL_3,
  input  [11:0] _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [2:0]  _EVAL_7,
  input  [1:0]  _EVAL_8,
  input  [9:0]  _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  input  [3:0]  _EVAL_14
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [575:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_15;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  reg [2:0] _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire [32:0] _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire [3:0] _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire [1:0] _EVAL_46;
  reg [1:0] _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire [31:0] _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  reg  _EVAL_56;
  wire  _EVAL_57;
  reg [2:0] _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire [1:0] _EVAL_69;
  wire  _EVAL_70;
  wire [575:0] _EVAL_71;
  wire [575:0] _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire [11:0] _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire [1023:0] _EVAL_87;
  reg [9:0] _EVAL_88;
  reg  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire [575:0] _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire [1:0] _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  reg [575:0] _EVAL_113;
  wire  _EVAL_114;
  reg [2:0] _EVAL_115;
  wire [1023:0] _EVAL_117;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire [12:0] _EVAL_121;
  wire [1:0] _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire [1:0] _EVAL_127;
  wire  _EVAL_128;
  wire [575:0] _EVAL_129;
  wire [575:0] _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire  _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  reg [11:0] _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire [1:0] _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire [12:0] _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  reg  _EVAL_158;
  wire  _EVAL_159;
  wire [1023:0] _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  reg [9:0] _EVAL_163;
  wire  _EVAL_164;
  wire [575:0] _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire [1:0] _EVAL_168;
  wire  _EVAL_169;
  wire [11:0] _EVAL_170;
  wire [1023:0] _EVAL_171;
  wire [3:0] _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  reg [31:0] _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire [12:0] _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  reg [1:0] _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire [575:0] _EVAL_202;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire [3:0] _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire [1:0] _EVAL_222;
  wire [4:0] _EVAL_223;
  wire  _EVAL_224;
  wire [3:0] _EVAL_225;
  wire  _EVAL_226;
  wire [575:0] _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  reg  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_179 = _EVAL_6 & _EVAL_20;
  assign _EVAL_76 = ~_EVAL_10;
  assign _EVAL_148 = _EVAL_219 | _EVAL_10;
  assign _EVAL_141 = ~_EVAL_156;
  assign _EVAL_175 = _EVAL_176 < plusarg_reader_out;
  assign _EVAL_186 = _EVAL_14 == _EVAL_225;
  assign _EVAL_33 = _EVAL_176 + 32'h1;
  assign _EVAL_210 = _EVAL_143 | _EVAL_10;
  assign _EVAL_37 = _EVAL_74 | _EVAL_10;
  assign _EVAL_24 = _EVAL_4[1];
  assign _EVAL_93 = _EVAL_147 | _EVAL_10;
  assign _EVAL_146 = _EVAL_46[0];
  assign _EVAL_237 = _EVAL_177 & _EVAL_98;
  assign _EVAL_206 = _EVAL_71[0];
  assign _EVAL_43 = _EVAL_13 & _EVAL_105;
  assign _EVAL_64 = _EVAL_112 | _EVAL_10;
  assign _EVAL_102 = _EVAL_172 == 4'h0;
  assign _EVAL_61 = _EVAL_13 & _EVAL_70;
  assign _EVAL_72 = _EVAL_113 | _EVAL_130;
  assign _EVAL_67 = ~_EVAL_215;
  assign _EVAL_215 = _EVAL_39 | _EVAL_10;
  assign _EVAL_134 = _EVAL_8 >= 2'h2;
  assign _EVAL_169 = _EVAL == 3'h0;
  assign _EVAL_156 = _EVAL_25 | _EVAL_10;
  assign _EVAL_92 = ~_EVAL_11;
  assign _EVAL_155 = {1'b0,$signed(_EVAL_4)};
  assign _EVAL_123 = ~_EVAL_110;
  assign _EVAL_159 = _EVAL_101 | _EVAL_10;
  assign _EVAL_234 = _EVAL_5 & _EVAL_13;
  assign _EVAL_84 = _EVAL_7 == 3'h2;
  assign _EVAL_197 = _EVAL_7 == 3'h4;
  assign _EVAL_184 = ~_EVAL_40;
  assign _EVAL_97 = _EVAL_7 == 3'h6;
  assign _EVAL_231 = ~_EVAL_93;
  assign _EVAL_46 = _EVAL_158 - 1'h1;
  assign _EVAL_22 = _EVAL_7 == 3'h5;
  assign _EVAL_45 = _EVAL_226 | _EVAL_10;
  assign _EVAL_105 = _EVAL_12 == 3'h2;
  assign _EVAL_145 = _EVAL_102 | _EVAL_10;
  assign _EVAL_152 = ~_EVAL_69;
  assign _EVAL_57 = _EVAL_229 | _EVAL_21;
  assign _EVAL_25 = _EVAL_9 <= 10'h23f;
  assign _EVAL_187 = plusarg_reader_out == 32'h0;
  assign _EVAL_213 = ~_EVAL_218;
  assign _EVAL_201 = _EVAL_122[0];
  assign _EVAL_60 = _EVAL_107 | _EVAL_10;
  assign _EVAL_153 = ~_EVAL_150;
  assign _EVAL_181 = _EVAL_234 & _EVAL_29;
  assign _EVAL_164 = ~_EVAL_190;
  assign _EVAL_48 = _EVAL_86 | _EVAL_114;
  assign _EVAL_228 = _EVAL_12 == 3'h0;
  assign _EVAL_191 = _EVAL_3 >= 2'h2;
  assign _EVAL_101 = _EVAL_2 == _EVAL_163;
  assign _EVAL_126 = _EVAL_127[1];
  assign _EVAL_229 = _EVAL_134 | _EVAL_63;
  assign _EVAL_162 = _EVAL <= 3'h3;
  assign _EVAL_121 = $signed(_EVAL_155) & 13'sh1000;
  assign _EVAL_183 = _EVAL_121;
  assign _EVAL_71 = _EVAL_113 >> _EVAL_9;
  assign _EVAL_107 = _EVAL_12 <= 3'h6;
  assign _EVAL_199 = _EVAL_236 | _EVAL_10;
  assign _EVAL_154 = ~_EVAL_37;
  assign _EVAL_143 = _EVAL != 3'h0;
  assign _EVAL_26 = ~_EVAL_31;
  assign _EVAL_223 = 5'h3 << _EVAL_8;
  assign _EVAL_81 = _EVAL_7 == 3'h3;
  assign _EVAL_217 = ~_EVAL_132;
  assign _EVAL_18 = ~_EVAL_180;
  assign _EVAL_230 = _EVAL_6 & _EVAL_22;
  assign _EVAL_220 = _EVAL_4[0];
  assign _EVAL_174 = _EVAL_92 | _EVAL_10;
  assign _EVAL_188 = ~_EVAL_60;
  assign _EVAL_226 = _EVAL <= 3'h4;
  assign _EVAL_127 = _EVAL_222 | 2'h1;
  assign _EVAL_133 = _EVAL_34 & _EVAL_216;
  assign _EVAL_74 = _EVAL_212 == 4'h0;
  assign _EVAL_190 = _EVAL_32 | _EVAL_10;
  assign _EVAL_35 = _EVAL_7 == 3'h0;
  assign _EVAL_136 = _EVAL_6 & _EVAL_197;
  assign _EVAL_211 = _EVAL_13 & _EVAL_42;
  assign _EVAL_114 = _EVAL_177 & _EVAL_77;
  assign _EVAL_173 = _EVAL <= 3'h1;
  assign _EVAL_204 = _EVAL_85 | _EVAL_10;
  assign _EVAL_178 = _EVAL_7 == 3'h1;
  assign _EVAL_160 = _EVAL_133 ? _EVAL_87 : 1024'h0;
  assign _EVAL_62 = ~_EVAL_128;
  assign _EVAL_40 = _EVAL_134 | _EVAL_10;
  assign _EVAL_63 = _EVAL_126 & _EVAL_24;
  assign _EVAL_144 = ~_EVAL_145;
  assign _EVAL_218 = _EVAL_169 | _EVAL_10;
  assign _EVAL_95 = ~_EVAL_210;
  assign _EVAL_20 = _EVAL_7 == 3'h7;
  assign _EVAL_17 = _EVAL_13 & _EVAL_119;
  assign _EVAL_75 = _EVAL_234 & _EVAL_44;
  assign _EVAL_39 = _EVAL <= 3'h2;
  assign _EVAL_165 = _EVAL_202 >> _EVAL_2;
  assign _EVAL_205 = _EVAL_12 == 3'h6;
  assign _EVAL_198 = _EVAL_125 | _EVAL_10;
  assign _EVAL_98 = _EVAL_24 & _EVAL_220;
  assign _EVAL_73 = _EVAL_86 | _EVAL_99;
  assign _EVAL_120 = _EVAL_6 & _EVAL_97;
  assign _EVAL_104 = _EVAL_34 | _EVAL_234;
  assign _EVAL_185 = _EVAL_6 & _EVAL_81;
  assign _EVAL_16 = _EVAL_139 | _EVAL_10;
  assign _EVAL_212 = ~_EVAL_14;
  assign _EVAL_70 = _EVAL_12 == 3'h1;
  assign _EVAL_19 = _EVAL_6 & _EVAL_178;
  assign _EVAL_222 = 2'h1 << _EVAL_28;
  assign _EVAL_85 = _EVAL_25 & _EVAL_36;
  assign _EVAL_51 = ~_EVAL_45;
  assign _EVAL_111 = _EVAL_75 & _EVAL_200;
  assign _EVAL_236 = _EVAL == _EVAL_23;
  assign _EVAL_209 = _EVAL_186 | _EVAL_10;
  assign _EVAL_54 = _EVAL_232 | _EVAL_10;
  assign _EVAL_208 = _EVAL_6 & _EVAL_84;
  assign _EVAL_172 = _EVAL_14 & _EVAL_38;
  assign _EVAL_32 = _EVAL_2 <= 10'h23f;
  assign _EVAL_128 = _EVAL_173 | _EVAL_10;
  assign _EVAL_167 = ~_EVAL_78;
  assign _EVAL_170 = _EVAL_4 & _EVAL_83;
  assign _EVAL_135 = ~_EVAL_195;
  assign _EVAL_110 = _EVAL_55 | _EVAL_10;
  assign _EVAL_232 = _EVAL_41 | _EVAL_175;
  assign _EVAL_86 = _EVAL_134 | _EVAL_137;
  assign _EVAL_119 = _EVAL_12 == 3'h4;
  assign _EVAL_161 = _EVAL_8 <= 2'h2;
  assign _EVAL_192 = _EVAL_13 & _EVAL_228;
  assign _EVAL_82 = ~_EVAL_206;
  assign _EVAL_59 = _EVAL_4 == _EVAL_149;
  assign _EVAL_195 = _EVAL_82 | _EVAL_10;
  assign _EVAL_66 = ~_EVAL_204;
  assign _EVAL_91 = _EVAL_79 | _EVAL_10;
  assign _EVAL_69 = _EVAL_223[1:0];
  assign _EVAL_166 = _EVAL_34 & _EVAL_78;
  assign _EVAL_138 = ~_EVAL_64;
  assign _EVAL_28 = _EVAL_8[0];
  assign _EVAL_87 = 1024'h1 << _EVAL_9;
  assign _EVAL_139 = _EVAL_12 == _EVAL_58;
  assign _EVAL_53 = _EVAL_33[31:0];
  assign _EVAL_137 = _EVAL_126 & _EVAL_193;
  assign _EVAL_49 = _EVAL_6 & _EVAL_35;
  assign _EVAL_122 = _EVAL_233 - 1'h1;
  assign _EVAL_34 = _EVAL_0 & _EVAL_6;
  assign _EVAL_130 = _EVAL_160[575:0];
  assign _EVAL_132 = _EVAL_162 | _EVAL_10;
  assign _EVAL_42 = ~_EVAL_29;
  assign _EVAL_216 = ~_EVAL_233;
  assign _EVAL_41 = _EVAL_52 | _EVAL_187;
  assign _EVAL_106 = _EVAL_13 & _EVAL_205;
  assign _EVAL_219 = _EVAL_170 == 12'h0;
  assign _EVAL_200 = ~_EVAL_205;
  assign _EVAL_202 = _EVAL_130 | _EVAL_113;
  assign _EVAL_168 = _EVAL_89 - 1'h1;
  assign _EVAL_100 = ~_EVAL_159;
  assign _EVAL_77 = _EVAL_193 & _EVAL_15;
  assign _EVAL_129 = _EVAL_171[575:0];
  assign _EVAL_193 = ~_EVAL_24;
  assign _EVAL_27 = ~_EVAL_54;
  assign _EVAL_44 = ~_EVAL_56;
  assign _EVAL_224 = _EVAL_103[0];
  assign _EVAL_171 = _EVAL_111 ? _EVAL_117 : 1024'h0;
  assign _EVAL_227 = ~_EVAL_129;
  assign _EVAL_214 = _EVAL_13 & _EVAL_221;
  assign _EVAL_235 = ~_EVAL_174;
  assign _EVAL_52 = ~_EVAL_151;
  assign _EVAL_207 = ~_EVAL_148;
  assign _EVAL_29 = ~_EVAL_89;
  assign _EVAL_140 = _EVAL_6 & _EVAL_167;
  assign _EVAL_96 = _EVAL_72 & _EVAL_227;
  assign _EVAL_90 = ~_EVAL_198;
  assign _EVAL_142 = _EVAL_193 & _EVAL_220;
  assign _EVAL_31 = _EVAL_191 | _EVAL_10;
  assign _EVAL_151 = |_EVAL_113;
  assign _EVAL_150 = _EVAL_59 | _EVAL_10;
  assign _EVAL_177 = _EVAL_127[0];
  assign _EVAL_157 = _EVAL_24 & _EVAL_15;
  assign _EVAL_125 = _EVAL_165[0];
  assign _EVAL_83 = {{10'd0}, _EVAL_152};
  assign _EVAL_36 = _EVAL_161 & _EVAL_108;
  assign _EVAL_68 = ~_EVAL_91;
  assign _EVAL_103 = _EVAL_56 - 1'h1;
  assign _EVAL_108 = $signed(_EVAL_183) == 13'sh0;
  assign _EVAL_194 = _EVAL_229 | _EVAL_237;
  assign _EVAL_131 = _EVAL_168[0];
  assign _EVAL_15 = ~_EVAL_220;
  assign _EVAL_80 = ~_EVAL_199;
  assign _EVAL_225 = {_EVAL_194,_EVAL_57,_EVAL_73,_EVAL_48};
  assign _EVAL_79 = _EVAL_9 == _EVAL_88;
  assign _EVAL_147 = _EVAL_3 == _EVAL_189;
  assign _EVAL_221 = _EVAL_12 == 3'h5;
  assign _EVAL_94 = ~_EVAL_16;
  assign _EVAL_65 = ~_EVAL_209;
  assign _EVAL_180 = _EVAL_36 | _EVAL_10;
  assign _EVAL_55 = _EVAL_7 == _EVAL_115;
  assign _EVAL_99 = _EVAL_177 & _EVAL_142;
  assign _EVAL_117 = 1024'h1 << _EVAL_2;
  assign _EVAL_112 = _EVAL_8 == _EVAL_47;
  assign _EVAL_21 = _EVAL_177 & _EVAL_157;
  assign _EVAL_78 = ~_EVAL_158;
  assign _EVAL_38 = ~_EVAL_225;
  always @(posedge _EVAL_1) begin
    if (_EVAL_166) begin
      _EVAL_23 <= _EVAL;
    end
    if (_EVAL_166) begin
      _EVAL_47 <= _EVAL_8;
    end
    if (_EVAL_10) begin
      _EVAL_56 <= 1'h0;
    end else if (_EVAL_234) begin
      if (_EVAL_44) begin
        _EVAL_56 <= 1'h0;
      end else begin
        _EVAL_56 <= _EVAL_224;
      end
    end
    if (_EVAL_181) begin
      _EVAL_58 <= _EVAL_12;
    end
    if (_EVAL_166) begin
      _EVAL_88 <= _EVAL_9;
    end
    if (_EVAL_10) begin
      _EVAL_89 <= 1'h0;
    end else if (_EVAL_234) begin
      if (_EVAL_29) begin
        _EVAL_89 <= 1'h0;
      end else begin
        _EVAL_89 <= _EVAL_131;
      end
    end
    if (_EVAL_10) begin
      _EVAL_113 <= 576'h0;
    end else begin
      _EVAL_113 <= _EVAL_96;
    end
    if (_EVAL_166) begin
      _EVAL_115 <= _EVAL_7;
    end
    if (_EVAL_166) begin
      _EVAL_149 <= _EVAL_4;
    end
    if (_EVAL_10) begin
      _EVAL_158 <= 1'h0;
    end else if (_EVAL_34) begin
      if (_EVAL_78) begin
        _EVAL_158 <= 1'h0;
      end else begin
        _EVAL_158 <= _EVAL_146;
      end
    end
    if (_EVAL_181) begin
      _EVAL_163 <= _EVAL_2;
    end
    if (_EVAL_10) begin
      _EVAL_176 <= 32'h0;
    end else if (_EVAL_104) begin
      _EVAL_176 <= 32'h0;
    end else begin
      _EVAL_176 <= _EVAL_53;
    end
    if (_EVAL_181) begin
      _EVAL_189 <= _EVAL_3;
    end
    if (_EVAL_10) begin
      _EVAL_233 <= 1'h0;
    end else if (_EVAL_34) begin
      if (_EVAL_216) begin
        _EVAL_233 <= 1'h0;
      end else begin
        _EVAL_233 <= _EVAL_201;
      end
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70e35f32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab22e21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a15206c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_144) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1564e979)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_80) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b14d46cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa907d5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7ee2d20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9afe0899)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_100) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52b8224e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8574b466)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_67) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff8f7ea9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6061a5e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff407ebd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_13 & _EVAL_188) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1660c443)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_90) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7cb045)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(793f1f1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1113997)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4de799a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_66) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e071cbaf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98d44a70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdf3a643)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_153) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(279ac5cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5fe7fd8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef9183a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_95) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed3ac213)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_13 & _EVAL_188) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(115d2930)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(194a04f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_100) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3332466)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2337dd7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_90) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffb809b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a97a87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30ac6e9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_213) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6faebcf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ece62ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2693eb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8299c87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56a315e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d767c5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d7c96ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_26) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_68) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be1e8ef3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_18) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae6878e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_153) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22e4dc0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa3e1bd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(56c0c883)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(746336ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_144) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ee5a155)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c0933ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3effe0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_65) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(483ffb65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_214 & _EVAL_26) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9cc4670)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_106 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e51e323f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_17 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(991eb578)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a450f9c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_135) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_95) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30bf14be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ffacf11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_67) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ed60927)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_80) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_133 & _EVAL_135) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb916d10)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_43 & _EVAL_164) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(53d65c59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ecedf2c1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_68) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc1cacb6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf6ed1aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_207) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a5dfeee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a130f1bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c436f45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_49 & _EVAL_66) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1e2db2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_120 & _EVAL_154) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e974ad59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62839c00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eab67122)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_136 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3de5cf70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_141) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8cef668)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4262a5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_65) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_140 & _EVAL_138) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6999d74a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_207) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_179 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff407ebd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_185 & _EVAL_141) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c5983d2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_213) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd7f2ff6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_19 & _EVAL_18) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_61 & _EVAL_164) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_23 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_47 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_56 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_58 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_88 = _RAND_4[9:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_89 = _RAND_5[0:0];
  _RAND_6 = {18{`RANDOM}};
  _EVAL_113 = _RAND_6[575:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_115 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_149 = _RAND_8[11:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_158 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_163 = _RAND_10[9:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_176 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_189 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_233 = _RAND_13[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
