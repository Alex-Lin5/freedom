//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module CoreIPSubsystemAllPortRAMTestHarness(
  input   clock,
  input   reset,
  output  io_success
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
`endif // RANDOMIZE_REG_INIT
  wire  system_clock;
  wire  system_reset;
  wire  system_external_source_for_core_0_clock;
  wire  system_external_source_for_core_0_reset;
  wire  system_halt_from_tile_0;
  wire  system_wfi_from_tile_0;
  wire  system_cease_from_tile_0;
  wire  system_debug_from_tile_0;
  wire  system_psd_test_clock_enable;
  wire  system_resetctrl_hartIsInReset_0;
  wire  system_debug_clock;
  wire  system_debug_reset;
  wire  system_debug_systemjtag_jtag_TCK;
  wire  system_debug_systemjtag_jtag_TMS;
  wire  system_debug_systemjtag_jtag_TDI;
  wire  system_debug_systemjtag_jtag_TDO_data;
  wire  system_debug_systemjtag_jtag_TDO_driven;
  wire  system_debug_systemjtag_reset;
  wire [10:0] system_debug_systemjtag_mfr_id;
  wire [15:0] system_debug_systemjtag_part_number;
  wire [3:0] system_debug_systemjtag_version;
  wire  system_debug_ndreset;
  wire  system_debug_dmactive;
  wire  system_debug_dmactiveAck;
  wire [31:0] system_reset_vector_0;
  wire  system_nmi_0_rnmi;
  wire [31:0] system_nmi_0_rnmi_interrupt_vector;
  wire [31:0] system_nmi_0_rnmi_exception_vector;
  wire  system_rtc_toggle;
  wire [126:0] system_global_interrupts;
  wire [15:0] system_local_interrupts_0;
  wire  system_sys_port_ahb_0_hmastlock;
  wire  system_sys_port_ahb_0_hready;
  wire [1:0] system_sys_port_ahb_0_htrans;
  wire [2:0] system_sys_port_ahb_0_hsize;
  wire [2:0] system_sys_port_ahb_0_hburst;
  wire  system_sys_port_ahb_0_hwrite;
  wire [3:0] system_sys_port_ahb_0_hprot;
  wire [30:0] system_sys_port_ahb_0_haddr;
  wire [31:0] system_sys_port_ahb_0_hwdata;
  wire  system_sys_port_ahb_0_hresp;
  wire [31:0] system_sys_port_ahb_0_hrdata;
  wire  system_periph_port_ahb_0_hmastlock;
  wire  system_periph_port_ahb_0_hready;
  wire [1:0] system_periph_port_ahb_0_htrans;
  wire [2:0] system_periph_port_ahb_0_hsize;
  wire [2:0] system_periph_port_ahb_0_hburst;
  wire  system_periph_port_ahb_0_hwrite;
  wire [3:0] system_periph_port_ahb_0_hprot;
  wire [29:0] system_periph_port_ahb_0_haddr;
  wire [31:0] system_periph_port_ahb_0_hwdata;
  wire  system_periph_port_ahb_0_hresp;
  wire [31:0] system_periph_port_ahb_0_hrdata;
  wire  system_front_port_ahb_0_hmastlock;
  wire  system_front_port_ahb_0_hsel;
  wire  system_front_port_ahb_0_hready;
  wire  system_front_port_ahb_0_hreadyout;
  wire [1:0] system_front_port_ahb_0_htrans;
  wire [2:0] system_front_port_ahb_0_hsize;
  wire [2:0] system_front_port_ahb_0_hburst;
  wire  system_front_port_ahb_0_hwrite;
  wire [3:0] system_front_port_ahb_0_hprot;
  wire [31:0] system_front_port_ahb_0_haddr;
  wire [31:0] system_front_port_ahb_0_hwdata;
  wire  system_front_port_ahb_0_hresp;
  wire [31:0] system_front_port_ahb_0_hrdata;
  wire  func_clock_clock;
  wire  func_clock_io_clock_out;
  wire  system_clock_divider_clock;
  wire  system_clock_divider_io_clock_out;
  wire  core_clocks_skew_clkin;
  wire  core_clocks_skew_clkout;
  wire  dpiClockGate_clock_in;
  wire  dpiClockGate_clock_out;
  wire [31:0] plusarg_reader_out;
  wire  c_core_reset_driver_clock;
  wire  c_core_reset_driver_out;
  wire  debug_compatibility_clock;
  wire  debug_compatibility_debug_outer_reset;
  wire  debug_compatibility_core_resets_in_0;
  wire  debug_compatibility_debug_clock;
  wire  debug_compatibility_debug_reset;
  wire  debug_compatibility_debug_dmactive;
  wire  debug_compatibility_debug_dmactiveAck;
  wire  debug_compatibility_debug_resetctrl_hartIsInReset_0;
  wire  debug_compatibility_core_resets_out_0;
  wire [31:0] plusarg_reader_1_out;
  wire  delayed_reset_count_and_driver_clock;
  wire  delayed_reset_count_and_driver_reset;
  wire  delayed_reset_count_and_driver_io_default_value;
  wire [15:0] delayed_reset_count_and_driver_io_count;
  wire  delayed_reset_count_and_driver_io_driven_value;
  wire  coreTraces_DataTap_10__0_clock;
  wire  coreTraces_DataTap_10__0_reset;
  wire  coreTraces_DataTap_10__0_excpt;
  wire [2:0] coreTraces_DataTap_10__0_priv_mode;
  wire [31:0] coreTraces_DataTap_10__0_hartid;
  wire [31:0] coreTraces_DataTap_10__0_timer;
  wire  coreTraces_DataTap_10__0_valid;
  wire [31:0] coreTraces_DataTap_10__0_pc;
  wire [4:0] coreTraces_DataTap_10__0_wrdst;
  wire [31:0] coreTraces_DataTap_10__0_wrdata;
  wire  coreTraces_DataTap_10__0_wrenx;
  wire  coreTraces_DataTap_10__0_wrenf;
  wire [4:0] coreTraces_DataTap_10__0_rd0src;
  wire [31:0] coreTraces_DataTap_10__0_rd0val;
  wire [4:0] coreTraces_DataTap_10__0_rd1src;
  wire [31:0] coreTraces_DataTap_10__0_rd1val;
  wire [31:0] coreTraces_DataTap_10__0_inst;
  wire  csrTraces_DataTap_1__9;
  wire  csrTraces_DataTap_1__8;
  wire  csrTraces_DataTap_1__7;
  wire  csrTraces_DataTap_1__6;
  wire [31:0] csrTraces_DataTap_1__5;
  wire [31:0] csrTraces_DataTap_1__4;
  wire [31:0] csrTraces_DataTap_1__3;
  wire [31:0] csrTraces_DataTap_1__2;
  wire [31:0] csrTraces_DataTap_1__1;
  wire  csrTraces_DataTap_1__0;
  wire  testRAM_clock;
  wire  testRAM_reset;
  wire  testRAM_io_ahb_0_hmastlock;
  wire  testRAM_io_ahb_0_hready;
  wire [1:0] testRAM_io_ahb_0_htrans;
  wire [2:0] testRAM_io_ahb_0_hsize;
  wire [2:0] testRAM_io_ahb_0_hburst;
  wire  testRAM_io_ahb_0_hwrite;
  wire [3:0] testRAM_io_ahb_0_hprot;
  wire [29:0] testRAM_io_ahb_0_haddr;
  wire [31:0] testRAM_io_ahb_0_hwdata;
  wire  testRAM_io_ahb_0_hresp;
  wire [31:0] testRAM_io_ahb_0_hrdata;
  wire  system_periph_port_ahb_0_hrdata_xs_valid;
  wire [31:0] system_periph_port_ahb_0_hrdata_xs_inp;
  wire [31:0] system_periph_port_ahb_0_hrdata_xs_outp;
  wire  system_periph_port_ahb_0_hresp_xs_valid;
  wire  system_periph_port_ahb_0_hresp_xs_inp;
  wire  system_periph_port_ahb_0_hresp_xs_outp;
  wire  testRAM_1_clock;
  wire  testRAM_1_reset;
  wire  testRAM_1_io_ahb_0_hmastlock;
  wire  testRAM_1_io_ahb_0_hready;
  wire [1:0] testRAM_1_io_ahb_0_htrans;
  wire [2:0] testRAM_1_io_ahb_0_hsize;
  wire [2:0] testRAM_1_io_ahb_0_hburst;
  wire  testRAM_1_io_ahb_0_hwrite;
  wire [3:0] testRAM_1_io_ahb_0_hprot;
  wire [30:0] testRAM_1_io_ahb_0_haddr;
  wire [31:0] testRAM_1_io_ahb_0_hwdata;
  wire  testRAM_1_io_ahb_0_hresp;
  wire [31:0] testRAM_1_io_ahb_0_hrdata;
  wire  system_sys_port_ahb_0_hrdata_xs_valid;
  wire [31:0] system_sys_port_ahb_0_hrdata_xs_inp;
  wire [31:0] system_sys_port_ahb_0_hrdata_xs_outp;
  wire  system_sys_port_ahb_0_hresp_xs_valid;
  wire  system_sys_port_ahb_0_hresp_xs_inp;
  wire  system_sys_port_ahb_0_hresp_xs_outp;
  wire  wfichecker_reset;
  wire  wfichecker_clock;
  wire  wfichecker_wfi;
  wire [31:0] wfichecker_csr_hartid;
  wire  wfichecker_excpt;
  wire  wfichecker_bus_err_int;
  wire  wfichecker_debug_int;
  wire  wfichecker_clint_int;
  wire  wfichecker_allow_wfi;
  wire  wfichecker_debug;
  wire  wfichecker_singleStep;
  wire [31:0] wfichecker_reg_mie;
  wire [31:0] wfichecker_reg_mip;
  wire [31:0] wfichecker_inst_hartid_0;
  wire  wfichecker_inst_vld_0;
  wire [31:0] wfichecker_pc_0;
  wire [31:0] wfichecker_inst_0;
  wire  core_monitor_m_0_clock;
  wire  core_monitor_m_0_reset;
  wire  core_monitor_m_0_excpt;
  wire [2:0] core_monitor_m_0_priv_mode;
  wire [31:0] core_monitor_m_0_hartid;
  wire [31:0] core_monitor_m_0_timer;
  wire  core_monitor_m_0_valid;
  wire [31:0] core_monitor_m_0_pc;
  wire [4:0] core_monitor_m_0_wrdst;
  wire [31:0] core_monitor_m_0_wrdata;
  wire  core_monitor_m_0_wrenx;
  wire  core_monitor_m_0_wrenf;
  wire [4:0] core_monitor_m_0_rd0src;
  wire [31:0] core_monitor_m_0_rd0val;
  wire [4:0] core_monitor_m_0_rd1src;
  wire [31:0] core_monitor_m_0_rd1val;
  wire [31:0] core_monitor_m_0_inst;
  wire  dpitbh_clock;
  wire  dpitbh_reset;
  wire [31:0] plusarg_reader_2_out;
  wire  dpi_driver_clock;
  wire  dpi_driver_reset;
  wire [126:0] dpi_driver_interrupts;
  wire [31:0] plusarg_reader_3_out;
  wire  dpi_drivers_0_clock;
  wire  dpi_drivers_0_reset;
  wire [31:0] dpi_drivers_0_interrupts;
  reg [4:0] count;
  reg  toggle;
  wire [4:0] _count_T_1 = count + 5'h1;
  wire  ram_reset = system_reset | reset;
  wire  ndm_reset = reset | system_debug_ndreset;
  reg  system_periph_port_ahb_0_hrdata_xs_io_valid_r;
  reg  system_periph_port_ahb_0_hrdata_xs_io_valid_r_1;
  reg  system_periph_port_ahb_0_hresp_xs_io_valid_r;
  reg  system_sys_port_ahb_0_hrdata_xs_io_valid_r;
  reg  system_sys_port_ahb_0_hrdata_xs_io_valid_r_1;
  reg  system_sys_port_ahb_0_hresp_xs_io_valid_r;
  reg [6:0] tick_value;
  wire  tick = tick_value == 7'h63;
  wire [6:0] _tick_value_T_1 = tick_value + 7'h1;
  wire [31:0] drive_interrupt_type = plusarg_reader_2_out;
  reg [6:0] system_global_interrupts_value;
  wire  system_global_interrupts_wrap_wrap = system_global_interrupts_value == 7'h7e;
  wire [6:0] _system_global_interrupts_wrap_value_T_1 = system_global_interrupts_value + 7'h1;
  wire [127:0] _system_global_interrupts_T_2 = 128'h1 << system_global_interrupts_value;
  reg [15:0] tickers_x3_lfsrReg;
  wire  tickers_x3_lfsrReg_hi = tickers_x3_lfsrReg[0] ^ tickers_x3_lfsrReg[2] ^ tickers_x3_lfsrReg[3] ^
    tickers_x3_lfsrReg[5];
  wire [14:0] tickers_x3_lfsrReg_lo = tickers_x3_lfsrReg[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_6 = {tickers_x3_lfsrReg_hi,tickers_x3_lfsrReg_lo};
  reg [15:0] tickers_x3_lfsrReg_1;
  wire  tickers_x3_lfsrReg_hi_1 = tickers_x3_lfsrReg_1[0] ^ tickers_x3_lfsrReg_1[2] ^ tickers_x3_lfsrReg_1[3] ^
    tickers_x3_lfsrReg_1[5];
  wire [14:0] tickers_x3_lfsrReg_lo_1 = tickers_x3_lfsrReg_1[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_13 = {tickers_x3_lfsrReg_hi_1,tickers_x3_lfsrReg_lo_1};
  reg [15:0] tickers_x3_lfsrReg_2;
  wire  tickers_x3_lfsrReg_hi_2 = tickers_x3_lfsrReg_2[0] ^ tickers_x3_lfsrReg_2[2] ^ tickers_x3_lfsrReg_2[3] ^
    tickers_x3_lfsrReg_2[5];
  wire [14:0] tickers_x3_lfsrReg_lo_2 = tickers_x3_lfsrReg_2[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_20 = {tickers_x3_lfsrReg_hi_2,tickers_x3_lfsrReg_lo_2};
  reg [15:0] tickers_x3_lfsrReg_3;
  wire  tickers_x3_lfsrReg_hi_3 = tickers_x3_lfsrReg_3[0] ^ tickers_x3_lfsrReg_3[2] ^ tickers_x3_lfsrReg_3[3] ^
    tickers_x3_lfsrReg_3[5];
  wire [14:0] tickers_x3_lfsrReg_lo_3 = tickers_x3_lfsrReg_3[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_27 = {tickers_x3_lfsrReg_hi_3,tickers_x3_lfsrReg_lo_3};
  reg [15:0] tickers_x3_lfsrReg_4;
  wire  tickers_x3_lfsrReg_hi_4 = tickers_x3_lfsrReg_4[0] ^ tickers_x3_lfsrReg_4[2] ^ tickers_x3_lfsrReg_4[3] ^
    tickers_x3_lfsrReg_4[5];
  wire [14:0] tickers_x3_lfsrReg_lo_4 = tickers_x3_lfsrReg_4[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_34 = {tickers_x3_lfsrReg_hi_4,tickers_x3_lfsrReg_lo_4};
  reg [15:0] tickers_x3_lfsrReg_5;
  wire  tickers_x3_lfsrReg_hi_5 = tickers_x3_lfsrReg_5[0] ^ tickers_x3_lfsrReg_5[2] ^ tickers_x3_lfsrReg_5[3] ^
    tickers_x3_lfsrReg_5[5];
  wire [14:0] tickers_x3_lfsrReg_lo_5 = tickers_x3_lfsrReg_5[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_41 = {tickers_x3_lfsrReg_hi_5,tickers_x3_lfsrReg_lo_5};
  reg [15:0] tickers_x3_lfsrReg_6;
  wire  tickers_x3_lfsrReg_hi_6 = tickers_x3_lfsrReg_6[0] ^ tickers_x3_lfsrReg_6[2] ^ tickers_x3_lfsrReg_6[3] ^
    tickers_x3_lfsrReg_6[5];
  wire [14:0] tickers_x3_lfsrReg_lo_6 = tickers_x3_lfsrReg_6[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_48 = {tickers_x3_lfsrReg_hi_6,tickers_x3_lfsrReg_lo_6};
  reg [15:0] tickers_x3_lfsrReg_7;
  wire  tickers_x3_lfsrReg_hi_7 = tickers_x3_lfsrReg_7[0] ^ tickers_x3_lfsrReg_7[2] ^ tickers_x3_lfsrReg_7[3] ^
    tickers_x3_lfsrReg_7[5];
  wire [14:0] tickers_x3_lfsrReg_lo_7 = tickers_x3_lfsrReg_7[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_55 = {tickers_x3_lfsrReg_hi_7,tickers_x3_lfsrReg_lo_7};
  reg [15:0] tickers_x3_lfsrReg_8;
  wire  tickers_x3_lfsrReg_hi_8 = tickers_x3_lfsrReg_8[0] ^ tickers_x3_lfsrReg_8[2] ^ tickers_x3_lfsrReg_8[3] ^
    tickers_x3_lfsrReg_8[5];
  wire [14:0] tickers_x3_lfsrReg_lo_8 = tickers_x3_lfsrReg_8[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_62 = {tickers_x3_lfsrReg_hi_8,tickers_x3_lfsrReg_lo_8};
  reg [15:0] tickers_x3_lfsrReg_9;
  wire  tickers_x3_lfsrReg_hi_9 = tickers_x3_lfsrReg_9[0] ^ tickers_x3_lfsrReg_9[2] ^ tickers_x3_lfsrReg_9[3] ^
    tickers_x3_lfsrReg_9[5];
  wire [14:0] tickers_x3_lfsrReg_lo_9 = tickers_x3_lfsrReg_9[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_69 = {tickers_x3_lfsrReg_hi_9,tickers_x3_lfsrReg_lo_9};
  reg [15:0] tickers_x3_lfsrReg_10;
  wire  tickers_x3_lfsrReg_hi_10 = tickers_x3_lfsrReg_10[0] ^ tickers_x3_lfsrReg_10[2] ^ tickers_x3_lfsrReg_10[3] ^
    tickers_x3_lfsrReg_10[5];
  wire [14:0] tickers_x3_lfsrReg_lo_10 = tickers_x3_lfsrReg_10[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_76 = {tickers_x3_lfsrReg_hi_10,tickers_x3_lfsrReg_lo_10};
  reg [15:0] tickers_x3_lfsrReg_11;
  wire  tickers_x3_lfsrReg_hi_11 = tickers_x3_lfsrReg_11[0] ^ tickers_x3_lfsrReg_11[2] ^ tickers_x3_lfsrReg_11[3] ^
    tickers_x3_lfsrReg_11[5];
  wire [14:0] tickers_x3_lfsrReg_lo_11 = tickers_x3_lfsrReg_11[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_83 = {tickers_x3_lfsrReg_hi_11,tickers_x3_lfsrReg_lo_11};
  reg [15:0] tickers_x3_lfsrReg_12;
  wire  tickers_x3_lfsrReg_hi_12 = tickers_x3_lfsrReg_12[0] ^ tickers_x3_lfsrReg_12[2] ^ tickers_x3_lfsrReg_12[3] ^
    tickers_x3_lfsrReg_12[5];
  wire [14:0] tickers_x3_lfsrReg_lo_12 = tickers_x3_lfsrReg_12[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_90 = {tickers_x3_lfsrReg_hi_12,tickers_x3_lfsrReg_lo_12};
  reg [15:0] tickers_x3_lfsrReg_13;
  wire  tickers_x3_lfsrReg_hi_13 = tickers_x3_lfsrReg_13[0] ^ tickers_x3_lfsrReg_13[2] ^ tickers_x3_lfsrReg_13[3] ^
    tickers_x3_lfsrReg_13[5];
  wire [14:0] tickers_x3_lfsrReg_lo_13 = tickers_x3_lfsrReg_13[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_97 = {tickers_x3_lfsrReg_hi_13,tickers_x3_lfsrReg_lo_13};
  reg [15:0] tickers_x3_lfsrReg_14;
  wire  tickers_x3_lfsrReg_hi_14 = tickers_x3_lfsrReg_14[0] ^ tickers_x3_lfsrReg_14[2] ^ tickers_x3_lfsrReg_14[3] ^
    tickers_x3_lfsrReg_14[5];
  wire [14:0] tickers_x3_lfsrReg_lo_14 = tickers_x3_lfsrReg_14[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_104 = {tickers_x3_lfsrReg_hi_14,tickers_x3_lfsrReg_lo_14};
  reg [15:0] tickers_x3_lfsrReg_15;
  wire  tickers_x3_lfsrReg_hi_15 = tickers_x3_lfsrReg_15[0] ^ tickers_x3_lfsrReg_15[2] ^ tickers_x3_lfsrReg_15[3] ^
    tickers_x3_lfsrReg_15[5];
  wire [14:0] tickers_x3_lfsrReg_lo_15 = tickers_x3_lfsrReg_15[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_111 = {tickers_x3_lfsrReg_hi_15,tickers_x3_lfsrReg_lo_15};
  reg [15:0] tickers_x3_lfsrReg_16;
  wire  tickers_x3_lfsrReg_hi_16 = tickers_x3_lfsrReg_16[0] ^ tickers_x3_lfsrReg_16[2] ^ tickers_x3_lfsrReg_16[3] ^
    tickers_x3_lfsrReg_16[5];
  wire [14:0] tickers_x3_lfsrReg_lo_16 = tickers_x3_lfsrReg_16[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_118 = {tickers_x3_lfsrReg_hi_16,tickers_x3_lfsrReg_lo_16};
  reg [15:0] tickers_x3_lfsrReg_17;
  wire  tickers_x3_lfsrReg_hi_17 = tickers_x3_lfsrReg_17[0] ^ tickers_x3_lfsrReg_17[2] ^ tickers_x3_lfsrReg_17[3] ^
    tickers_x3_lfsrReg_17[5];
  wire [14:0] tickers_x3_lfsrReg_lo_17 = tickers_x3_lfsrReg_17[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_125 = {tickers_x3_lfsrReg_hi_17,tickers_x3_lfsrReg_lo_17};
  reg [15:0] tickers_x3_lfsrReg_18;
  wire  tickers_x3_lfsrReg_hi_18 = tickers_x3_lfsrReg_18[0] ^ tickers_x3_lfsrReg_18[2] ^ tickers_x3_lfsrReg_18[3] ^
    tickers_x3_lfsrReg_18[5];
  wire [14:0] tickers_x3_lfsrReg_lo_18 = tickers_x3_lfsrReg_18[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_132 = {tickers_x3_lfsrReg_hi_18,tickers_x3_lfsrReg_lo_18};
  reg [15:0] tickers_x3_lfsrReg_19;
  wire  tickers_x3_lfsrReg_hi_19 = tickers_x3_lfsrReg_19[0] ^ tickers_x3_lfsrReg_19[2] ^ tickers_x3_lfsrReg_19[3] ^
    tickers_x3_lfsrReg_19[5];
  wire [14:0] tickers_x3_lfsrReg_lo_19 = tickers_x3_lfsrReg_19[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_139 = {tickers_x3_lfsrReg_hi_19,tickers_x3_lfsrReg_lo_19};
  reg [15:0] tickers_x3_lfsrReg_20;
  wire  tickers_x3_lfsrReg_hi_20 = tickers_x3_lfsrReg_20[0] ^ tickers_x3_lfsrReg_20[2] ^ tickers_x3_lfsrReg_20[3] ^
    tickers_x3_lfsrReg_20[5];
  wire [14:0] tickers_x3_lfsrReg_lo_20 = tickers_x3_lfsrReg_20[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_146 = {tickers_x3_lfsrReg_hi_20,tickers_x3_lfsrReg_lo_20};
  reg [15:0] tickers_x3_lfsrReg_21;
  wire  tickers_x3_lfsrReg_hi_21 = tickers_x3_lfsrReg_21[0] ^ tickers_x3_lfsrReg_21[2] ^ tickers_x3_lfsrReg_21[3] ^
    tickers_x3_lfsrReg_21[5];
  wire [14:0] tickers_x3_lfsrReg_lo_21 = tickers_x3_lfsrReg_21[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_153 = {tickers_x3_lfsrReg_hi_21,tickers_x3_lfsrReg_lo_21};
  reg [15:0] tickers_x3_lfsrReg_22;
  wire  tickers_x3_lfsrReg_hi_22 = tickers_x3_lfsrReg_22[0] ^ tickers_x3_lfsrReg_22[2] ^ tickers_x3_lfsrReg_22[3] ^
    tickers_x3_lfsrReg_22[5];
  wire [14:0] tickers_x3_lfsrReg_lo_22 = tickers_x3_lfsrReg_22[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_160 = {tickers_x3_lfsrReg_hi_22,tickers_x3_lfsrReg_lo_22};
  reg [15:0] tickers_x3_lfsrReg_23;
  wire  tickers_x3_lfsrReg_hi_23 = tickers_x3_lfsrReg_23[0] ^ tickers_x3_lfsrReg_23[2] ^ tickers_x3_lfsrReg_23[3] ^
    tickers_x3_lfsrReg_23[5];
  wire [14:0] tickers_x3_lfsrReg_lo_23 = tickers_x3_lfsrReg_23[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_167 = {tickers_x3_lfsrReg_hi_23,tickers_x3_lfsrReg_lo_23};
  reg [15:0] tickers_x3_lfsrReg_24;
  wire  tickers_x3_lfsrReg_hi_24 = tickers_x3_lfsrReg_24[0] ^ tickers_x3_lfsrReg_24[2] ^ tickers_x3_lfsrReg_24[3] ^
    tickers_x3_lfsrReg_24[5];
  wire [14:0] tickers_x3_lfsrReg_lo_24 = tickers_x3_lfsrReg_24[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_174 = {tickers_x3_lfsrReg_hi_24,tickers_x3_lfsrReg_lo_24};
  reg [15:0] tickers_x3_lfsrReg_25;
  wire  tickers_x3_lfsrReg_hi_25 = tickers_x3_lfsrReg_25[0] ^ tickers_x3_lfsrReg_25[2] ^ tickers_x3_lfsrReg_25[3] ^
    tickers_x3_lfsrReg_25[5];
  wire [14:0] tickers_x3_lfsrReg_lo_25 = tickers_x3_lfsrReg_25[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_181 = {tickers_x3_lfsrReg_hi_25,tickers_x3_lfsrReg_lo_25};
  reg [15:0] tickers_x3_lfsrReg_26;
  wire  tickers_x3_lfsrReg_hi_26 = tickers_x3_lfsrReg_26[0] ^ tickers_x3_lfsrReg_26[2] ^ tickers_x3_lfsrReg_26[3] ^
    tickers_x3_lfsrReg_26[5];
  wire [14:0] tickers_x3_lfsrReg_lo_26 = tickers_x3_lfsrReg_26[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_188 = {tickers_x3_lfsrReg_hi_26,tickers_x3_lfsrReg_lo_26};
  reg [15:0] tickers_x3_lfsrReg_27;
  wire  tickers_x3_lfsrReg_hi_27 = tickers_x3_lfsrReg_27[0] ^ tickers_x3_lfsrReg_27[2] ^ tickers_x3_lfsrReg_27[3] ^
    tickers_x3_lfsrReg_27[5];
  wire [14:0] tickers_x3_lfsrReg_lo_27 = tickers_x3_lfsrReg_27[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_195 = {tickers_x3_lfsrReg_hi_27,tickers_x3_lfsrReg_lo_27};
  reg [15:0] tickers_x3_lfsrReg_28;
  wire  tickers_x3_lfsrReg_hi_28 = tickers_x3_lfsrReg_28[0] ^ tickers_x3_lfsrReg_28[2] ^ tickers_x3_lfsrReg_28[3] ^
    tickers_x3_lfsrReg_28[5];
  wire [14:0] tickers_x3_lfsrReg_lo_28 = tickers_x3_lfsrReg_28[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_202 = {tickers_x3_lfsrReg_hi_28,tickers_x3_lfsrReg_lo_28};
  reg [15:0] tickers_x3_lfsrReg_29;
  wire  tickers_x3_lfsrReg_hi_29 = tickers_x3_lfsrReg_29[0] ^ tickers_x3_lfsrReg_29[2] ^ tickers_x3_lfsrReg_29[3] ^
    tickers_x3_lfsrReg_29[5];
  wire [14:0] tickers_x3_lfsrReg_lo_29 = tickers_x3_lfsrReg_29[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_209 = {tickers_x3_lfsrReg_hi_29,tickers_x3_lfsrReg_lo_29};
  reg [15:0] tickers_x3_lfsrReg_30;
  wire  tickers_x3_lfsrReg_hi_30 = tickers_x3_lfsrReg_30[0] ^ tickers_x3_lfsrReg_30[2] ^ tickers_x3_lfsrReg_30[3] ^
    tickers_x3_lfsrReg_30[5];
  wire [14:0] tickers_x3_lfsrReg_lo_30 = tickers_x3_lfsrReg_30[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_216 = {tickers_x3_lfsrReg_hi_30,tickers_x3_lfsrReg_lo_30};
  reg [15:0] tickers_x3_lfsrReg_31;
  wire  tickers_x3_lfsrReg_hi_31 = tickers_x3_lfsrReg_31[0] ^ tickers_x3_lfsrReg_31[2] ^ tickers_x3_lfsrReg_31[3] ^
    tickers_x3_lfsrReg_31[5];
  wire [14:0] tickers_x3_lfsrReg_lo_31 = tickers_x3_lfsrReg_31[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_223 = {tickers_x3_lfsrReg_hi_31,tickers_x3_lfsrReg_lo_31};
  reg [15:0] tickers_x3_lfsrReg_32;
  wire  tickers_x3_lfsrReg_hi_32 = tickers_x3_lfsrReg_32[0] ^ tickers_x3_lfsrReg_32[2] ^ tickers_x3_lfsrReg_32[3] ^
    tickers_x3_lfsrReg_32[5];
  wire [14:0] tickers_x3_lfsrReg_lo_32 = tickers_x3_lfsrReg_32[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_230 = {tickers_x3_lfsrReg_hi_32,tickers_x3_lfsrReg_lo_32};
  reg [15:0] tickers_x3_lfsrReg_33;
  wire  tickers_x3_lfsrReg_hi_33 = tickers_x3_lfsrReg_33[0] ^ tickers_x3_lfsrReg_33[2] ^ tickers_x3_lfsrReg_33[3] ^
    tickers_x3_lfsrReg_33[5];
  wire [14:0] tickers_x3_lfsrReg_lo_33 = tickers_x3_lfsrReg_33[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_237 = {tickers_x3_lfsrReg_hi_33,tickers_x3_lfsrReg_lo_33};
  reg [15:0] tickers_x3_lfsrReg_34;
  wire  tickers_x3_lfsrReg_hi_34 = tickers_x3_lfsrReg_34[0] ^ tickers_x3_lfsrReg_34[2] ^ tickers_x3_lfsrReg_34[3] ^
    tickers_x3_lfsrReg_34[5];
  wire [14:0] tickers_x3_lfsrReg_lo_34 = tickers_x3_lfsrReg_34[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_244 = {tickers_x3_lfsrReg_hi_34,tickers_x3_lfsrReg_lo_34};
  reg [15:0] tickers_x3_lfsrReg_35;
  wire  tickers_x3_lfsrReg_hi_35 = tickers_x3_lfsrReg_35[0] ^ tickers_x3_lfsrReg_35[2] ^ tickers_x3_lfsrReg_35[3] ^
    tickers_x3_lfsrReg_35[5];
  wire [14:0] tickers_x3_lfsrReg_lo_35 = tickers_x3_lfsrReg_35[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_251 = {tickers_x3_lfsrReg_hi_35,tickers_x3_lfsrReg_lo_35};
  reg [15:0] tickers_x3_lfsrReg_36;
  wire  tickers_x3_lfsrReg_hi_36 = tickers_x3_lfsrReg_36[0] ^ tickers_x3_lfsrReg_36[2] ^ tickers_x3_lfsrReg_36[3] ^
    tickers_x3_lfsrReg_36[5];
  wire [14:0] tickers_x3_lfsrReg_lo_36 = tickers_x3_lfsrReg_36[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_258 = {tickers_x3_lfsrReg_hi_36,tickers_x3_lfsrReg_lo_36};
  reg [15:0] tickers_x3_lfsrReg_37;
  wire  tickers_x3_lfsrReg_hi_37 = tickers_x3_lfsrReg_37[0] ^ tickers_x3_lfsrReg_37[2] ^ tickers_x3_lfsrReg_37[3] ^
    tickers_x3_lfsrReg_37[5];
  wire [14:0] tickers_x3_lfsrReg_lo_37 = tickers_x3_lfsrReg_37[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_265 = {tickers_x3_lfsrReg_hi_37,tickers_x3_lfsrReg_lo_37};
  reg [15:0] tickers_x3_lfsrReg_38;
  wire  tickers_x3_lfsrReg_hi_38 = tickers_x3_lfsrReg_38[0] ^ tickers_x3_lfsrReg_38[2] ^ tickers_x3_lfsrReg_38[3] ^
    tickers_x3_lfsrReg_38[5];
  wire [14:0] tickers_x3_lfsrReg_lo_38 = tickers_x3_lfsrReg_38[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_272 = {tickers_x3_lfsrReg_hi_38,tickers_x3_lfsrReg_lo_38};
  reg [15:0] tickers_x3_lfsrReg_39;
  wire  tickers_x3_lfsrReg_hi_39 = tickers_x3_lfsrReg_39[0] ^ tickers_x3_lfsrReg_39[2] ^ tickers_x3_lfsrReg_39[3] ^
    tickers_x3_lfsrReg_39[5];
  wire [14:0] tickers_x3_lfsrReg_lo_39 = tickers_x3_lfsrReg_39[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_279 = {tickers_x3_lfsrReg_hi_39,tickers_x3_lfsrReg_lo_39};
  reg [15:0] tickers_x3_lfsrReg_40;
  wire  tickers_x3_lfsrReg_hi_40 = tickers_x3_lfsrReg_40[0] ^ tickers_x3_lfsrReg_40[2] ^ tickers_x3_lfsrReg_40[3] ^
    tickers_x3_lfsrReg_40[5];
  wire [14:0] tickers_x3_lfsrReg_lo_40 = tickers_x3_lfsrReg_40[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_286 = {tickers_x3_lfsrReg_hi_40,tickers_x3_lfsrReg_lo_40};
  reg [15:0] tickers_x3_lfsrReg_41;
  wire  tickers_x3_lfsrReg_hi_41 = tickers_x3_lfsrReg_41[0] ^ tickers_x3_lfsrReg_41[2] ^ tickers_x3_lfsrReg_41[3] ^
    tickers_x3_lfsrReg_41[5];
  wire [14:0] tickers_x3_lfsrReg_lo_41 = tickers_x3_lfsrReg_41[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_293 = {tickers_x3_lfsrReg_hi_41,tickers_x3_lfsrReg_lo_41};
  reg [15:0] tickers_x3_lfsrReg_42;
  wire  tickers_x3_lfsrReg_hi_42 = tickers_x3_lfsrReg_42[0] ^ tickers_x3_lfsrReg_42[2] ^ tickers_x3_lfsrReg_42[3] ^
    tickers_x3_lfsrReg_42[5];
  wire [14:0] tickers_x3_lfsrReg_lo_42 = tickers_x3_lfsrReg_42[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_300 = {tickers_x3_lfsrReg_hi_42,tickers_x3_lfsrReg_lo_42};
  reg [15:0] tickers_x3_lfsrReg_43;
  wire  tickers_x3_lfsrReg_hi_43 = tickers_x3_lfsrReg_43[0] ^ tickers_x3_lfsrReg_43[2] ^ tickers_x3_lfsrReg_43[3] ^
    tickers_x3_lfsrReg_43[5];
  wire [14:0] tickers_x3_lfsrReg_lo_43 = tickers_x3_lfsrReg_43[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_307 = {tickers_x3_lfsrReg_hi_43,tickers_x3_lfsrReg_lo_43};
  reg [15:0] tickers_x3_lfsrReg_44;
  wire  tickers_x3_lfsrReg_hi_44 = tickers_x3_lfsrReg_44[0] ^ tickers_x3_lfsrReg_44[2] ^ tickers_x3_lfsrReg_44[3] ^
    tickers_x3_lfsrReg_44[5];
  wire [14:0] tickers_x3_lfsrReg_lo_44 = tickers_x3_lfsrReg_44[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_314 = {tickers_x3_lfsrReg_hi_44,tickers_x3_lfsrReg_lo_44};
  reg [15:0] tickers_x3_lfsrReg_45;
  wire  tickers_x3_lfsrReg_hi_45 = tickers_x3_lfsrReg_45[0] ^ tickers_x3_lfsrReg_45[2] ^ tickers_x3_lfsrReg_45[3] ^
    tickers_x3_lfsrReg_45[5];
  wire [14:0] tickers_x3_lfsrReg_lo_45 = tickers_x3_lfsrReg_45[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_321 = {tickers_x3_lfsrReg_hi_45,tickers_x3_lfsrReg_lo_45};
  reg [15:0] tickers_x3_lfsrReg_46;
  wire  tickers_x3_lfsrReg_hi_46 = tickers_x3_lfsrReg_46[0] ^ tickers_x3_lfsrReg_46[2] ^ tickers_x3_lfsrReg_46[3] ^
    tickers_x3_lfsrReg_46[5];
  wire [14:0] tickers_x3_lfsrReg_lo_46 = tickers_x3_lfsrReg_46[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_328 = {tickers_x3_lfsrReg_hi_46,tickers_x3_lfsrReg_lo_46};
  reg [15:0] tickers_x3_lfsrReg_47;
  wire  tickers_x3_lfsrReg_hi_47 = tickers_x3_lfsrReg_47[0] ^ tickers_x3_lfsrReg_47[2] ^ tickers_x3_lfsrReg_47[3] ^
    tickers_x3_lfsrReg_47[5];
  wire [14:0] tickers_x3_lfsrReg_lo_47 = tickers_x3_lfsrReg_47[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_335 = {tickers_x3_lfsrReg_hi_47,tickers_x3_lfsrReg_lo_47};
  reg [15:0] tickers_x3_lfsrReg_48;
  wire  tickers_x3_lfsrReg_hi_48 = tickers_x3_lfsrReg_48[0] ^ tickers_x3_lfsrReg_48[2] ^ tickers_x3_lfsrReg_48[3] ^
    tickers_x3_lfsrReg_48[5];
  wire [14:0] tickers_x3_lfsrReg_lo_48 = tickers_x3_lfsrReg_48[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_342 = {tickers_x3_lfsrReg_hi_48,tickers_x3_lfsrReg_lo_48};
  reg [15:0] tickers_x3_lfsrReg_49;
  wire  tickers_x3_lfsrReg_hi_49 = tickers_x3_lfsrReg_49[0] ^ tickers_x3_lfsrReg_49[2] ^ tickers_x3_lfsrReg_49[3] ^
    tickers_x3_lfsrReg_49[5];
  wire [14:0] tickers_x3_lfsrReg_lo_49 = tickers_x3_lfsrReg_49[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_349 = {tickers_x3_lfsrReg_hi_49,tickers_x3_lfsrReg_lo_49};
  reg [15:0] tickers_x3_lfsrReg_50;
  wire  tickers_x3_lfsrReg_hi_50 = tickers_x3_lfsrReg_50[0] ^ tickers_x3_lfsrReg_50[2] ^ tickers_x3_lfsrReg_50[3] ^
    tickers_x3_lfsrReg_50[5];
  wire [14:0] tickers_x3_lfsrReg_lo_50 = tickers_x3_lfsrReg_50[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_356 = {tickers_x3_lfsrReg_hi_50,tickers_x3_lfsrReg_lo_50};
  reg [15:0] tickers_x3_lfsrReg_51;
  wire  tickers_x3_lfsrReg_hi_51 = tickers_x3_lfsrReg_51[0] ^ tickers_x3_lfsrReg_51[2] ^ tickers_x3_lfsrReg_51[3] ^
    tickers_x3_lfsrReg_51[5];
  wire [14:0] tickers_x3_lfsrReg_lo_51 = tickers_x3_lfsrReg_51[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_363 = {tickers_x3_lfsrReg_hi_51,tickers_x3_lfsrReg_lo_51};
  reg [15:0] tickers_x3_lfsrReg_52;
  wire  tickers_x3_lfsrReg_hi_52 = tickers_x3_lfsrReg_52[0] ^ tickers_x3_lfsrReg_52[2] ^ tickers_x3_lfsrReg_52[3] ^
    tickers_x3_lfsrReg_52[5];
  wire [14:0] tickers_x3_lfsrReg_lo_52 = tickers_x3_lfsrReg_52[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_370 = {tickers_x3_lfsrReg_hi_52,tickers_x3_lfsrReg_lo_52};
  reg [15:0] tickers_x3_lfsrReg_53;
  wire  tickers_x3_lfsrReg_hi_53 = tickers_x3_lfsrReg_53[0] ^ tickers_x3_lfsrReg_53[2] ^ tickers_x3_lfsrReg_53[3] ^
    tickers_x3_lfsrReg_53[5];
  wire [14:0] tickers_x3_lfsrReg_lo_53 = tickers_x3_lfsrReg_53[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_377 = {tickers_x3_lfsrReg_hi_53,tickers_x3_lfsrReg_lo_53};
  reg [15:0] tickers_x3_lfsrReg_54;
  wire  tickers_x3_lfsrReg_hi_54 = tickers_x3_lfsrReg_54[0] ^ tickers_x3_lfsrReg_54[2] ^ tickers_x3_lfsrReg_54[3] ^
    tickers_x3_lfsrReg_54[5];
  wire [14:0] tickers_x3_lfsrReg_lo_54 = tickers_x3_lfsrReg_54[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_384 = {tickers_x3_lfsrReg_hi_54,tickers_x3_lfsrReg_lo_54};
  reg [15:0] tickers_x3_lfsrReg_55;
  wire  tickers_x3_lfsrReg_hi_55 = tickers_x3_lfsrReg_55[0] ^ tickers_x3_lfsrReg_55[2] ^ tickers_x3_lfsrReg_55[3] ^
    tickers_x3_lfsrReg_55[5];
  wire [14:0] tickers_x3_lfsrReg_lo_55 = tickers_x3_lfsrReg_55[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_391 = {tickers_x3_lfsrReg_hi_55,tickers_x3_lfsrReg_lo_55};
  reg [15:0] tickers_x3_lfsrReg_56;
  wire  tickers_x3_lfsrReg_hi_56 = tickers_x3_lfsrReg_56[0] ^ tickers_x3_lfsrReg_56[2] ^ tickers_x3_lfsrReg_56[3] ^
    tickers_x3_lfsrReg_56[5];
  wire [14:0] tickers_x3_lfsrReg_lo_56 = tickers_x3_lfsrReg_56[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_398 = {tickers_x3_lfsrReg_hi_56,tickers_x3_lfsrReg_lo_56};
  reg [15:0] tickers_x3_lfsrReg_57;
  wire  tickers_x3_lfsrReg_hi_57 = tickers_x3_lfsrReg_57[0] ^ tickers_x3_lfsrReg_57[2] ^ tickers_x3_lfsrReg_57[3] ^
    tickers_x3_lfsrReg_57[5];
  wire [14:0] tickers_x3_lfsrReg_lo_57 = tickers_x3_lfsrReg_57[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_405 = {tickers_x3_lfsrReg_hi_57,tickers_x3_lfsrReg_lo_57};
  reg [15:0] tickers_x3_lfsrReg_58;
  wire  tickers_x3_lfsrReg_hi_58 = tickers_x3_lfsrReg_58[0] ^ tickers_x3_lfsrReg_58[2] ^ tickers_x3_lfsrReg_58[3] ^
    tickers_x3_lfsrReg_58[5];
  wire [14:0] tickers_x3_lfsrReg_lo_58 = tickers_x3_lfsrReg_58[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_412 = {tickers_x3_lfsrReg_hi_58,tickers_x3_lfsrReg_lo_58};
  reg [15:0] tickers_x3_lfsrReg_59;
  wire  tickers_x3_lfsrReg_hi_59 = tickers_x3_lfsrReg_59[0] ^ tickers_x3_lfsrReg_59[2] ^ tickers_x3_lfsrReg_59[3] ^
    tickers_x3_lfsrReg_59[5];
  wire [14:0] tickers_x3_lfsrReg_lo_59 = tickers_x3_lfsrReg_59[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_419 = {tickers_x3_lfsrReg_hi_59,tickers_x3_lfsrReg_lo_59};
  reg [15:0] tickers_x3_lfsrReg_60;
  wire  tickers_x3_lfsrReg_hi_60 = tickers_x3_lfsrReg_60[0] ^ tickers_x3_lfsrReg_60[2] ^ tickers_x3_lfsrReg_60[3] ^
    tickers_x3_lfsrReg_60[5];
  wire [14:0] tickers_x3_lfsrReg_lo_60 = tickers_x3_lfsrReg_60[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_426 = {tickers_x3_lfsrReg_hi_60,tickers_x3_lfsrReg_lo_60};
  reg [15:0] tickers_x3_lfsrReg_61;
  wire  tickers_x3_lfsrReg_hi_61 = tickers_x3_lfsrReg_61[0] ^ tickers_x3_lfsrReg_61[2] ^ tickers_x3_lfsrReg_61[3] ^
    tickers_x3_lfsrReg_61[5];
  wire [14:0] tickers_x3_lfsrReg_lo_61 = tickers_x3_lfsrReg_61[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_433 = {tickers_x3_lfsrReg_hi_61,tickers_x3_lfsrReg_lo_61};
  reg [15:0] tickers_x3_lfsrReg_62;
  wire  tickers_x3_lfsrReg_hi_62 = tickers_x3_lfsrReg_62[0] ^ tickers_x3_lfsrReg_62[2] ^ tickers_x3_lfsrReg_62[3] ^
    tickers_x3_lfsrReg_62[5];
  wire [14:0] tickers_x3_lfsrReg_lo_62 = tickers_x3_lfsrReg_62[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_440 = {tickers_x3_lfsrReg_hi_62,tickers_x3_lfsrReg_lo_62};
  reg [15:0] tickers_x3_lfsrReg_63;
  wire  tickers_x3_lfsrReg_hi_63 = tickers_x3_lfsrReg_63[0] ^ tickers_x3_lfsrReg_63[2] ^ tickers_x3_lfsrReg_63[3] ^
    tickers_x3_lfsrReg_63[5];
  wire [14:0] tickers_x3_lfsrReg_lo_63 = tickers_x3_lfsrReg_63[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_447 = {tickers_x3_lfsrReg_hi_63,tickers_x3_lfsrReg_lo_63};
  reg [15:0] tickers_x3_lfsrReg_64;
  wire  tickers_x3_lfsrReg_hi_64 = tickers_x3_lfsrReg_64[0] ^ tickers_x3_lfsrReg_64[2] ^ tickers_x3_lfsrReg_64[3] ^
    tickers_x3_lfsrReg_64[5];
  wire [14:0] tickers_x3_lfsrReg_lo_64 = tickers_x3_lfsrReg_64[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_454 = {tickers_x3_lfsrReg_hi_64,tickers_x3_lfsrReg_lo_64};
  reg [15:0] tickers_x3_lfsrReg_65;
  wire  tickers_x3_lfsrReg_hi_65 = tickers_x3_lfsrReg_65[0] ^ tickers_x3_lfsrReg_65[2] ^ tickers_x3_lfsrReg_65[3] ^
    tickers_x3_lfsrReg_65[5];
  wire [14:0] tickers_x3_lfsrReg_lo_65 = tickers_x3_lfsrReg_65[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_461 = {tickers_x3_lfsrReg_hi_65,tickers_x3_lfsrReg_lo_65};
  reg [15:0] tickers_x3_lfsrReg_66;
  wire  tickers_x3_lfsrReg_hi_66 = tickers_x3_lfsrReg_66[0] ^ tickers_x3_lfsrReg_66[2] ^ tickers_x3_lfsrReg_66[3] ^
    tickers_x3_lfsrReg_66[5];
  wire [14:0] tickers_x3_lfsrReg_lo_66 = tickers_x3_lfsrReg_66[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_468 = {tickers_x3_lfsrReg_hi_66,tickers_x3_lfsrReg_lo_66};
  reg [15:0] tickers_x3_lfsrReg_67;
  wire  tickers_x3_lfsrReg_hi_67 = tickers_x3_lfsrReg_67[0] ^ tickers_x3_lfsrReg_67[2] ^ tickers_x3_lfsrReg_67[3] ^
    tickers_x3_lfsrReg_67[5];
  wire [14:0] tickers_x3_lfsrReg_lo_67 = tickers_x3_lfsrReg_67[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_475 = {tickers_x3_lfsrReg_hi_67,tickers_x3_lfsrReg_lo_67};
  reg [15:0] tickers_x3_lfsrReg_68;
  wire  tickers_x3_lfsrReg_hi_68 = tickers_x3_lfsrReg_68[0] ^ tickers_x3_lfsrReg_68[2] ^ tickers_x3_lfsrReg_68[3] ^
    tickers_x3_lfsrReg_68[5];
  wire [14:0] tickers_x3_lfsrReg_lo_68 = tickers_x3_lfsrReg_68[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_482 = {tickers_x3_lfsrReg_hi_68,tickers_x3_lfsrReg_lo_68};
  reg [15:0] tickers_x3_lfsrReg_69;
  wire  tickers_x3_lfsrReg_hi_69 = tickers_x3_lfsrReg_69[0] ^ tickers_x3_lfsrReg_69[2] ^ tickers_x3_lfsrReg_69[3] ^
    tickers_x3_lfsrReg_69[5];
  wire [14:0] tickers_x3_lfsrReg_lo_69 = tickers_x3_lfsrReg_69[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_489 = {tickers_x3_lfsrReg_hi_69,tickers_x3_lfsrReg_lo_69};
  reg [15:0] tickers_x3_lfsrReg_70;
  wire  tickers_x3_lfsrReg_hi_70 = tickers_x3_lfsrReg_70[0] ^ tickers_x3_lfsrReg_70[2] ^ tickers_x3_lfsrReg_70[3] ^
    tickers_x3_lfsrReg_70[5];
  wire [14:0] tickers_x3_lfsrReg_lo_70 = tickers_x3_lfsrReg_70[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_496 = {tickers_x3_lfsrReg_hi_70,tickers_x3_lfsrReg_lo_70};
  reg [15:0] tickers_x3_lfsrReg_71;
  wire  tickers_x3_lfsrReg_hi_71 = tickers_x3_lfsrReg_71[0] ^ tickers_x3_lfsrReg_71[2] ^ tickers_x3_lfsrReg_71[3] ^
    tickers_x3_lfsrReg_71[5];
  wire [14:0] tickers_x3_lfsrReg_lo_71 = tickers_x3_lfsrReg_71[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_503 = {tickers_x3_lfsrReg_hi_71,tickers_x3_lfsrReg_lo_71};
  reg [15:0] tickers_x3_lfsrReg_72;
  wire  tickers_x3_lfsrReg_hi_72 = tickers_x3_lfsrReg_72[0] ^ tickers_x3_lfsrReg_72[2] ^ tickers_x3_lfsrReg_72[3] ^
    tickers_x3_lfsrReg_72[5];
  wire [14:0] tickers_x3_lfsrReg_lo_72 = tickers_x3_lfsrReg_72[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_510 = {tickers_x3_lfsrReg_hi_72,tickers_x3_lfsrReg_lo_72};
  reg [15:0] tickers_x3_lfsrReg_73;
  wire  tickers_x3_lfsrReg_hi_73 = tickers_x3_lfsrReg_73[0] ^ tickers_x3_lfsrReg_73[2] ^ tickers_x3_lfsrReg_73[3] ^
    tickers_x3_lfsrReg_73[5];
  wire [14:0] tickers_x3_lfsrReg_lo_73 = tickers_x3_lfsrReg_73[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_517 = {tickers_x3_lfsrReg_hi_73,tickers_x3_lfsrReg_lo_73};
  reg [15:0] tickers_x3_lfsrReg_74;
  wire  tickers_x3_lfsrReg_hi_74 = tickers_x3_lfsrReg_74[0] ^ tickers_x3_lfsrReg_74[2] ^ tickers_x3_lfsrReg_74[3] ^
    tickers_x3_lfsrReg_74[5];
  wire [14:0] tickers_x3_lfsrReg_lo_74 = tickers_x3_lfsrReg_74[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_524 = {tickers_x3_lfsrReg_hi_74,tickers_x3_lfsrReg_lo_74};
  reg [15:0] tickers_x3_lfsrReg_75;
  wire  tickers_x3_lfsrReg_hi_75 = tickers_x3_lfsrReg_75[0] ^ tickers_x3_lfsrReg_75[2] ^ tickers_x3_lfsrReg_75[3] ^
    tickers_x3_lfsrReg_75[5];
  wire [14:0] tickers_x3_lfsrReg_lo_75 = tickers_x3_lfsrReg_75[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_531 = {tickers_x3_lfsrReg_hi_75,tickers_x3_lfsrReg_lo_75};
  reg [15:0] tickers_x3_lfsrReg_76;
  wire  tickers_x3_lfsrReg_hi_76 = tickers_x3_lfsrReg_76[0] ^ tickers_x3_lfsrReg_76[2] ^ tickers_x3_lfsrReg_76[3] ^
    tickers_x3_lfsrReg_76[5];
  wire [14:0] tickers_x3_lfsrReg_lo_76 = tickers_x3_lfsrReg_76[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_538 = {tickers_x3_lfsrReg_hi_76,tickers_x3_lfsrReg_lo_76};
  reg [15:0] tickers_x3_lfsrReg_77;
  wire  tickers_x3_lfsrReg_hi_77 = tickers_x3_lfsrReg_77[0] ^ tickers_x3_lfsrReg_77[2] ^ tickers_x3_lfsrReg_77[3] ^
    tickers_x3_lfsrReg_77[5];
  wire [14:0] tickers_x3_lfsrReg_lo_77 = tickers_x3_lfsrReg_77[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_545 = {tickers_x3_lfsrReg_hi_77,tickers_x3_lfsrReg_lo_77};
  reg [15:0] tickers_x3_lfsrReg_78;
  wire  tickers_x3_lfsrReg_hi_78 = tickers_x3_lfsrReg_78[0] ^ tickers_x3_lfsrReg_78[2] ^ tickers_x3_lfsrReg_78[3] ^
    tickers_x3_lfsrReg_78[5];
  wire [14:0] tickers_x3_lfsrReg_lo_78 = tickers_x3_lfsrReg_78[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_552 = {tickers_x3_lfsrReg_hi_78,tickers_x3_lfsrReg_lo_78};
  reg [15:0] tickers_x3_lfsrReg_79;
  wire  tickers_x3_lfsrReg_hi_79 = tickers_x3_lfsrReg_79[0] ^ tickers_x3_lfsrReg_79[2] ^ tickers_x3_lfsrReg_79[3] ^
    tickers_x3_lfsrReg_79[5];
  wire [14:0] tickers_x3_lfsrReg_lo_79 = tickers_x3_lfsrReg_79[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_559 = {tickers_x3_lfsrReg_hi_79,tickers_x3_lfsrReg_lo_79};
  reg [15:0] tickers_x3_lfsrReg_80;
  wire  tickers_x3_lfsrReg_hi_80 = tickers_x3_lfsrReg_80[0] ^ tickers_x3_lfsrReg_80[2] ^ tickers_x3_lfsrReg_80[3] ^
    tickers_x3_lfsrReg_80[5];
  wire [14:0] tickers_x3_lfsrReg_lo_80 = tickers_x3_lfsrReg_80[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_566 = {tickers_x3_lfsrReg_hi_80,tickers_x3_lfsrReg_lo_80};
  reg [15:0] tickers_x3_lfsrReg_81;
  wire  tickers_x3_lfsrReg_hi_81 = tickers_x3_lfsrReg_81[0] ^ tickers_x3_lfsrReg_81[2] ^ tickers_x3_lfsrReg_81[3] ^
    tickers_x3_lfsrReg_81[5];
  wire [14:0] tickers_x3_lfsrReg_lo_81 = tickers_x3_lfsrReg_81[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_573 = {tickers_x3_lfsrReg_hi_81,tickers_x3_lfsrReg_lo_81};
  reg [15:0] tickers_x3_lfsrReg_82;
  wire  tickers_x3_lfsrReg_hi_82 = tickers_x3_lfsrReg_82[0] ^ tickers_x3_lfsrReg_82[2] ^ tickers_x3_lfsrReg_82[3] ^
    tickers_x3_lfsrReg_82[5];
  wire [14:0] tickers_x3_lfsrReg_lo_82 = tickers_x3_lfsrReg_82[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_580 = {tickers_x3_lfsrReg_hi_82,tickers_x3_lfsrReg_lo_82};
  reg [15:0] tickers_x3_lfsrReg_83;
  wire  tickers_x3_lfsrReg_hi_83 = tickers_x3_lfsrReg_83[0] ^ tickers_x3_lfsrReg_83[2] ^ tickers_x3_lfsrReg_83[3] ^
    tickers_x3_lfsrReg_83[5];
  wire [14:0] tickers_x3_lfsrReg_lo_83 = tickers_x3_lfsrReg_83[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_587 = {tickers_x3_lfsrReg_hi_83,tickers_x3_lfsrReg_lo_83};
  reg [15:0] tickers_x3_lfsrReg_84;
  wire  tickers_x3_lfsrReg_hi_84 = tickers_x3_lfsrReg_84[0] ^ tickers_x3_lfsrReg_84[2] ^ tickers_x3_lfsrReg_84[3] ^
    tickers_x3_lfsrReg_84[5];
  wire [14:0] tickers_x3_lfsrReg_lo_84 = tickers_x3_lfsrReg_84[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_594 = {tickers_x3_lfsrReg_hi_84,tickers_x3_lfsrReg_lo_84};
  reg [15:0] tickers_x3_lfsrReg_85;
  wire  tickers_x3_lfsrReg_hi_85 = tickers_x3_lfsrReg_85[0] ^ tickers_x3_lfsrReg_85[2] ^ tickers_x3_lfsrReg_85[3] ^
    tickers_x3_lfsrReg_85[5];
  wire [14:0] tickers_x3_lfsrReg_lo_85 = tickers_x3_lfsrReg_85[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_601 = {tickers_x3_lfsrReg_hi_85,tickers_x3_lfsrReg_lo_85};
  reg [15:0] tickers_x3_lfsrReg_86;
  wire  tickers_x3_lfsrReg_hi_86 = tickers_x3_lfsrReg_86[0] ^ tickers_x3_lfsrReg_86[2] ^ tickers_x3_lfsrReg_86[3] ^
    tickers_x3_lfsrReg_86[5];
  wire [14:0] tickers_x3_lfsrReg_lo_86 = tickers_x3_lfsrReg_86[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_608 = {tickers_x3_lfsrReg_hi_86,tickers_x3_lfsrReg_lo_86};
  reg [15:0] tickers_x3_lfsrReg_87;
  wire  tickers_x3_lfsrReg_hi_87 = tickers_x3_lfsrReg_87[0] ^ tickers_x3_lfsrReg_87[2] ^ tickers_x3_lfsrReg_87[3] ^
    tickers_x3_lfsrReg_87[5];
  wire [14:0] tickers_x3_lfsrReg_lo_87 = tickers_x3_lfsrReg_87[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_615 = {tickers_x3_lfsrReg_hi_87,tickers_x3_lfsrReg_lo_87};
  reg [15:0] tickers_x3_lfsrReg_88;
  wire  tickers_x3_lfsrReg_hi_88 = tickers_x3_lfsrReg_88[0] ^ tickers_x3_lfsrReg_88[2] ^ tickers_x3_lfsrReg_88[3] ^
    tickers_x3_lfsrReg_88[5];
  wire [14:0] tickers_x3_lfsrReg_lo_88 = tickers_x3_lfsrReg_88[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_622 = {tickers_x3_lfsrReg_hi_88,tickers_x3_lfsrReg_lo_88};
  reg [15:0] tickers_x3_lfsrReg_89;
  wire  tickers_x3_lfsrReg_hi_89 = tickers_x3_lfsrReg_89[0] ^ tickers_x3_lfsrReg_89[2] ^ tickers_x3_lfsrReg_89[3] ^
    tickers_x3_lfsrReg_89[5];
  wire [14:0] tickers_x3_lfsrReg_lo_89 = tickers_x3_lfsrReg_89[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_629 = {tickers_x3_lfsrReg_hi_89,tickers_x3_lfsrReg_lo_89};
  reg [15:0] tickers_x3_lfsrReg_90;
  wire  tickers_x3_lfsrReg_hi_90 = tickers_x3_lfsrReg_90[0] ^ tickers_x3_lfsrReg_90[2] ^ tickers_x3_lfsrReg_90[3] ^
    tickers_x3_lfsrReg_90[5];
  wire [14:0] tickers_x3_lfsrReg_lo_90 = tickers_x3_lfsrReg_90[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_636 = {tickers_x3_lfsrReg_hi_90,tickers_x3_lfsrReg_lo_90};
  reg [15:0] tickers_x3_lfsrReg_91;
  wire  tickers_x3_lfsrReg_hi_91 = tickers_x3_lfsrReg_91[0] ^ tickers_x3_lfsrReg_91[2] ^ tickers_x3_lfsrReg_91[3] ^
    tickers_x3_lfsrReg_91[5];
  wire [14:0] tickers_x3_lfsrReg_lo_91 = tickers_x3_lfsrReg_91[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_643 = {tickers_x3_lfsrReg_hi_91,tickers_x3_lfsrReg_lo_91};
  reg [15:0] tickers_x3_lfsrReg_92;
  wire  tickers_x3_lfsrReg_hi_92 = tickers_x3_lfsrReg_92[0] ^ tickers_x3_lfsrReg_92[2] ^ tickers_x3_lfsrReg_92[3] ^
    tickers_x3_lfsrReg_92[5];
  wire [14:0] tickers_x3_lfsrReg_lo_92 = tickers_x3_lfsrReg_92[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_650 = {tickers_x3_lfsrReg_hi_92,tickers_x3_lfsrReg_lo_92};
  reg [15:0] tickers_x3_lfsrReg_93;
  wire  tickers_x3_lfsrReg_hi_93 = tickers_x3_lfsrReg_93[0] ^ tickers_x3_lfsrReg_93[2] ^ tickers_x3_lfsrReg_93[3] ^
    tickers_x3_lfsrReg_93[5];
  wire [14:0] tickers_x3_lfsrReg_lo_93 = tickers_x3_lfsrReg_93[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_657 = {tickers_x3_lfsrReg_hi_93,tickers_x3_lfsrReg_lo_93};
  reg [15:0] tickers_x3_lfsrReg_94;
  wire  tickers_x3_lfsrReg_hi_94 = tickers_x3_lfsrReg_94[0] ^ tickers_x3_lfsrReg_94[2] ^ tickers_x3_lfsrReg_94[3] ^
    tickers_x3_lfsrReg_94[5];
  wire [14:0] tickers_x3_lfsrReg_lo_94 = tickers_x3_lfsrReg_94[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_664 = {tickers_x3_lfsrReg_hi_94,tickers_x3_lfsrReg_lo_94};
  reg [15:0] tickers_x3_lfsrReg_95;
  wire  tickers_x3_lfsrReg_hi_95 = tickers_x3_lfsrReg_95[0] ^ tickers_x3_lfsrReg_95[2] ^ tickers_x3_lfsrReg_95[3] ^
    tickers_x3_lfsrReg_95[5];
  wire [14:0] tickers_x3_lfsrReg_lo_95 = tickers_x3_lfsrReg_95[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_671 = {tickers_x3_lfsrReg_hi_95,tickers_x3_lfsrReg_lo_95};
  reg [15:0] tickers_x3_lfsrReg_96;
  wire  tickers_x3_lfsrReg_hi_96 = tickers_x3_lfsrReg_96[0] ^ tickers_x3_lfsrReg_96[2] ^ tickers_x3_lfsrReg_96[3] ^
    tickers_x3_lfsrReg_96[5];
  wire [14:0] tickers_x3_lfsrReg_lo_96 = tickers_x3_lfsrReg_96[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_678 = {tickers_x3_lfsrReg_hi_96,tickers_x3_lfsrReg_lo_96};
  reg [15:0] tickers_x3_lfsrReg_97;
  wire  tickers_x3_lfsrReg_hi_97 = tickers_x3_lfsrReg_97[0] ^ tickers_x3_lfsrReg_97[2] ^ tickers_x3_lfsrReg_97[3] ^
    tickers_x3_lfsrReg_97[5];
  wire [14:0] tickers_x3_lfsrReg_lo_97 = tickers_x3_lfsrReg_97[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_685 = {tickers_x3_lfsrReg_hi_97,tickers_x3_lfsrReg_lo_97};
  reg [15:0] tickers_x3_lfsrReg_98;
  wire  tickers_x3_lfsrReg_hi_98 = tickers_x3_lfsrReg_98[0] ^ tickers_x3_lfsrReg_98[2] ^ tickers_x3_lfsrReg_98[3] ^
    tickers_x3_lfsrReg_98[5];
  wire [14:0] tickers_x3_lfsrReg_lo_98 = tickers_x3_lfsrReg_98[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_692 = {tickers_x3_lfsrReg_hi_98,tickers_x3_lfsrReg_lo_98};
  reg [15:0] tickers_x3_lfsrReg_99;
  wire  tickers_x3_lfsrReg_hi_99 = tickers_x3_lfsrReg_99[0] ^ tickers_x3_lfsrReg_99[2] ^ tickers_x3_lfsrReg_99[3] ^
    tickers_x3_lfsrReg_99[5];
  wire [14:0] tickers_x3_lfsrReg_lo_99 = tickers_x3_lfsrReg_99[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_699 = {tickers_x3_lfsrReg_hi_99,tickers_x3_lfsrReg_lo_99};
  reg [15:0] tickers_x3_lfsrReg_100;
  wire  tickers_x3_lfsrReg_hi_100 = tickers_x3_lfsrReg_100[0] ^ tickers_x3_lfsrReg_100[2] ^ tickers_x3_lfsrReg_100[3] ^
    tickers_x3_lfsrReg_100[5];
  wire [14:0] tickers_x3_lfsrReg_lo_100 = tickers_x3_lfsrReg_100[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_706 = {tickers_x3_lfsrReg_hi_100,tickers_x3_lfsrReg_lo_100};
  reg [15:0] tickers_x3_lfsrReg_101;
  wire  tickers_x3_lfsrReg_hi_101 = tickers_x3_lfsrReg_101[0] ^ tickers_x3_lfsrReg_101[2] ^ tickers_x3_lfsrReg_101[3] ^
    tickers_x3_lfsrReg_101[5];
  wire [14:0] tickers_x3_lfsrReg_lo_101 = tickers_x3_lfsrReg_101[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_713 = {tickers_x3_lfsrReg_hi_101,tickers_x3_lfsrReg_lo_101};
  reg [15:0] tickers_x3_lfsrReg_102;
  wire  tickers_x3_lfsrReg_hi_102 = tickers_x3_lfsrReg_102[0] ^ tickers_x3_lfsrReg_102[2] ^ tickers_x3_lfsrReg_102[3] ^
    tickers_x3_lfsrReg_102[5];
  wire [14:0] tickers_x3_lfsrReg_lo_102 = tickers_x3_lfsrReg_102[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_720 = {tickers_x3_lfsrReg_hi_102,tickers_x3_lfsrReg_lo_102};
  reg [15:0] tickers_x3_lfsrReg_103;
  wire  tickers_x3_lfsrReg_hi_103 = tickers_x3_lfsrReg_103[0] ^ tickers_x3_lfsrReg_103[2] ^ tickers_x3_lfsrReg_103[3] ^
    tickers_x3_lfsrReg_103[5];
  wire [14:0] tickers_x3_lfsrReg_lo_103 = tickers_x3_lfsrReg_103[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_727 = {tickers_x3_lfsrReg_hi_103,tickers_x3_lfsrReg_lo_103};
  reg [15:0] tickers_x3_lfsrReg_104;
  wire  tickers_x3_lfsrReg_hi_104 = tickers_x3_lfsrReg_104[0] ^ tickers_x3_lfsrReg_104[2] ^ tickers_x3_lfsrReg_104[3] ^
    tickers_x3_lfsrReg_104[5];
  wire [14:0] tickers_x3_lfsrReg_lo_104 = tickers_x3_lfsrReg_104[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_734 = {tickers_x3_lfsrReg_hi_104,tickers_x3_lfsrReg_lo_104};
  reg [15:0] tickers_x3_lfsrReg_105;
  wire  tickers_x3_lfsrReg_hi_105 = tickers_x3_lfsrReg_105[0] ^ tickers_x3_lfsrReg_105[2] ^ tickers_x3_lfsrReg_105[3] ^
    tickers_x3_lfsrReg_105[5];
  wire [14:0] tickers_x3_lfsrReg_lo_105 = tickers_x3_lfsrReg_105[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_741 = {tickers_x3_lfsrReg_hi_105,tickers_x3_lfsrReg_lo_105};
  reg [15:0] tickers_x3_lfsrReg_106;
  wire  tickers_x3_lfsrReg_hi_106 = tickers_x3_lfsrReg_106[0] ^ tickers_x3_lfsrReg_106[2] ^ tickers_x3_lfsrReg_106[3] ^
    tickers_x3_lfsrReg_106[5];
  wire [14:0] tickers_x3_lfsrReg_lo_106 = tickers_x3_lfsrReg_106[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_748 = {tickers_x3_lfsrReg_hi_106,tickers_x3_lfsrReg_lo_106};
  reg [15:0] tickers_x3_lfsrReg_107;
  wire  tickers_x3_lfsrReg_hi_107 = tickers_x3_lfsrReg_107[0] ^ tickers_x3_lfsrReg_107[2] ^ tickers_x3_lfsrReg_107[3] ^
    tickers_x3_lfsrReg_107[5];
  wire [14:0] tickers_x3_lfsrReg_lo_107 = tickers_x3_lfsrReg_107[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_755 = {tickers_x3_lfsrReg_hi_107,tickers_x3_lfsrReg_lo_107};
  reg [15:0] tickers_x3_lfsrReg_108;
  wire  tickers_x3_lfsrReg_hi_108 = tickers_x3_lfsrReg_108[0] ^ tickers_x3_lfsrReg_108[2] ^ tickers_x3_lfsrReg_108[3] ^
    tickers_x3_lfsrReg_108[5];
  wire [14:0] tickers_x3_lfsrReg_lo_108 = tickers_x3_lfsrReg_108[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_762 = {tickers_x3_lfsrReg_hi_108,tickers_x3_lfsrReg_lo_108};
  reg [15:0] tickers_x3_lfsrReg_109;
  wire  tickers_x3_lfsrReg_hi_109 = tickers_x3_lfsrReg_109[0] ^ tickers_x3_lfsrReg_109[2] ^ tickers_x3_lfsrReg_109[3] ^
    tickers_x3_lfsrReg_109[5];
  wire [14:0] tickers_x3_lfsrReg_lo_109 = tickers_x3_lfsrReg_109[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_769 = {tickers_x3_lfsrReg_hi_109,tickers_x3_lfsrReg_lo_109};
  reg [15:0] tickers_x3_lfsrReg_110;
  wire  tickers_x3_lfsrReg_hi_110 = tickers_x3_lfsrReg_110[0] ^ tickers_x3_lfsrReg_110[2] ^ tickers_x3_lfsrReg_110[3] ^
    tickers_x3_lfsrReg_110[5];
  wire [14:0] tickers_x3_lfsrReg_lo_110 = tickers_x3_lfsrReg_110[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_776 = {tickers_x3_lfsrReg_hi_110,tickers_x3_lfsrReg_lo_110};
  reg [15:0] tickers_x3_lfsrReg_111;
  wire  tickers_x3_lfsrReg_hi_111 = tickers_x3_lfsrReg_111[0] ^ tickers_x3_lfsrReg_111[2] ^ tickers_x3_lfsrReg_111[3] ^
    tickers_x3_lfsrReg_111[5];
  wire [14:0] tickers_x3_lfsrReg_lo_111 = tickers_x3_lfsrReg_111[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_783 = {tickers_x3_lfsrReg_hi_111,tickers_x3_lfsrReg_lo_111};
  reg [15:0] tickers_x3_lfsrReg_112;
  wire  tickers_x3_lfsrReg_hi_112 = tickers_x3_lfsrReg_112[0] ^ tickers_x3_lfsrReg_112[2] ^ tickers_x3_lfsrReg_112[3] ^
    tickers_x3_lfsrReg_112[5];
  wire [14:0] tickers_x3_lfsrReg_lo_112 = tickers_x3_lfsrReg_112[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_790 = {tickers_x3_lfsrReg_hi_112,tickers_x3_lfsrReg_lo_112};
  reg [15:0] tickers_x3_lfsrReg_113;
  wire  tickers_x3_lfsrReg_hi_113 = tickers_x3_lfsrReg_113[0] ^ tickers_x3_lfsrReg_113[2] ^ tickers_x3_lfsrReg_113[3] ^
    tickers_x3_lfsrReg_113[5];
  wire [14:0] tickers_x3_lfsrReg_lo_113 = tickers_x3_lfsrReg_113[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_797 = {tickers_x3_lfsrReg_hi_113,tickers_x3_lfsrReg_lo_113};
  reg [15:0] tickers_x3_lfsrReg_114;
  wire  tickers_x3_lfsrReg_hi_114 = tickers_x3_lfsrReg_114[0] ^ tickers_x3_lfsrReg_114[2] ^ tickers_x3_lfsrReg_114[3] ^
    tickers_x3_lfsrReg_114[5];
  wire [14:0] tickers_x3_lfsrReg_lo_114 = tickers_x3_lfsrReg_114[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_804 = {tickers_x3_lfsrReg_hi_114,tickers_x3_lfsrReg_lo_114};
  reg [15:0] tickers_x3_lfsrReg_115;
  wire  tickers_x3_lfsrReg_hi_115 = tickers_x3_lfsrReg_115[0] ^ tickers_x3_lfsrReg_115[2] ^ tickers_x3_lfsrReg_115[3] ^
    tickers_x3_lfsrReg_115[5];
  wire [14:0] tickers_x3_lfsrReg_lo_115 = tickers_x3_lfsrReg_115[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_811 = {tickers_x3_lfsrReg_hi_115,tickers_x3_lfsrReg_lo_115};
  reg [15:0] tickers_x3_lfsrReg_116;
  wire  tickers_x3_lfsrReg_hi_116 = tickers_x3_lfsrReg_116[0] ^ tickers_x3_lfsrReg_116[2] ^ tickers_x3_lfsrReg_116[3] ^
    tickers_x3_lfsrReg_116[5];
  wire [14:0] tickers_x3_lfsrReg_lo_116 = tickers_x3_lfsrReg_116[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_818 = {tickers_x3_lfsrReg_hi_116,tickers_x3_lfsrReg_lo_116};
  reg [15:0] tickers_x3_lfsrReg_117;
  wire  tickers_x3_lfsrReg_hi_117 = tickers_x3_lfsrReg_117[0] ^ tickers_x3_lfsrReg_117[2] ^ tickers_x3_lfsrReg_117[3] ^
    tickers_x3_lfsrReg_117[5];
  wire [14:0] tickers_x3_lfsrReg_lo_117 = tickers_x3_lfsrReg_117[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_825 = {tickers_x3_lfsrReg_hi_117,tickers_x3_lfsrReg_lo_117};
  reg [15:0] tickers_x3_lfsrReg_118;
  wire  tickers_x3_lfsrReg_hi_118 = tickers_x3_lfsrReg_118[0] ^ tickers_x3_lfsrReg_118[2] ^ tickers_x3_lfsrReg_118[3] ^
    tickers_x3_lfsrReg_118[5];
  wire [14:0] tickers_x3_lfsrReg_lo_118 = tickers_x3_lfsrReg_118[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_832 = {tickers_x3_lfsrReg_hi_118,tickers_x3_lfsrReg_lo_118};
  reg [15:0] tickers_x3_lfsrReg_119;
  wire  tickers_x3_lfsrReg_hi_119 = tickers_x3_lfsrReg_119[0] ^ tickers_x3_lfsrReg_119[2] ^ tickers_x3_lfsrReg_119[3] ^
    tickers_x3_lfsrReg_119[5];
  wire [14:0] tickers_x3_lfsrReg_lo_119 = tickers_x3_lfsrReg_119[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_839 = {tickers_x3_lfsrReg_hi_119,tickers_x3_lfsrReg_lo_119};
  reg [15:0] tickers_x3_lfsrReg_120;
  wire  tickers_x3_lfsrReg_hi_120 = tickers_x3_lfsrReg_120[0] ^ tickers_x3_lfsrReg_120[2] ^ tickers_x3_lfsrReg_120[3] ^
    tickers_x3_lfsrReg_120[5];
  wire [14:0] tickers_x3_lfsrReg_lo_120 = tickers_x3_lfsrReg_120[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_846 = {tickers_x3_lfsrReg_hi_120,tickers_x3_lfsrReg_lo_120};
  reg [15:0] tickers_x3_lfsrReg_121;
  wire  tickers_x3_lfsrReg_hi_121 = tickers_x3_lfsrReg_121[0] ^ tickers_x3_lfsrReg_121[2] ^ tickers_x3_lfsrReg_121[3] ^
    tickers_x3_lfsrReg_121[5];
  wire [14:0] tickers_x3_lfsrReg_lo_121 = tickers_x3_lfsrReg_121[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_853 = {tickers_x3_lfsrReg_hi_121,tickers_x3_lfsrReg_lo_121};
  reg [15:0] tickers_x3_lfsrReg_122;
  wire  tickers_x3_lfsrReg_hi_122 = tickers_x3_lfsrReg_122[0] ^ tickers_x3_lfsrReg_122[2] ^ tickers_x3_lfsrReg_122[3] ^
    tickers_x3_lfsrReg_122[5];
  wire [14:0] tickers_x3_lfsrReg_lo_122 = tickers_x3_lfsrReg_122[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_860 = {tickers_x3_lfsrReg_hi_122,tickers_x3_lfsrReg_lo_122};
  reg [15:0] tickers_x3_lfsrReg_123;
  wire  tickers_x3_lfsrReg_hi_123 = tickers_x3_lfsrReg_123[0] ^ tickers_x3_lfsrReg_123[2] ^ tickers_x3_lfsrReg_123[3] ^
    tickers_x3_lfsrReg_123[5];
  wire [14:0] tickers_x3_lfsrReg_lo_123 = tickers_x3_lfsrReg_123[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_867 = {tickers_x3_lfsrReg_hi_123,tickers_x3_lfsrReg_lo_123};
  reg [15:0] tickers_x3_lfsrReg_124;
  wire  tickers_x3_lfsrReg_hi_124 = tickers_x3_lfsrReg_124[0] ^ tickers_x3_lfsrReg_124[2] ^ tickers_x3_lfsrReg_124[3] ^
    tickers_x3_lfsrReg_124[5];
  wire [14:0] tickers_x3_lfsrReg_lo_124 = tickers_x3_lfsrReg_124[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_874 = {tickers_x3_lfsrReg_hi_124,tickers_x3_lfsrReg_lo_124};
  reg [15:0] tickers_x3_lfsrReg_125;
  wire  tickers_x3_lfsrReg_hi_125 = tickers_x3_lfsrReg_125[0] ^ tickers_x3_lfsrReg_125[2] ^ tickers_x3_lfsrReg_125[3] ^
    tickers_x3_lfsrReg_125[5];
  wire [14:0] tickers_x3_lfsrReg_lo_125 = tickers_x3_lfsrReg_125[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_881 = {tickers_x3_lfsrReg_hi_125,tickers_x3_lfsrReg_lo_125};
  reg [15:0] tickers_x3_lfsrReg_126;
  wire  tickers_x3_lfsrReg_hi_126 = tickers_x3_lfsrReg_126[0] ^ tickers_x3_lfsrReg_126[2] ^ tickers_x3_lfsrReg_126[3] ^
    tickers_x3_lfsrReg_126[5];
  wire [14:0] tickers_x3_lfsrReg_lo_126 = tickers_x3_lfsrReg_126[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_888 = {tickers_x3_lfsrReg_hi_126,tickers_x3_lfsrReg_lo_126};
  reg [15:0] system_global_interrupts_x5_lfsrReg;
  wire  system_global_interrupts_x5_lfsrReg_hi = system_global_interrupts_x5_lfsrReg[0] ^
    system_global_interrupts_x5_lfsrReg[2] ^ system_global_interrupts_x5_lfsrReg[3] ^
    system_global_interrupts_x5_lfsrReg[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo = system_global_interrupts_x5_lfsrReg[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_6 = {system_global_interrupts_x5_lfsrReg_hi,
    system_global_interrupts_x5_lfsrReg_lo};
  reg [15:0] system_global_interrupts_x5_lfsrReg_1;
  wire  system_global_interrupts_x5_lfsrReg_hi_1 = system_global_interrupts_x5_lfsrReg_1[0] ^
    system_global_interrupts_x5_lfsrReg_1[2] ^ system_global_interrupts_x5_lfsrReg_1[3] ^
    system_global_interrupts_x5_lfsrReg_1[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_1 = system_global_interrupts_x5_lfsrReg_1[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_13 = {system_global_interrupts_x5_lfsrReg_hi_1,
    system_global_interrupts_x5_lfsrReg_lo_1};
  reg [15:0] system_global_interrupts_x5_lfsrReg_2;
  wire  system_global_interrupts_x5_lfsrReg_hi_2 = system_global_interrupts_x5_lfsrReg_2[0] ^
    system_global_interrupts_x5_lfsrReg_2[2] ^ system_global_interrupts_x5_lfsrReg_2[3] ^
    system_global_interrupts_x5_lfsrReg_2[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_2 = system_global_interrupts_x5_lfsrReg_2[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_20 = {system_global_interrupts_x5_lfsrReg_hi_2,
    system_global_interrupts_x5_lfsrReg_lo_2};
  reg [15:0] system_global_interrupts_x5_lfsrReg_3;
  wire  system_global_interrupts_x5_lfsrReg_hi_3 = system_global_interrupts_x5_lfsrReg_3[0] ^
    system_global_interrupts_x5_lfsrReg_3[2] ^ system_global_interrupts_x5_lfsrReg_3[3] ^
    system_global_interrupts_x5_lfsrReg_3[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_3 = system_global_interrupts_x5_lfsrReg_3[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_27 = {system_global_interrupts_x5_lfsrReg_hi_3,
    system_global_interrupts_x5_lfsrReg_lo_3};
  reg [15:0] system_global_interrupts_x5_lfsrReg_4;
  wire  system_global_interrupts_x5_lfsrReg_hi_4 = system_global_interrupts_x5_lfsrReg_4[0] ^
    system_global_interrupts_x5_lfsrReg_4[2] ^ system_global_interrupts_x5_lfsrReg_4[3] ^
    system_global_interrupts_x5_lfsrReg_4[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_4 = system_global_interrupts_x5_lfsrReg_4[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_34 = {system_global_interrupts_x5_lfsrReg_hi_4,
    system_global_interrupts_x5_lfsrReg_lo_4};
  reg [15:0] system_global_interrupts_x5_lfsrReg_5;
  wire  system_global_interrupts_x5_lfsrReg_hi_5 = system_global_interrupts_x5_lfsrReg_5[0] ^
    system_global_interrupts_x5_lfsrReg_5[2] ^ system_global_interrupts_x5_lfsrReg_5[3] ^
    system_global_interrupts_x5_lfsrReg_5[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_5 = system_global_interrupts_x5_lfsrReg_5[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_41 = {system_global_interrupts_x5_lfsrReg_hi_5,
    system_global_interrupts_x5_lfsrReg_lo_5};
  reg [15:0] system_global_interrupts_x5_lfsrReg_6;
  wire  system_global_interrupts_x5_lfsrReg_hi_6 = system_global_interrupts_x5_lfsrReg_6[0] ^
    system_global_interrupts_x5_lfsrReg_6[2] ^ system_global_interrupts_x5_lfsrReg_6[3] ^
    system_global_interrupts_x5_lfsrReg_6[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_6 = system_global_interrupts_x5_lfsrReg_6[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_48 = {system_global_interrupts_x5_lfsrReg_hi_6,
    system_global_interrupts_x5_lfsrReg_lo_6};
  reg [15:0] system_global_interrupts_x5_lfsrReg_7;
  wire  system_global_interrupts_x5_lfsrReg_hi_7 = system_global_interrupts_x5_lfsrReg_7[0] ^
    system_global_interrupts_x5_lfsrReg_7[2] ^ system_global_interrupts_x5_lfsrReg_7[3] ^
    system_global_interrupts_x5_lfsrReg_7[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_7 = system_global_interrupts_x5_lfsrReg_7[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_55 = {system_global_interrupts_x5_lfsrReg_hi_7,
    system_global_interrupts_x5_lfsrReg_lo_7};
  reg [15:0] system_global_interrupts_x5_lfsrReg_8;
  wire  system_global_interrupts_x5_lfsrReg_hi_8 = system_global_interrupts_x5_lfsrReg_8[0] ^
    system_global_interrupts_x5_lfsrReg_8[2] ^ system_global_interrupts_x5_lfsrReg_8[3] ^
    system_global_interrupts_x5_lfsrReg_8[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_8 = system_global_interrupts_x5_lfsrReg_8[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_62 = {system_global_interrupts_x5_lfsrReg_hi_8,
    system_global_interrupts_x5_lfsrReg_lo_8};
  reg [15:0] system_global_interrupts_x5_lfsrReg_9;
  wire  system_global_interrupts_x5_lfsrReg_hi_9 = system_global_interrupts_x5_lfsrReg_9[0] ^
    system_global_interrupts_x5_lfsrReg_9[2] ^ system_global_interrupts_x5_lfsrReg_9[3] ^
    system_global_interrupts_x5_lfsrReg_9[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_9 = system_global_interrupts_x5_lfsrReg_9[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_69 = {system_global_interrupts_x5_lfsrReg_hi_9,
    system_global_interrupts_x5_lfsrReg_lo_9};
  reg [15:0] system_global_interrupts_x5_lfsrReg_10;
  wire  system_global_interrupts_x5_lfsrReg_hi_10 = system_global_interrupts_x5_lfsrReg_10[0] ^
    system_global_interrupts_x5_lfsrReg_10[2] ^ system_global_interrupts_x5_lfsrReg_10[3] ^
    system_global_interrupts_x5_lfsrReg_10[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_10 = system_global_interrupts_x5_lfsrReg_10[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_76 = {system_global_interrupts_x5_lfsrReg_hi_10,
    system_global_interrupts_x5_lfsrReg_lo_10};
  reg [15:0] system_global_interrupts_x5_lfsrReg_11;
  wire  system_global_interrupts_x5_lfsrReg_hi_11 = system_global_interrupts_x5_lfsrReg_11[0] ^
    system_global_interrupts_x5_lfsrReg_11[2] ^ system_global_interrupts_x5_lfsrReg_11[3] ^
    system_global_interrupts_x5_lfsrReg_11[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_11 = system_global_interrupts_x5_lfsrReg_11[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_83 = {system_global_interrupts_x5_lfsrReg_hi_11,
    system_global_interrupts_x5_lfsrReg_lo_11};
  reg [15:0] system_global_interrupts_x5_lfsrReg_12;
  wire  system_global_interrupts_x5_lfsrReg_hi_12 = system_global_interrupts_x5_lfsrReg_12[0] ^
    system_global_interrupts_x5_lfsrReg_12[2] ^ system_global_interrupts_x5_lfsrReg_12[3] ^
    system_global_interrupts_x5_lfsrReg_12[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_12 = system_global_interrupts_x5_lfsrReg_12[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_90 = {system_global_interrupts_x5_lfsrReg_hi_12,
    system_global_interrupts_x5_lfsrReg_lo_12};
  reg [15:0] system_global_interrupts_x5_lfsrReg_13;
  wire  system_global_interrupts_x5_lfsrReg_hi_13 = system_global_interrupts_x5_lfsrReg_13[0] ^
    system_global_interrupts_x5_lfsrReg_13[2] ^ system_global_interrupts_x5_lfsrReg_13[3] ^
    system_global_interrupts_x5_lfsrReg_13[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_13 = system_global_interrupts_x5_lfsrReg_13[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_97 = {system_global_interrupts_x5_lfsrReg_hi_13,
    system_global_interrupts_x5_lfsrReg_lo_13};
  reg [15:0] system_global_interrupts_x5_lfsrReg_14;
  wire  system_global_interrupts_x5_lfsrReg_hi_14 = system_global_interrupts_x5_lfsrReg_14[0] ^
    system_global_interrupts_x5_lfsrReg_14[2] ^ system_global_interrupts_x5_lfsrReg_14[3] ^
    system_global_interrupts_x5_lfsrReg_14[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_14 = system_global_interrupts_x5_lfsrReg_14[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_104 = {system_global_interrupts_x5_lfsrReg_hi_14,
    system_global_interrupts_x5_lfsrReg_lo_14};
  reg [15:0] system_global_interrupts_x5_lfsrReg_15;
  wire  system_global_interrupts_x5_lfsrReg_hi_15 = system_global_interrupts_x5_lfsrReg_15[0] ^
    system_global_interrupts_x5_lfsrReg_15[2] ^ system_global_interrupts_x5_lfsrReg_15[3] ^
    system_global_interrupts_x5_lfsrReg_15[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_15 = system_global_interrupts_x5_lfsrReg_15[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_111 = {system_global_interrupts_x5_lfsrReg_hi_15,
    system_global_interrupts_x5_lfsrReg_lo_15};
  reg [15:0] system_global_interrupts_x5_lfsrReg_16;
  wire  system_global_interrupts_x5_lfsrReg_hi_16 = system_global_interrupts_x5_lfsrReg_16[0] ^
    system_global_interrupts_x5_lfsrReg_16[2] ^ system_global_interrupts_x5_lfsrReg_16[3] ^
    system_global_interrupts_x5_lfsrReg_16[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_16 = system_global_interrupts_x5_lfsrReg_16[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_118 = {system_global_interrupts_x5_lfsrReg_hi_16,
    system_global_interrupts_x5_lfsrReg_lo_16};
  reg [15:0] system_global_interrupts_x5_lfsrReg_17;
  wire  system_global_interrupts_x5_lfsrReg_hi_17 = system_global_interrupts_x5_lfsrReg_17[0] ^
    system_global_interrupts_x5_lfsrReg_17[2] ^ system_global_interrupts_x5_lfsrReg_17[3] ^
    system_global_interrupts_x5_lfsrReg_17[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_17 = system_global_interrupts_x5_lfsrReg_17[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_125 = {system_global_interrupts_x5_lfsrReg_hi_17,
    system_global_interrupts_x5_lfsrReg_lo_17};
  reg [15:0] system_global_interrupts_x5_lfsrReg_18;
  wire  system_global_interrupts_x5_lfsrReg_hi_18 = system_global_interrupts_x5_lfsrReg_18[0] ^
    system_global_interrupts_x5_lfsrReg_18[2] ^ system_global_interrupts_x5_lfsrReg_18[3] ^
    system_global_interrupts_x5_lfsrReg_18[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_18 = system_global_interrupts_x5_lfsrReg_18[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_132 = {system_global_interrupts_x5_lfsrReg_hi_18,
    system_global_interrupts_x5_lfsrReg_lo_18};
  reg [15:0] system_global_interrupts_x5_lfsrReg_19;
  wire  system_global_interrupts_x5_lfsrReg_hi_19 = system_global_interrupts_x5_lfsrReg_19[0] ^
    system_global_interrupts_x5_lfsrReg_19[2] ^ system_global_interrupts_x5_lfsrReg_19[3] ^
    system_global_interrupts_x5_lfsrReg_19[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_19 = system_global_interrupts_x5_lfsrReg_19[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_139 = {system_global_interrupts_x5_lfsrReg_hi_19,
    system_global_interrupts_x5_lfsrReg_lo_19};
  reg [15:0] system_global_interrupts_x5_lfsrReg_20;
  wire  system_global_interrupts_x5_lfsrReg_hi_20 = system_global_interrupts_x5_lfsrReg_20[0] ^
    system_global_interrupts_x5_lfsrReg_20[2] ^ system_global_interrupts_x5_lfsrReg_20[3] ^
    system_global_interrupts_x5_lfsrReg_20[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_20 = system_global_interrupts_x5_lfsrReg_20[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_146 = {system_global_interrupts_x5_lfsrReg_hi_20,
    system_global_interrupts_x5_lfsrReg_lo_20};
  reg [15:0] system_global_interrupts_x5_lfsrReg_21;
  wire  system_global_interrupts_x5_lfsrReg_hi_21 = system_global_interrupts_x5_lfsrReg_21[0] ^
    system_global_interrupts_x5_lfsrReg_21[2] ^ system_global_interrupts_x5_lfsrReg_21[3] ^
    system_global_interrupts_x5_lfsrReg_21[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_21 = system_global_interrupts_x5_lfsrReg_21[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_153 = {system_global_interrupts_x5_lfsrReg_hi_21,
    system_global_interrupts_x5_lfsrReg_lo_21};
  reg [15:0] system_global_interrupts_x5_lfsrReg_22;
  wire  system_global_interrupts_x5_lfsrReg_hi_22 = system_global_interrupts_x5_lfsrReg_22[0] ^
    system_global_interrupts_x5_lfsrReg_22[2] ^ system_global_interrupts_x5_lfsrReg_22[3] ^
    system_global_interrupts_x5_lfsrReg_22[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_22 = system_global_interrupts_x5_lfsrReg_22[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_160 = {system_global_interrupts_x5_lfsrReg_hi_22,
    system_global_interrupts_x5_lfsrReg_lo_22};
  reg [15:0] system_global_interrupts_x5_lfsrReg_23;
  wire  system_global_interrupts_x5_lfsrReg_hi_23 = system_global_interrupts_x5_lfsrReg_23[0] ^
    system_global_interrupts_x5_lfsrReg_23[2] ^ system_global_interrupts_x5_lfsrReg_23[3] ^
    system_global_interrupts_x5_lfsrReg_23[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_23 = system_global_interrupts_x5_lfsrReg_23[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_167 = {system_global_interrupts_x5_lfsrReg_hi_23,
    system_global_interrupts_x5_lfsrReg_lo_23};
  reg [15:0] system_global_interrupts_x5_lfsrReg_24;
  wire  system_global_interrupts_x5_lfsrReg_hi_24 = system_global_interrupts_x5_lfsrReg_24[0] ^
    system_global_interrupts_x5_lfsrReg_24[2] ^ system_global_interrupts_x5_lfsrReg_24[3] ^
    system_global_interrupts_x5_lfsrReg_24[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_24 = system_global_interrupts_x5_lfsrReg_24[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_174 = {system_global_interrupts_x5_lfsrReg_hi_24,
    system_global_interrupts_x5_lfsrReg_lo_24};
  reg [15:0] system_global_interrupts_x5_lfsrReg_25;
  wire  system_global_interrupts_x5_lfsrReg_hi_25 = system_global_interrupts_x5_lfsrReg_25[0] ^
    system_global_interrupts_x5_lfsrReg_25[2] ^ system_global_interrupts_x5_lfsrReg_25[3] ^
    system_global_interrupts_x5_lfsrReg_25[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_25 = system_global_interrupts_x5_lfsrReg_25[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_181 = {system_global_interrupts_x5_lfsrReg_hi_25,
    system_global_interrupts_x5_lfsrReg_lo_25};
  reg [15:0] system_global_interrupts_x5_lfsrReg_26;
  wire  system_global_interrupts_x5_lfsrReg_hi_26 = system_global_interrupts_x5_lfsrReg_26[0] ^
    system_global_interrupts_x5_lfsrReg_26[2] ^ system_global_interrupts_x5_lfsrReg_26[3] ^
    system_global_interrupts_x5_lfsrReg_26[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_26 = system_global_interrupts_x5_lfsrReg_26[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_188 = {system_global_interrupts_x5_lfsrReg_hi_26,
    system_global_interrupts_x5_lfsrReg_lo_26};
  reg [15:0] system_global_interrupts_x5_lfsrReg_27;
  wire  system_global_interrupts_x5_lfsrReg_hi_27 = system_global_interrupts_x5_lfsrReg_27[0] ^
    system_global_interrupts_x5_lfsrReg_27[2] ^ system_global_interrupts_x5_lfsrReg_27[3] ^
    system_global_interrupts_x5_lfsrReg_27[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_27 = system_global_interrupts_x5_lfsrReg_27[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_195 = {system_global_interrupts_x5_lfsrReg_hi_27,
    system_global_interrupts_x5_lfsrReg_lo_27};
  reg [15:0] system_global_interrupts_x5_lfsrReg_28;
  wire  system_global_interrupts_x5_lfsrReg_hi_28 = system_global_interrupts_x5_lfsrReg_28[0] ^
    system_global_interrupts_x5_lfsrReg_28[2] ^ system_global_interrupts_x5_lfsrReg_28[3] ^
    system_global_interrupts_x5_lfsrReg_28[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_28 = system_global_interrupts_x5_lfsrReg_28[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_202 = {system_global_interrupts_x5_lfsrReg_hi_28,
    system_global_interrupts_x5_lfsrReg_lo_28};
  reg [15:0] system_global_interrupts_x5_lfsrReg_29;
  wire  system_global_interrupts_x5_lfsrReg_hi_29 = system_global_interrupts_x5_lfsrReg_29[0] ^
    system_global_interrupts_x5_lfsrReg_29[2] ^ system_global_interrupts_x5_lfsrReg_29[3] ^
    system_global_interrupts_x5_lfsrReg_29[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_29 = system_global_interrupts_x5_lfsrReg_29[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_209 = {system_global_interrupts_x5_lfsrReg_hi_29,
    system_global_interrupts_x5_lfsrReg_lo_29};
  reg [15:0] system_global_interrupts_x5_lfsrReg_30;
  wire  system_global_interrupts_x5_lfsrReg_hi_30 = system_global_interrupts_x5_lfsrReg_30[0] ^
    system_global_interrupts_x5_lfsrReg_30[2] ^ system_global_interrupts_x5_lfsrReg_30[3] ^
    system_global_interrupts_x5_lfsrReg_30[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_30 = system_global_interrupts_x5_lfsrReg_30[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_216 = {system_global_interrupts_x5_lfsrReg_hi_30,
    system_global_interrupts_x5_lfsrReg_lo_30};
  reg [15:0] system_global_interrupts_x5_lfsrReg_31;
  wire  system_global_interrupts_x5_lfsrReg_hi_31 = system_global_interrupts_x5_lfsrReg_31[0] ^
    system_global_interrupts_x5_lfsrReg_31[2] ^ system_global_interrupts_x5_lfsrReg_31[3] ^
    system_global_interrupts_x5_lfsrReg_31[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_31 = system_global_interrupts_x5_lfsrReg_31[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_223 = {system_global_interrupts_x5_lfsrReg_hi_31,
    system_global_interrupts_x5_lfsrReg_lo_31};
  reg [15:0] system_global_interrupts_x5_lfsrReg_32;
  wire  system_global_interrupts_x5_lfsrReg_hi_32 = system_global_interrupts_x5_lfsrReg_32[0] ^
    system_global_interrupts_x5_lfsrReg_32[2] ^ system_global_interrupts_x5_lfsrReg_32[3] ^
    system_global_interrupts_x5_lfsrReg_32[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_32 = system_global_interrupts_x5_lfsrReg_32[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_230 = {system_global_interrupts_x5_lfsrReg_hi_32,
    system_global_interrupts_x5_lfsrReg_lo_32};
  reg [15:0] system_global_interrupts_x5_lfsrReg_33;
  wire  system_global_interrupts_x5_lfsrReg_hi_33 = system_global_interrupts_x5_lfsrReg_33[0] ^
    system_global_interrupts_x5_lfsrReg_33[2] ^ system_global_interrupts_x5_lfsrReg_33[3] ^
    system_global_interrupts_x5_lfsrReg_33[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_33 = system_global_interrupts_x5_lfsrReg_33[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_237 = {system_global_interrupts_x5_lfsrReg_hi_33,
    system_global_interrupts_x5_lfsrReg_lo_33};
  reg [15:0] system_global_interrupts_x5_lfsrReg_34;
  wire  system_global_interrupts_x5_lfsrReg_hi_34 = system_global_interrupts_x5_lfsrReg_34[0] ^
    system_global_interrupts_x5_lfsrReg_34[2] ^ system_global_interrupts_x5_lfsrReg_34[3] ^
    system_global_interrupts_x5_lfsrReg_34[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_34 = system_global_interrupts_x5_lfsrReg_34[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_244 = {system_global_interrupts_x5_lfsrReg_hi_34,
    system_global_interrupts_x5_lfsrReg_lo_34};
  reg [15:0] system_global_interrupts_x5_lfsrReg_35;
  wire  system_global_interrupts_x5_lfsrReg_hi_35 = system_global_interrupts_x5_lfsrReg_35[0] ^
    system_global_interrupts_x5_lfsrReg_35[2] ^ system_global_interrupts_x5_lfsrReg_35[3] ^
    system_global_interrupts_x5_lfsrReg_35[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_35 = system_global_interrupts_x5_lfsrReg_35[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_251 = {system_global_interrupts_x5_lfsrReg_hi_35,
    system_global_interrupts_x5_lfsrReg_lo_35};
  reg [15:0] system_global_interrupts_x5_lfsrReg_36;
  wire  system_global_interrupts_x5_lfsrReg_hi_36 = system_global_interrupts_x5_lfsrReg_36[0] ^
    system_global_interrupts_x5_lfsrReg_36[2] ^ system_global_interrupts_x5_lfsrReg_36[3] ^
    system_global_interrupts_x5_lfsrReg_36[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_36 = system_global_interrupts_x5_lfsrReg_36[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_258 = {system_global_interrupts_x5_lfsrReg_hi_36,
    system_global_interrupts_x5_lfsrReg_lo_36};
  reg [15:0] system_global_interrupts_x5_lfsrReg_37;
  wire  system_global_interrupts_x5_lfsrReg_hi_37 = system_global_interrupts_x5_lfsrReg_37[0] ^
    system_global_interrupts_x5_lfsrReg_37[2] ^ system_global_interrupts_x5_lfsrReg_37[3] ^
    system_global_interrupts_x5_lfsrReg_37[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_37 = system_global_interrupts_x5_lfsrReg_37[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_265 = {system_global_interrupts_x5_lfsrReg_hi_37,
    system_global_interrupts_x5_lfsrReg_lo_37};
  reg [15:0] system_global_interrupts_x5_lfsrReg_38;
  wire  system_global_interrupts_x5_lfsrReg_hi_38 = system_global_interrupts_x5_lfsrReg_38[0] ^
    system_global_interrupts_x5_lfsrReg_38[2] ^ system_global_interrupts_x5_lfsrReg_38[3] ^
    system_global_interrupts_x5_lfsrReg_38[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_38 = system_global_interrupts_x5_lfsrReg_38[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_272 = {system_global_interrupts_x5_lfsrReg_hi_38,
    system_global_interrupts_x5_lfsrReg_lo_38};
  reg [15:0] system_global_interrupts_x5_lfsrReg_39;
  wire  system_global_interrupts_x5_lfsrReg_hi_39 = system_global_interrupts_x5_lfsrReg_39[0] ^
    system_global_interrupts_x5_lfsrReg_39[2] ^ system_global_interrupts_x5_lfsrReg_39[3] ^
    system_global_interrupts_x5_lfsrReg_39[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_39 = system_global_interrupts_x5_lfsrReg_39[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_279 = {system_global_interrupts_x5_lfsrReg_hi_39,
    system_global_interrupts_x5_lfsrReg_lo_39};
  reg [15:0] system_global_interrupts_x5_lfsrReg_40;
  wire  system_global_interrupts_x5_lfsrReg_hi_40 = system_global_interrupts_x5_lfsrReg_40[0] ^
    system_global_interrupts_x5_lfsrReg_40[2] ^ system_global_interrupts_x5_lfsrReg_40[3] ^
    system_global_interrupts_x5_lfsrReg_40[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_40 = system_global_interrupts_x5_lfsrReg_40[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_286 = {system_global_interrupts_x5_lfsrReg_hi_40,
    system_global_interrupts_x5_lfsrReg_lo_40};
  reg [15:0] system_global_interrupts_x5_lfsrReg_41;
  wire  system_global_interrupts_x5_lfsrReg_hi_41 = system_global_interrupts_x5_lfsrReg_41[0] ^
    system_global_interrupts_x5_lfsrReg_41[2] ^ system_global_interrupts_x5_lfsrReg_41[3] ^
    system_global_interrupts_x5_lfsrReg_41[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_41 = system_global_interrupts_x5_lfsrReg_41[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_293 = {system_global_interrupts_x5_lfsrReg_hi_41,
    system_global_interrupts_x5_lfsrReg_lo_41};
  reg [15:0] system_global_interrupts_x5_lfsrReg_42;
  wire  system_global_interrupts_x5_lfsrReg_hi_42 = system_global_interrupts_x5_lfsrReg_42[0] ^
    system_global_interrupts_x5_lfsrReg_42[2] ^ system_global_interrupts_x5_lfsrReg_42[3] ^
    system_global_interrupts_x5_lfsrReg_42[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_42 = system_global_interrupts_x5_lfsrReg_42[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_300 = {system_global_interrupts_x5_lfsrReg_hi_42,
    system_global_interrupts_x5_lfsrReg_lo_42};
  reg [15:0] system_global_interrupts_x5_lfsrReg_43;
  wire  system_global_interrupts_x5_lfsrReg_hi_43 = system_global_interrupts_x5_lfsrReg_43[0] ^
    system_global_interrupts_x5_lfsrReg_43[2] ^ system_global_interrupts_x5_lfsrReg_43[3] ^
    system_global_interrupts_x5_lfsrReg_43[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_43 = system_global_interrupts_x5_lfsrReg_43[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_307 = {system_global_interrupts_x5_lfsrReg_hi_43,
    system_global_interrupts_x5_lfsrReg_lo_43};
  reg [15:0] system_global_interrupts_x5_lfsrReg_44;
  wire  system_global_interrupts_x5_lfsrReg_hi_44 = system_global_interrupts_x5_lfsrReg_44[0] ^
    system_global_interrupts_x5_lfsrReg_44[2] ^ system_global_interrupts_x5_lfsrReg_44[3] ^
    system_global_interrupts_x5_lfsrReg_44[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_44 = system_global_interrupts_x5_lfsrReg_44[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_314 = {system_global_interrupts_x5_lfsrReg_hi_44,
    system_global_interrupts_x5_lfsrReg_lo_44};
  reg [15:0] system_global_interrupts_x5_lfsrReg_45;
  wire  system_global_interrupts_x5_lfsrReg_hi_45 = system_global_interrupts_x5_lfsrReg_45[0] ^
    system_global_interrupts_x5_lfsrReg_45[2] ^ system_global_interrupts_x5_lfsrReg_45[3] ^
    system_global_interrupts_x5_lfsrReg_45[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_45 = system_global_interrupts_x5_lfsrReg_45[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_321 = {system_global_interrupts_x5_lfsrReg_hi_45,
    system_global_interrupts_x5_lfsrReg_lo_45};
  reg [15:0] system_global_interrupts_x5_lfsrReg_46;
  wire  system_global_interrupts_x5_lfsrReg_hi_46 = system_global_interrupts_x5_lfsrReg_46[0] ^
    system_global_interrupts_x5_lfsrReg_46[2] ^ system_global_interrupts_x5_lfsrReg_46[3] ^
    system_global_interrupts_x5_lfsrReg_46[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_46 = system_global_interrupts_x5_lfsrReg_46[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_328 = {system_global_interrupts_x5_lfsrReg_hi_46,
    system_global_interrupts_x5_lfsrReg_lo_46};
  reg [15:0] system_global_interrupts_x5_lfsrReg_47;
  wire  system_global_interrupts_x5_lfsrReg_hi_47 = system_global_interrupts_x5_lfsrReg_47[0] ^
    system_global_interrupts_x5_lfsrReg_47[2] ^ system_global_interrupts_x5_lfsrReg_47[3] ^
    system_global_interrupts_x5_lfsrReg_47[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_47 = system_global_interrupts_x5_lfsrReg_47[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_335 = {system_global_interrupts_x5_lfsrReg_hi_47,
    system_global_interrupts_x5_lfsrReg_lo_47};
  reg [15:0] system_global_interrupts_x5_lfsrReg_48;
  wire  system_global_interrupts_x5_lfsrReg_hi_48 = system_global_interrupts_x5_lfsrReg_48[0] ^
    system_global_interrupts_x5_lfsrReg_48[2] ^ system_global_interrupts_x5_lfsrReg_48[3] ^
    system_global_interrupts_x5_lfsrReg_48[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_48 = system_global_interrupts_x5_lfsrReg_48[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_342 = {system_global_interrupts_x5_lfsrReg_hi_48,
    system_global_interrupts_x5_lfsrReg_lo_48};
  reg [15:0] system_global_interrupts_x5_lfsrReg_49;
  wire  system_global_interrupts_x5_lfsrReg_hi_49 = system_global_interrupts_x5_lfsrReg_49[0] ^
    system_global_interrupts_x5_lfsrReg_49[2] ^ system_global_interrupts_x5_lfsrReg_49[3] ^
    system_global_interrupts_x5_lfsrReg_49[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_49 = system_global_interrupts_x5_lfsrReg_49[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_349 = {system_global_interrupts_x5_lfsrReg_hi_49,
    system_global_interrupts_x5_lfsrReg_lo_49};
  reg [15:0] system_global_interrupts_x5_lfsrReg_50;
  wire  system_global_interrupts_x5_lfsrReg_hi_50 = system_global_interrupts_x5_lfsrReg_50[0] ^
    system_global_interrupts_x5_lfsrReg_50[2] ^ system_global_interrupts_x5_lfsrReg_50[3] ^
    system_global_interrupts_x5_lfsrReg_50[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_50 = system_global_interrupts_x5_lfsrReg_50[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_356 = {system_global_interrupts_x5_lfsrReg_hi_50,
    system_global_interrupts_x5_lfsrReg_lo_50};
  reg [15:0] system_global_interrupts_x5_lfsrReg_51;
  wire  system_global_interrupts_x5_lfsrReg_hi_51 = system_global_interrupts_x5_lfsrReg_51[0] ^
    system_global_interrupts_x5_lfsrReg_51[2] ^ system_global_interrupts_x5_lfsrReg_51[3] ^
    system_global_interrupts_x5_lfsrReg_51[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_51 = system_global_interrupts_x5_lfsrReg_51[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_363 = {system_global_interrupts_x5_lfsrReg_hi_51,
    system_global_interrupts_x5_lfsrReg_lo_51};
  reg [15:0] system_global_interrupts_x5_lfsrReg_52;
  wire  system_global_interrupts_x5_lfsrReg_hi_52 = system_global_interrupts_x5_lfsrReg_52[0] ^
    system_global_interrupts_x5_lfsrReg_52[2] ^ system_global_interrupts_x5_lfsrReg_52[3] ^
    system_global_interrupts_x5_lfsrReg_52[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_52 = system_global_interrupts_x5_lfsrReg_52[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_370 = {system_global_interrupts_x5_lfsrReg_hi_52,
    system_global_interrupts_x5_lfsrReg_lo_52};
  reg [15:0] system_global_interrupts_x5_lfsrReg_53;
  wire  system_global_interrupts_x5_lfsrReg_hi_53 = system_global_interrupts_x5_lfsrReg_53[0] ^
    system_global_interrupts_x5_lfsrReg_53[2] ^ system_global_interrupts_x5_lfsrReg_53[3] ^
    system_global_interrupts_x5_lfsrReg_53[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_53 = system_global_interrupts_x5_lfsrReg_53[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_377 = {system_global_interrupts_x5_lfsrReg_hi_53,
    system_global_interrupts_x5_lfsrReg_lo_53};
  reg [15:0] system_global_interrupts_x5_lfsrReg_54;
  wire  system_global_interrupts_x5_lfsrReg_hi_54 = system_global_interrupts_x5_lfsrReg_54[0] ^
    system_global_interrupts_x5_lfsrReg_54[2] ^ system_global_interrupts_x5_lfsrReg_54[3] ^
    system_global_interrupts_x5_lfsrReg_54[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_54 = system_global_interrupts_x5_lfsrReg_54[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_384 = {system_global_interrupts_x5_lfsrReg_hi_54,
    system_global_interrupts_x5_lfsrReg_lo_54};
  reg [15:0] system_global_interrupts_x5_lfsrReg_55;
  wire  system_global_interrupts_x5_lfsrReg_hi_55 = system_global_interrupts_x5_lfsrReg_55[0] ^
    system_global_interrupts_x5_lfsrReg_55[2] ^ system_global_interrupts_x5_lfsrReg_55[3] ^
    system_global_interrupts_x5_lfsrReg_55[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_55 = system_global_interrupts_x5_lfsrReg_55[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_391 = {system_global_interrupts_x5_lfsrReg_hi_55,
    system_global_interrupts_x5_lfsrReg_lo_55};
  reg [15:0] system_global_interrupts_x5_lfsrReg_56;
  wire  system_global_interrupts_x5_lfsrReg_hi_56 = system_global_interrupts_x5_lfsrReg_56[0] ^
    system_global_interrupts_x5_lfsrReg_56[2] ^ system_global_interrupts_x5_lfsrReg_56[3] ^
    system_global_interrupts_x5_lfsrReg_56[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_56 = system_global_interrupts_x5_lfsrReg_56[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_398 = {system_global_interrupts_x5_lfsrReg_hi_56,
    system_global_interrupts_x5_lfsrReg_lo_56};
  reg [15:0] system_global_interrupts_x5_lfsrReg_57;
  wire  system_global_interrupts_x5_lfsrReg_hi_57 = system_global_interrupts_x5_lfsrReg_57[0] ^
    system_global_interrupts_x5_lfsrReg_57[2] ^ system_global_interrupts_x5_lfsrReg_57[3] ^
    system_global_interrupts_x5_lfsrReg_57[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_57 = system_global_interrupts_x5_lfsrReg_57[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_405 = {system_global_interrupts_x5_lfsrReg_hi_57,
    system_global_interrupts_x5_lfsrReg_lo_57};
  reg [15:0] system_global_interrupts_x5_lfsrReg_58;
  wire  system_global_interrupts_x5_lfsrReg_hi_58 = system_global_interrupts_x5_lfsrReg_58[0] ^
    system_global_interrupts_x5_lfsrReg_58[2] ^ system_global_interrupts_x5_lfsrReg_58[3] ^
    system_global_interrupts_x5_lfsrReg_58[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_58 = system_global_interrupts_x5_lfsrReg_58[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_412 = {system_global_interrupts_x5_lfsrReg_hi_58,
    system_global_interrupts_x5_lfsrReg_lo_58};
  reg [15:0] system_global_interrupts_x5_lfsrReg_59;
  wire  system_global_interrupts_x5_lfsrReg_hi_59 = system_global_interrupts_x5_lfsrReg_59[0] ^
    system_global_interrupts_x5_lfsrReg_59[2] ^ system_global_interrupts_x5_lfsrReg_59[3] ^
    system_global_interrupts_x5_lfsrReg_59[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_59 = system_global_interrupts_x5_lfsrReg_59[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_419 = {system_global_interrupts_x5_lfsrReg_hi_59,
    system_global_interrupts_x5_lfsrReg_lo_59};
  reg [15:0] system_global_interrupts_x5_lfsrReg_60;
  wire  system_global_interrupts_x5_lfsrReg_hi_60 = system_global_interrupts_x5_lfsrReg_60[0] ^
    system_global_interrupts_x5_lfsrReg_60[2] ^ system_global_interrupts_x5_lfsrReg_60[3] ^
    system_global_interrupts_x5_lfsrReg_60[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_60 = system_global_interrupts_x5_lfsrReg_60[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_426 = {system_global_interrupts_x5_lfsrReg_hi_60,
    system_global_interrupts_x5_lfsrReg_lo_60};
  reg [15:0] system_global_interrupts_x5_lfsrReg_61;
  wire  system_global_interrupts_x5_lfsrReg_hi_61 = system_global_interrupts_x5_lfsrReg_61[0] ^
    system_global_interrupts_x5_lfsrReg_61[2] ^ system_global_interrupts_x5_lfsrReg_61[3] ^
    system_global_interrupts_x5_lfsrReg_61[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_61 = system_global_interrupts_x5_lfsrReg_61[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_433 = {system_global_interrupts_x5_lfsrReg_hi_61,
    system_global_interrupts_x5_lfsrReg_lo_61};
  reg [15:0] system_global_interrupts_x5_lfsrReg_62;
  wire  system_global_interrupts_x5_lfsrReg_hi_62 = system_global_interrupts_x5_lfsrReg_62[0] ^
    system_global_interrupts_x5_lfsrReg_62[2] ^ system_global_interrupts_x5_lfsrReg_62[3] ^
    system_global_interrupts_x5_lfsrReg_62[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_62 = system_global_interrupts_x5_lfsrReg_62[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_440 = {system_global_interrupts_x5_lfsrReg_hi_62,
    system_global_interrupts_x5_lfsrReg_lo_62};
  reg [15:0] system_global_interrupts_x5_lfsrReg_63;
  wire  system_global_interrupts_x5_lfsrReg_hi_63 = system_global_interrupts_x5_lfsrReg_63[0] ^
    system_global_interrupts_x5_lfsrReg_63[2] ^ system_global_interrupts_x5_lfsrReg_63[3] ^
    system_global_interrupts_x5_lfsrReg_63[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_63 = system_global_interrupts_x5_lfsrReg_63[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_447 = {system_global_interrupts_x5_lfsrReg_hi_63,
    system_global_interrupts_x5_lfsrReg_lo_63};
  reg [15:0] system_global_interrupts_x5_lfsrReg_64;
  wire  system_global_interrupts_x5_lfsrReg_hi_64 = system_global_interrupts_x5_lfsrReg_64[0] ^
    system_global_interrupts_x5_lfsrReg_64[2] ^ system_global_interrupts_x5_lfsrReg_64[3] ^
    system_global_interrupts_x5_lfsrReg_64[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_64 = system_global_interrupts_x5_lfsrReg_64[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_454 = {system_global_interrupts_x5_lfsrReg_hi_64,
    system_global_interrupts_x5_lfsrReg_lo_64};
  reg [15:0] system_global_interrupts_x5_lfsrReg_65;
  wire  system_global_interrupts_x5_lfsrReg_hi_65 = system_global_interrupts_x5_lfsrReg_65[0] ^
    system_global_interrupts_x5_lfsrReg_65[2] ^ system_global_interrupts_x5_lfsrReg_65[3] ^
    system_global_interrupts_x5_lfsrReg_65[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_65 = system_global_interrupts_x5_lfsrReg_65[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_461 = {system_global_interrupts_x5_lfsrReg_hi_65,
    system_global_interrupts_x5_lfsrReg_lo_65};
  reg [15:0] system_global_interrupts_x5_lfsrReg_66;
  wire  system_global_interrupts_x5_lfsrReg_hi_66 = system_global_interrupts_x5_lfsrReg_66[0] ^
    system_global_interrupts_x5_lfsrReg_66[2] ^ system_global_interrupts_x5_lfsrReg_66[3] ^
    system_global_interrupts_x5_lfsrReg_66[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_66 = system_global_interrupts_x5_lfsrReg_66[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_468 = {system_global_interrupts_x5_lfsrReg_hi_66,
    system_global_interrupts_x5_lfsrReg_lo_66};
  reg [15:0] system_global_interrupts_x5_lfsrReg_67;
  wire  system_global_interrupts_x5_lfsrReg_hi_67 = system_global_interrupts_x5_lfsrReg_67[0] ^
    system_global_interrupts_x5_lfsrReg_67[2] ^ system_global_interrupts_x5_lfsrReg_67[3] ^
    system_global_interrupts_x5_lfsrReg_67[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_67 = system_global_interrupts_x5_lfsrReg_67[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_475 = {system_global_interrupts_x5_lfsrReg_hi_67,
    system_global_interrupts_x5_lfsrReg_lo_67};
  reg [15:0] system_global_interrupts_x5_lfsrReg_68;
  wire  system_global_interrupts_x5_lfsrReg_hi_68 = system_global_interrupts_x5_lfsrReg_68[0] ^
    system_global_interrupts_x5_lfsrReg_68[2] ^ system_global_interrupts_x5_lfsrReg_68[3] ^
    system_global_interrupts_x5_lfsrReg_68[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_68 = system_global_interrupts_x5_lfsrReg_68[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_482 = {system_global_interrupts_x5_lfsrReg_hi_68,
    system_global_interrupts_x5_lfsrReg_lo_68};
  reg [15:0] system_global_interrupts_x5_lfsrReg_69;
  wire  system_global_interrupts_x5_lfsrReg_hi_69 = system_global_interrupts_x5_lfsrReg_69[0] ^
    system_global_interrupts_x5_lfsrReg_69[2] ^ system_global_interrupts_x5_lfsrReg_69[3] ^
    system_global_interrupts_x5_lfsrReg_69[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_69 = system_global_interrupts_x5_lfsrReg_69[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_489 = {system_global_interrupts_x5_lfsrReg_hi_69,
    system_global_interrupts_x5_lfsrReg_lo_69};
  reg [15:0] system_global_interrupts_x5_lfsrReg_70;
  wire  system_global_interrupts_x5_lfsrReg_hi_70 = system_global_interrupts_x5_lfsrReg_70[0] ^
    system_global_interrupts_x5_lfsrReg_70[2] ^ system_global_interrupts_x5_lfsrReg_70[3] ^
    system_global_interrupts_x5_lfsrReg_70[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_70 = system_global_interrupts_x5_lfsrReg_70[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_496 = {system_global_interrupts_x5_lfsrReg_hi_70,
    system_global_interrupts_x5_lfsrReg_lo_70};
  reg [15:0] system_global_interrupts_x5_lfsrReg_71;
  wire  system_global_interrupts_x5_lfsrReg_hi_71 = system_global_interrupts_x5_lfsrReg_71[0] ^
    system_global_interrupts_x5_lfsrReg_71[2] ^ system_global_interrupts_x5_lfsrReg_71[3] ^
    system_global_interrupts_x5_lfsrReg_71[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_71 = system_global_interrupts_x5_lfsrReg_71[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_503 = {system_global_interrupts_x5_lfsrReg_hi_71,
    system_global_interrupts_x5_lfsrReg_lo_71};
  reg [15:0] system_global_interrupts_x5_lfsrReg_72;
  wire  system_global_interrupts_x5_lfsrReg_hi_72 = system_global_interrupts_x5_lfsrReg_72[0] ^
    system_global_interrupts_x5_lfsrReg_72[2] ^ system_global_interrupts_x5_lfsrReg_72[3] ^
    system_global_interrupts_x5_lfsrReg_72[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_72 = system_global_interrupts_x5_lfsrReg_72[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_510 = {system_global_interrupts_x5_lfsrReg_hi_72,
    system_global_interrupts_x5_lfsrReg_lo_72};
  reg [15:0] system_global_interrupts_x5_lfsrReg_73;
  wire  system_global_interrupts_x5_lfsrReg_hi_73 = system_global_interrupts_x5_lfsrReg_73[0] ^
    system_global_interrupts_x5_lfsrReg_73[2] ^ system_global_interrupts_x5_lfsrReg_73[3] ^
    system_global_interrupts_x5_lfsrReg_73[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_73 = system_global_interrupts_x5_lfsrReg_73[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_517 = {system_global_interrupts_x5_lfsrReg_hi_73,
    system_global_interrupts_x5_lfsrReg_lo_73};
  reg [15:0] system_global_interrupts_x5_lfsrReg_74;
  wire  system_global_interrupts_x5_lfsrReg_hi_74 = system_global_interrupts_x5_lfsrReg_74[0] ^
    system_global_interrupts_x5_lfsrReg_74[2] ^ system_global_interrupts_x5_lfsrReg_74[3] ^
    system_global_interrupts_x5_lfsrReg_74[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_74 = system_global_interrupts_x5_lfsrReg_74[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_524 = {system_global_interrupts_x5_lfsrReg_hi_74,
    system_global_interrupts_x5_lfsrReg_lo_74};
  reg [15:0] system_global_interrupts_x5_lfsrReg_75;
  wire  system_global_interrupts_x5_lfsrReg_hi_75 = system_global_interrupts_x5_lfsrReg_75[0] ^
    system_global_interrupts_x5_lfsrReg_75[2] ^ system_global_interrupts_x5_lfsrReg_75[3] ^
    system_global_interrupts_x5_lfsrReg_75[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_75 = system_global_interrupts_x5_lfsrReg_75[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_531 = {system_global_interrupts_x5_lfsrReg_hi_75,
    system_global_interrupts_x5_lfsrReg_lo_75};
  reg [15:0] system_global_interrupts_x5_lfsrReg_76;
  wire  system_global_interrupts_x5_lfsrReg_hi_76 = system_global_interrupts_x5_lfsrReg_76[0] ^
    system_global_interrupts_x5_lfsrReg_76[2] ^ system_global_interrupts_x5_lfsrReg_76[3] ^
    system_global_interrupts_x5_lfsrReg_76[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_76 = system_global_interrupts_x5_lfsrReg_76[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_538 = {system_global_interrupts_x5_lfsrReg_hi_76,
    system_global_interrupts_x5_lfsrReg_lo_76};
  reg [15:0] system_global_interrupts_x5_lfsrReg_77;
  wire  system_global_interrupts_x5_lfsrReg_hi_77 = system_global_interrupts_x5_lfsrReg_77[0] ^
    system_global_interrupts_x5_lfsrReg_77[2] ^ system_global_interrupts_x5_lfsrReg_77[3] ^
    system_global_interrupts_x5_lfsrReg_77[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_77 = system_global_interrupts_x5_lfsrReg_77[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_545 = {system_global_interrupts_x5_lfsrReg_hi_77,
    system_global_interrupts_x5_lfsrReg_lo_77};
  reg [15:0] system_global_interrupts_x5_lfsrReg_78;
  wire  system_global_interrupts_x5_lfsrReg_hi_78 = system_global_interrupts_x5_lfsrReg_78[0] ^
    system_global_interrupts_x5_lfsrReg_78[2] ^ system_global_interrupts_x5_lfsrReg_78[3] ^
    system_global_interrupts_x5_lfsrReg_78[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_78 = system_global_interrupts_x5_lfsrReg_78[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_552 = {system_global_interrupts_x5_lfsrReg_hi_78,
    system_global_interrupts_x5_lfsrReg_lo_78};
  reg [15:0] system_global_interrupts_x5_lfsrReg_79;
  wire  system_global_interrupts_x5_lfsrReg_hi_79 = system_global_interrupts_x5_lfsrReg_79[0] ^
    system_global_interrupts_x5_lfsrReg_79[2] ^ system_global_interrupts_x5_lfsrReg_79[3] ^
    system_global_interrupts_x5_lfsrReg_79[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_79 = system_global_interrupts_x5_lfsrReg_79[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_559 = {system_global_interrupts_x5_lfsrReg_hi_79,
    system_global_interrupts_x5_lfsrReg_lo_79};
  reg [15:0] system_global_interrupts_x5_lfsrReg_80;
  wire  system_global_interrupts_x5_lfsrReg_hi_80 = system_global_interrupts_x5_lfsrReg_80[0] ^
    system_global_interrupts_x5_lfsrReg_80[2] ^ system_global_interrupts_x5_lfsrReg_80[3] ^
    system_global_interrupts_x5_lfsrReg_80[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_80 = system_global_interrupts_x5_lfsrReg_80[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_566 = {system_global_interrupts_x5_lfsrReg_hi_80,
    system_global_interrupts_x5_lfsrReg_lo_80};
  reg [15:0] system_global_interrupts_x5_lfsrReg_81;
  wire  system_global_interrupts_x5_lfsrReg_hi_81 = system_global_interrupts_x5_lfsrReg_81[0] ^
    system_global_interrupts_x5_lfsrReg_81[2] ^ system_global_interrupts_x5_lfsrReg_81[3] ^
    system_global_interrupts_x5_lfsrReg_81[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_81 = system_global_interrupts_x5_lfsrReg_81[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_573 = {system_global_interrupts_x5_lfsrReg_hi_81,
    system_global_interrupts_x5_lfsrReg_lo_81};
  reg [15:0] system_global_interrupts_x5_lfsrReg_82;
  wire  system_global_interrupts_x5_lfsrReg_hi_82 = system_global_interrupts_x5_lfsrReg_82[0] ^
    system_global_interrupts_x5_lfsrReg_82[2] ^ system_global_interrupts_x5_lfsrReg_82[3] ^
    system_global_interrupts_x5_lfsrReg_82[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_82 = system_global_interrupts_x5_lfsrReg_82[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_580 = {system_global_interrupts_x5_lfsrReg_hi_82,
    system_global_interrupts_x5_lfsrReg_lo_82};
  reg [15:0] system_global_interrupts_x5_lfsrReg_83;
  wire  system_global_interrupts_x5_lfsrReg_hi_83 = system_global_interrupts_x5_lfsrReg_83[0] ^
    system_global_interrupts_x5_lfsrReg_83[2] ^ system_global_interrupts_x5_lfsrReg_83[3] ^
    system_global_interrupts_x5_lfsrReg_83[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_83 = system_global_interrupts_x5_lfsrReg_83[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_587 = {system_global_interrupts_x5_lfsrReg_hi_83,
    system_global_interrupts_x5_lfsrReg_lo_83};
  reg [15:0] system_global_interrupts_x5_lfsrReg_84;
  wire  system_global_interrupts_x5_lfsrReg_hi_84 = system_global_interrupts_x5_lfsrReg_84[0] ^
    system_global_interrupts_x5_lfsrReg_84[2] ^ system_global_interrupts_x5_lfsrReg_84[3] ^
    system_global_interrupts_x5_lfsrReg_84[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_84 = system_global_interrupts_x5_lfsrReg_84[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_594 = {system_global_interrupts_x5_lfsrReg_hi_84,
    system_global_interrupts_x5_lfsrReg_lo_84};
  reg [15:0] system_global_interrupts_x5_lfsrReg_85;
  wire  system_global_interrupts_x5_lfsrReg_hi_85 = system_global_interrupts_x5_lfsrReg_85[0] ^
    system_global_interrupts_x5_lfsrReg_85[2] ^ system_global_interrupts_x5_lfsrReg_85[3] ^
    system_global_interrupts_x5_lfsrReg_85[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_85 = system_global_interrupts_x5_lfsrReg_85[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_601 = {system_global_interrupts_x5_lfsrReg_hi_85,
    system_global_interrupts_x5_lfsrReg_lo_85};
  reg [15:0] system_global_interrupts_x5_lfsrReg_86;
  wire  system_global_interrupts_x5_lfsrReg_hi_86 = system_global_interrupts_x5_lfsrReg_86[0] ^
    system_global_interrupts_x5_lfsrReg_86[2] ^ system_global_interrupts_x5_lfsrReg_86[3] ^
    system_global_interrupts_x5_lfsrReg_86[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_86 = system_global_interrupts_x5_lfsrReg_86[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_608 = {system_global_interrupts_x5_lfsrReg_hi_86,
    system_global_interrupts_x5_lfsrReg_lo_86};
  reg [15:0] system_global_interrupts_x5_lfsrReg_87;
  wire  system_global_interrupts_x5_lfsrReg_hi_87 = system_global_interrupts_x5_lfsrReg_87[0] ^
    system_global_interrupts_x5_lfsrReg_87[2] ^ system_global_interrupts_x5_lfsrReg_87[3] ^
    system_global_interrupts_x5_lfsrReg_87[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_87 = system_global_interrupts_x5_lfsrReg_87[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_615 = {system_global_interrupts_x5_lfsrReg_hi_87,
    system_global_interrupts_x5_lfsrReg_lo_87};
  reg [15:0] system_global_interrupts_x5_lfsrReg_88;
  wire  system_global_interrupts_x5_lfsrReg_hi_88 = system_global_interrupts_x5_lfsrReg_88[0] ^
    system_global_interrupts_x5_lfsrReg_88[2] ^ system_global_interrupts_x5_lfsrReg_88[3] ^
    system_global_interrupts_x5_lfsrReg_88[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_88 = system_global_interrupts_x5_lfsrReg_88[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_622 = {system_global_interrupts_x5_lfsrReg_hi_88,
    system_global_interrupts_x5_lfsrReg_lo_88};
  reg [15:0] system_global_interrupts_x5_lfsrReg_89;
  wire  system_global_interrupts_x5_lfsrReg_hi_89 = system_global_interrupts_x5_lfsrReg_89[0] ^
    system_global_interrupts_x5_lfsrReg_89[2] ^ system_global_interrupts_x5_lfsrReg_89[3] ^
    system_global_interrupts_x5_lfsrReg_89[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_89 = system_global_interrupts_x5_lfsrReg_89[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_629 = {system_global_interrupts_x5_lfsrReg_hi_89,
    system_global_interrupts_x5_lfsrReg_lo_89};
  reg [15:0] system_global_interrupts_x5_lfsrReg_90;
  wire  system_global_interrupts_x5_lfsrReg_hi_90 = system_global_interrupts_x5_lfsrReg_90[0] ^
    system_global_interrupts_x5_lfsrReg_90[2] ^ system_global_interrupts_x5_lfsrReg_90[3] ^
    system_global_interrupts_x5_lfsrReg_90[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_90 = system_global_interrupts_x5_lfsrReg_90[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_636 = {system_global_interrupts_x5_lfsrReg_hi_90,
    system_global_interrupts_x5_lfsrReg_lo_90};
  reg [15:0] system_global_interrupts_x5_lfsrReg_91;
  wire  system_global_interrupts_x5_lfsrReg_hi_91 = system_global_interrupts_x5_lfsrReg_91[0] ^
    system_global_interrupts_x5_lfsrReg_91[2] ^ system_global_interrupts_x5_lfsrReg_91[3] ^
    system_global_interrupts_x5_lfsrReg_91[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_91 = system_global_interrupts_x5_lfsrReg_91[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_643 = {system_global_interrupts_x5_lfsrReg_hi_91,
    system_global_interrupts_x5_lfsrReg_lo_91};
  reg [15:0] system_global_interrupts_x5_lfsrReg_92;
  wire  system_global_interrupts_x5_lfsrReg_hi_92 = system_global_interrupts_x5_lfsrReg_92[0] ^
    system_global_interrupts_x5_lfsrReg_92[2] ^ system_global_interrupts_x5_lfsrReg_92[3] ^
    system_global_interrupts_x5_lfsrReg_92[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_92 = system_global_interrupts_x5_lfsrReg_92[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_650 = {system_global_interrupts_x5_lfsrReg_hi_92,
    system_global_interrupts_x5_lfsrReg_lo_92};
  reg [15:0] system_global_interrupts_x5_lfsrReg_93;
  wire  system_global_interrupts_x5_lfsrReg_hi_93 = system_global_interrupts_x5_lfsrReg_93[0] ^
    system_global_interrupts_x5_lfsrReg_93[2] ^ system_global_interrupts_x5_lfsrReg_93[3] ^
    system_global_interrupts_x5_lfsrReg_93[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_93 = system_global_interrupts_x5_lfsrReg_93[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_657 = {system_global_interrupts_x5_lfsrReg_hi_93,
    system_global_interrupts_x5_lfsrReg_lo_93};
  reg [15:0] system_global_interrupts_x5_lfsrReg_94;
  wire  system_global_interrupts_x5_lfsrReg_hi_94 = system_global_interrupts_x5_lfsrReg_94[0] ^
    system_global_interrupts_x5_lfsrReg_94[2] ^ system_global_interrupts_x5_lfsrReg_94[3] ^
    system_global_interrupts_x5_lfsrReg_94[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_94 = system_global_interrupts_x5_lfsrReg_94[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_664 = {system_global_interrupts_x5_lfsrReg_hi_94,
    system_global_interrupts_x5_lfsrReg_lo_94};
  reg [15:0] system_global_interrupts_x5_lfsrReg_95;
  wire  system_global_interrupts_x5_lfsrReg_hi_95 = system_global_interrupts_x5_lfsrReg_95[0] ^
    system_global_interrupts_x5_lfsrReg_95[2] ^ system_global_interrupts_x5_lfsrReg_95[3] ^
    system_global_interrupts_x5_lfsrReg_95[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_95 = system_global_interrupts_x5_lfsrReg_95[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_671 = {system_global_interrupts_x5_lfsrReg_hi_95,
    system_global_interrupts_x5_lfsrReg_lo_95};
  reg [15:0] system_global_interrupts_x5_lfsrReg_96;
  wire  system_global_interrupts_x5_lfsrReg_hi_96 = system_global_interrupts_x5_lfsrReg_96[0] ^
    system_global_interrupts_x5_lfsrReg_96[2] ^ system_global_interrupts_x5_lfsrReg_96[3] ^
    system_global_interrupts_x5_lfsrReg_96[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_96 = system_global_interrupts_x5_lfsrReg_96[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_678 = {system_global_interrupts_x5_lfsrReg_hi_96,
    system_global_interrupts_x5_lfsrReg_lo_96};
  reg [15:0] system_global_interrupts_x5_lfsrReg_97;
  wire  system_global_interrupts_x5_lfsrReg_hi_97 = system_global_interrupts_x5_lfsrReg_97[0] ^
    system_global_interrupts_x5_lfsrReg_97[2] ^ system_global_interrupts_x5_lfsrReg_97[3] ^
    system_global_interrupts_x5_lfsrReg_97[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_97 = system_global_interrupts_x5_lfsrReg_97[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_685 = {system_global_interrupts_x5_lfsrReg_hi_97,
    system_global_interrupts_x5_lfsrReg_lo_97};
  reg [15:0] system_global_interrupts_x5_lfsrReg_98;
  wire  system_global_interrupts_x5_lfsrReg_hi_98 = system_global_interrupts_x5_lfsrReg_98[0] ^
    system_global_interrupts_x5_lfsrReg_98[2] ^ system_global_interrupts_x5_lfsrReg_98[3] ^
    system_global_interrupts_x5_lfsrReg_98[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_98 = system_global_interrupts_x5_lfsrReg_98[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_692 = {system_global_interrupts_x5_lfsrReg_hi_98,
    system_global_interrupts_x5_lfsrReg_lo_98};
  reg [15:0] system_global_interrupts_x5_lfsrReg_99;
  wire  system_global_interrupts_x5_lfsrReg_hi_99 = system_global_interrupts_x5_lfsrReg_99[0] ^
    system_global_interrupts_x5_lfsrReg_99[2] ^ system_global_interrupts_x5_lfsrReg_99[3] ^
    system_global_interrupts_x5_lfsrReg_99[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_99 = system_global_interrupts_x5_lfsrReg_99[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_699 = {system_global_interrupts_x5_lfsrReg_hi_99,
    system_global_interrupts_x5_lfsrReg_lo_99};
  reg [15:0] system_global_interrupts_x5_lfsrReg_100;
  wire  system_global_interrupts_x5_lfsrReg_hi_100 = system_global_interrupts_x5_lfsrReg_100[0] ^
    system_global_interrupts_x5_lfsrReg_100[2] ^ system_global_interrupts_x5_lfsrReg_100[3] ^
    system_global_interrupts_x5_lfsrReg_100[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_100 = system_global_interrupts_x5_lfsrReg_100[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_706 = {system_global_interrupts_x5_lfsrReg_hi_100,
    system_global_interrupts_x5_lfsrReg_lo_100};
  reg [15:0] system_global_interrupts_x5_lfsrReg_101;
  wire  system_global_interrupts_x5_lfsrReg_hi_101 = system_global_interrupts_x5_lfsrReg_101[0] ^
    system_global_interrupts_x5_lfsrReg_101[2] ^ system_global_interrupts_x5_lfsrReg_101[3] ^
    system_global_interrupts_x5_lfsrReg_101[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_101 = system_global_interrupts_x5_lfsrReg_101[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_713 = {system_global_interrupts_x5_lfsrReg_hi_101,
    system_global_interrupts_x5_lfsrReg_lo_101};
  reg [15:0] system_global_interrupts_x5_lfsrReg_102;
  wire  system_global_interrupts_x5_lfsrReg_hi_102 = system_global_interrupts_x5_lfsrReg_102[0] ^
    system_global_interrupts_x5_lfsrReg_102[2] ^ system_global_interrupts_x5_lfsrReg_102[3] ^
    system_global_interrupts_x5_lfsrReg_102[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_102 = system_global_interrupts_x5_lfsrReg_102[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_720 = {system_global_interrupts_x5_lfsrReg_hi_102,
    system_global_interrupts_x5_lfsrReg_lo_102};
  reg [15:0] system_global_interrupts_x5_lfsrReg_103;
  wire  system_global_interrupts_x5_lfsrReg_hi_103 = system_global_interrupts_x5_lfsrReg_103[0] ^
    system_global_interrupts_x5_lfsrReg_103[2] ^ system_global_interrupts_x5_lfsrReg_103[3] ^
    system_global_interrupts_x5_lfsrReg_103[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_103 = system_global_interrupts_x5_lfsrReg_103[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_727 = {system_global_interrupts_x5_lfsrReg_hi_103,
    system_global_interrupts_x5_lfsrReg_lo_103};
  reg [15:0] system_global_interrupts_x5_lfsrReg_104;
  wire  system_global_interrupts_x5_lfsrReg_hi_104 = system_global_interrupts_x5_lfsrReg_104[0] ^
    system_global_interrupts_x5_lfsrReg_104[2] ^ system_global_interrupts_x5_lfsrReg_104[3] ^
    system_global_interrupts_x5_lfsrReg_104[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_104 = system_global_interrupts_x5_lfsrReg_104[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_734 = {system_global_interrupts_x5_lfsrReg_hi_104,
    system_global_interrupts_x5_lfsrReg_lo_104};
  reg [15:0] system_global_interrupts_x5_lfsrReg_105;
  wire  system_global_interrupts_x5_lfsrReg_hi_105 = system_global_interrupts_x5_lfsrReg_105[0] ^
    system_global_interrupts_x5_lfsrReg_105[2] ^ system_global_interrupts_x5_lfsrReg_105[3] ^
    system_global_interrupts_x5_lfsrReg_105[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_105 = system_global_interrupts_x5_lfsrReg_105[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_741 = {system_global_interrupts_x5_lfsrReg_hi_105,
    system_global_interrupts_x5_lfsrReg_lo_105};
  reg [15:0] system_global_interrupts_x5_lfsrReg_106;
  wire  system_global_interrupts_x5_lfsrReg_hi_106 = system_global_interrupts_x5_lfsrReg_106[0] ^
    system_global_interrupts_x5_lfsrReg_106[2] ^ system_global_interrupts_x5_lfsrReg_106[3] ^
    system_global_interrupts_x5_lfsrReg_106[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_106 = system_global_interrupts_x5_lfsrReg_106[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_748 = {system_global_interrupts_x5_lfsrReg_hi_106,
    system_global_interrupts_x5_lfsrReg_lo_106};
  reg [15:0] system_global_interrupts_x5_lfsrReg_107;
  wire  system_global_interrupts_x5_lfsrReg_hi_107 = system_global_interrupts_x5_lfsrReg_107[0] ^
    system_global_interrupts_x5_lfsrReg_107[2] ^ system_global_interrupts_x5_lfsrReg_107[3] ^
    system_global_interrupts_x5_lfsrReg_107[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_107 = system_global_interrupts_x5_lfsrReg_107[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_755 = {system_global_interrupts_x5_lfsrReg_hi_107,
    system_global_interrupts_x5_lfsrReg_lo_107};
  reg [15:0] system_global_interrupts_x5_lfsrReg_108;
  wire  system_global_interrupts_x5_lfsrReg_hi_108 = system_global_interrupts_x5_lfsrReg_108[0] ^
    system_global_interrupts_x5_lfsrReg_108[2] ^ system_global_interrupts_x5_lfsrReg_108[3] ^
    system_global_interrupts_x5_lfsrReg_108[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_108 = system_global_interrupts_x5_lfsrReg_108[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_762 = {system_global_interrupts_x5_lfsrReg_hi_108,
    system_global_interrupts_x5_lfsrReg_lo_108};
  reg [15:0] system_global_interrupts_x5_lfsrReg_109;
  wire  system_global_interrupts_x5_lfsrReg_hi_109 = system_global_interrupts_x5_lfsrReg_109[0] ^
    system_global_interrupts_x5_lfsrReg_109[2] ^ system_global_interrupts_x5_lfsrReg_109[3] ^
    system_global_interrupts_x5_lfsrReg_109[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_109 = system_global_interrupts_x5_lfsrReg_109[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_769 = {system_global_interrupts_x5_lfsrReg_hi_109,
    system_global_interrupts_x5_lfsrReg_lo_109};
  reg [15:0] system_global_interrupts_x5_lfsrReg_110;
  wire  system_global_interrupts_x5_lfsrReg_hi_110 = system_global_interrupts_x5_lfsrReg_110[0] ^
    system_global_interrupts_x5_lfsrReg_110[2] ^ system_global_interrupts_x5_lfsrReg_110[3] ^
    system_global_interrupts_x5_lfsrReg_110[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_110 = system_global_interrupts_x5_lfsrReg_110[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_776 = {system_global_interrupts_x5_lfsrReg_hi_110,
    system_global_interrupts_x5_lfsrReg_lo_110};
  reg [15:0] system_global_interrupts_x5_lfsrReg_111;
  wire  system_global_interrupts_x5_lfsrReg_hi_111 = system_global_interrupts_x5_lfsrReg_111[0] ^
    system_global_interrupts_x5_lfsrReg_111[2] ^ system_global_interrupts_x5_lfsrReg_111[3] ^
    system_global_interrupts_x5_lfsrReg_111[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_111 = system_global_interrupts_x5_lfsrReg_111[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_783 = {system_global_interrupts_x5_lfsrReg_hi_111,
    system_global_interrupts_x5_lfsrReg_lo_111};
  reg [15:0] system_global_interrupts_x5_lfsrReg_112;
  wire  system_global_interrupts_x5_lfsrReg_hi_112 = system_global_interrupts_x5_lfsrReg_112[0] ^
    system_global_interrupts_x5_lfsrReg_112[2] ^ system_global_interrupts_x5_lfsrReg_112[3] ^
    system_global_interrupts_x5_lfsrReg_112[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_112 = system_global_interrupts_x5_lfsrReg_112[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_790 = {system_global_interrupts_x5_lfsrReg_hi_112,
    system_global_interrupts_x5_lfsrReg_lo_112};
  reg [15:0] system_global_interrupts_x5_lfsrReg_113;
  wire  system_global_interrupts_x5_lfsrReg_hi_113 = system_global_interrupts_x5_lfsrReg_113[0] ^
    system_global_interrupts_x5_lfsrReg_113[2] ^ system_global_interrupts_x5_lfsrReg_113[3] ^
    system_global_interrupts_x5_lfsrReg_113[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_113 = system_global_interrupts_x5_lfsrReg_113[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_797 = {system_global_interrupts_x5_lfsrReg_hi_113,
    system_global_interrupts_x5_lfsrReg_lo_113};
  reg [15:0] system_global_interrupts_x5_lfsrReg_114;
  wire  system_global_interrupts_x5_lfsrReg_hi_114 = system_global_interrupts_x5_lfsrReg_114[0] ^
    system_global_interrupts_x5_lfsrReg_114[2] ^ system_global_interrupts_x5_lfsrReg_114[3] ^
    system_global_interrupts_x5_lfsrReg_114[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_114 = system_global_interrupts_x5_lfsrReg_114[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_804 = {system_global_interrupts_x5_lfsrReg_hi_114,
    system_global_interrupts_x5_lfsrReg_lo_114};
  reg [15:0] system_global_interrupts_x5_lfsrReg_115;
  wire  system_global_interrupts_x5_lfsrReg_hi_115 = system_global_interrupts_x5_lfsrReg_115[0] ^
    system_global_interrupts_x5_lfsrReg_115[2] ^ system_global_interrupts_x5_lfsrReg_115[3] ^
    system_global_interrupts_x5_lfsrReg_115[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_115 = system_global_interrupts_x5_lfsrReg_115[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_811 = {system_global_interrupts_x5_lfsrReg_hi_115,
    system_global_interrupts_x5_lfsrReg_lo_115};
  reg [15:0] system_global_interrupts_x5_lfsrReg_116;
  wire  system_global_interrupts_x5_lfsrReg_hi_116 = system_global_interrupts_x5_lfsrReg_116[0] ^
    system_global_interrupts_x5_lfsrReg_116[2] ^ system_global_interrupts_x5_lfsrReg_116[3] ^
    system_global_interrupts_x5_lfsrReg_116[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_116 = system_global_interrupts_x5_lfsrReg_116[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_818 = {system_global_interrupts_x5_lfsrReg_hi_116,
    system_global_interrupts_x5_lfsrReg_lo_116};
  reg [15:0] system_global_interrupts_x5_lfsrReg_117;
  wire  system_global_interrupts_x5_lfsrReg_hi_117 = system_global_interrupts_x5_lfsrReg_117[0] ^
    system_global_interrupts_x5_lfsrReg_117[2] ^ system_global_interrupts_x5_lfsrReg_117[3] ^
    system_global_interrupts_x5_lfsrReg_117[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_117 = system_global_interrupts_x5_lfsrReg_117[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_825 = {system_global_interrupts_x5_lfsrReg_hi_117,
    system_global_interrupts_x5_lfsrReg_lo_117};
  reg [15:0] system_global_interrupts_x5_lfsrReg_118;
  wire  system_global_interrupts_x5_lfsrReg_hi_118 = system_global_interrupts_x5_lfsrReg_118[0] ^
    system_global_interrupts_x5_lfsrReg_118[2] ^ system_global_interrupts_x5_lfsrReg_118[3] ^
    system_global_interrupts_x5_lfsrReg_118[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_118 = system_global_interrupts_x5_lfsrReg_118[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_832 = {system_global_interrupts_x5_lfsrReg_hi_118,
    system_global_interrupts_x5_lfsrReg_lo_118};
  reg [15:0] system_global_interrupts_x5_lfsrReg_119;
  wire  system_global_interrupts_x5_lfsrReg_hi_119 = system_global_interrupts_x5_lfsrReg_119[0] ^
    system_global_interrupts_x5_lfsrReg_119[2] ^ system_global_interrupts_x5_lfsrReg_119[3] ^
    system_global_interrupts_x5_lfsrReg_119[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_119 = system_global_interrupts_x5_lfsrReg_119[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_839 = {system_global_interrupts_x5_lfsrReg_hi_119,
    system_global_interrupts_x5_lfsrReg_lo_119};
  reg [15:0] system_global_interrupts_x5_lfsrReg_120;
  wire  system_global_interrupts_x5_lfsrReg_hi_120 = system_global_interrupts_x5_lfsrReg_120[0] ^
    system_global_interrupts_x5_lfsrReg_120[2] ^ system_global_interrupts_x5_lfsrReg_120[3] ^
    system_global_interrupts_x5_lfsrReg_120[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_120 = system_global_interrupts_x5_lfsrReg_120[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_846 = {system_global_interrupts_x5_lfsrReg_hi_120,
    system_global_interrupts_x5_lfsrReg_lo_120};
  reg [15:0] system_global_interrupts_x5_lfsrReg_121;
  wire  system_global_interrupts_x5_lfsrReg_hi_121 = system_global_interrupts_x5_lfsrReg_121[0] ^
    system_global_interrupts_x5_lfsrReg_121[2] ^ system_global_interrupts_x5_lfsrReg_121[3] ^
    system_global_interrupts_x5_lfsrReg_121[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_121 = system_global_interrupts_x5_lfsrReg_121[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_853 = {system_global_interrupts_x5_lfsrReg_hi_121,
    system_global_interrupts_x5_lfsrReg_lo_121};
  reg [15:0] system_global_interrupts_x5_lfsrReg_122;
  wire  system_global_interrupts_x5_lfsrReg_hi_122 = system_global_interrupts_x5_lfsrReg_122[0] ^
    system_global_interrupts_x5_lfsrReg_122[2] ^ system_global_interrupts_x5_lfsrReg_122[3] ^
    system_global_interrupts_x5_lfsrReg_122[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_122 = system_global_interrupts_x5_lfsrReg_122[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_860 = {system_global_interrupts_x5_lfsrReg_hi_122,
    system_global_interrupts_x5_lfsrReg_lo_122};
  reg [15:0] system_global_interrupts_x5_lfsrReg_123;
  wire  system_global_interrupts_x5_lfsrReg_hi_123 = system_global_interrupts_x5_lfsrReg_123[0] ^
    system_global_interrupts_x5_lfsrReg_123[2] ^ system_global_interrupts_x5_lfsrReg_123[3] ^
    system_global_interrupts_x5_lfsrReg_123[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_123 = system_global_interrupts_x5_lfsrReg_123[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_867 = {system_global_interrupts_x5_lfsrReg_hi_123,
    system_global_interrupts_x5_lfsrReg_lo_123};
  reg [15:0] system_global_interrupts_x5_lfsrReg_124;
  wire  system_global_interrupts_x5_lfsrReg_hi_124 = system_global_interrupts_x5_lfsrReg_124[0] ^
    system_global_interrupts_x5_lfsrReg_124[2] ^ system_global_interrupts_x5_lfsrReg_124[3] ^
    system_global_interrupts_x5_lfsrReg_124[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_124 = system_global_interrupts_x5_lfsrReg_124[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_874 = {system_global_interrupts_x5_lfsrReg_hi_124,
    system_global_interrupts_x5_lfsrReg_lo_124};
  reg [15:0] system_global_interrupts_x5_lfsrReg_125;
  wire  system_global_interrupts_x5_lfsrReg_hi_125 = system_global_interrupts_x5_lfsrReg_125[0] ^
    system_global_interrupts_x5_lfsrReg_125[2] ^ system_global_interrupts_x5_lfsrReg_125[3] ^
    system_global_interrupts_x5_lfsrReg_125[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_125 = system_global_interrupts_x5_lfsrReg_125[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_881 = {system_global_interrupts_x5_lfsrReg_hi_125,
    system_global_interrupts_x5_lfsrReg_lo_125};
  reg [15:0] system_global_interrupts_x5_lfsrReg_126;
  wire  system_global_interrupts_x5_lfsrReg_hi_126 = system_global_interrupts_x5_lfsrReg_126[0] ^
    system_global_interrupts_x5_lfsrReg_126[2] ^ system_global_interrupts_x5_lfsrReg_126[3] ^
    system_global_interrupts_x5_lfsrReg_126[5];
  wire [14:0] system_global_interrupts_x5_lfsrReg_lo_126 = system_global_interrupts_x5_lfsrReg_126[15:1];
  wire [15:0] _system_global_interrupts_x5_lfsrReg_T_888 = {system_global_interrupts_x5_lfsrReg_hi_126,
    system_global_interrupts_x5_lfsrReg_lo_126};
  wire [6:0] system_global_interrupts_lo_lo_lo_lo_1 = {system_global_interrupts_x5_lfsrReg_6[0],
    system_global_interrupts_x5_lfsrReg_5[0],system_global_interrupts_x5_lfsrReg_4[0],
    system_global_interrupts_x5_lfsrReg_3[0],system_global_interrupts_x5_lfsrReg_2[0],
    system_global_interrupts_x5_lfsrReg_1[0],system_global_interrupts_x5_lfsrReg[0]};
  wire [14:0] system_global_interrupts_lo_lo_lo_1 = {system_global_interrupts_x5_lfsrReg_14[0],
    system_global_interrupts_x5_lfsrReg_13[0],system_global_interrupts_x5_lfsrReg_12[0],
    system_global_interrupts_x5_lfsrReg_11[0],system_global_interrupts_x5_lfsrReg_10[0],
    system_global_interrupts_x5_lfsrReg_9[0],system_global_interrupts_x5_lfsrReg_8[0],
    system_global_interrupts_x5_lfsrReg_7[0],system_global_interrupts_lo_lo_lo_lo_1};
  wire [7:0] system_global_interrupts_lo_lo_hi_lo_1 = {system_global_interrupts_x5_lfsrReg_22[0],
    system_global_interrupts_x5_lfsrReg_21[0],system_global_interrupts_x5_lfsrReg_20[0],
    system_global_interrupts_x5_lfsrReg_19[0],system_global_interrupts_x5_lfsrReg_18[0],
    system_global_interrupts_x5_lfsrReg_17[0],system_global_interrupts_x5_lfsrReg_16[0],
    system_global_interrupts_x5_lfsrReg_15[0]};
  wire [30:0] system_global_interrupts_lo_lo_1 = {system_global_interrupts_x5_lfsrReg_30[0],
    system_global_interrupts_x5_lfsrReg_29[0],system_global_interrupts_x5_lfsrReg_28[0],
    system_global_interrupts_x5_lfsrReg_27[0],system_global_interrupts_x5_lfsrReg_26[0],
    system_global_interrupts_x5_lfsrReg_25[0],system_global_interrupts_x5_lfsrReg_24[0],
    system_global_interrupts_x5_lfsrReg_23[0],system_global_interrupts_lo_lo_hi_lo_1,system_global_interrupts_lo_lo_lo_1
    };
  wire [7:0] system_global_interrupts_lo_hi_lo_lo_1 = {system_global_interrupts_x5_lfsrReg_38[0],
    system_global_interrupts_x5_lfsrReg_37[0],system_global_interrupts_x5_lfsrReg_36[0],
    system_global_interrupts_x5_lfsrReg_35[0],system_global_interrupts_x5_lfsrReg_34[0],
    system_global_interrupts_x5_lfsrReg_33[0],system_global_interrupts_x5_lfsrReg_32[0],
    system_global_interrupts_x5_lfsrReg_31[0]};
  wire [15:0] system_global_interrupts_lo_hi_lo_1 = {system_global_interrupts_x5_lfsrReg_46[0],
    system_global_interrupts_x5_lfsrReg_45[0],system_global_interrupts_x5_lfsrReg_44[0],
    system_global_interrupts_x5_lfsrReg_43[0],system_global_interrupts_x5_lfsrReg_42[0],
    system_global_interrupts_x5_lfsrReg_41[0],system_global_interrupts_x5_lfsrReg_40[0],
    system_global_interrupts_x5_lfsrReg_39[0],system_global_interrupts_lo_hi_lo_lo_1};
  wire [7:0] system_global_interrupts_lo_hi_hi_lo_1 = {system_global_interrupts_x5_lfsrReg_54[0],
    system_global_interrupts_x5_lfsrReg_53[0],system_global_interrupts_x5_lfsrReg_52[0],
    system_global_interrupts_x5_lfsrReg_51[0],system_global_interrupts_x5_lfsrReg_50[0],
    system_global_interrupts_x5_lfsrReg_49[0],system_global_interrupts_x5_lfsrReg_48[0],
    system_global_interrupts_x5_lfsrReg_47[0]};
  wire [31:0] system_global_interrupts_lo_hi_1 = {system_global_interrupts_x5_lfsrReg_62[0],
    system_global_interrupts_x5_lfsrReg_61[0],system_global_interrupts_x5_lfsrReg_60[0],
    system_global_interrupts_x5_lfsrReg_59[0],system_global_interrupts_x5_lfsrReg_58[0],
    system_global_interrupts_x5_lfsrReg_57[0],system_global_interrupts_x5_lfsrReg_56[0],
    system_global_interrupts_x5_lfsrReg_55[0],system_global_interrupts_lo_hi_hi_lo_1,system_global_interrupts_lo_hi_lo_1
    };
  wire [7:0] system_global_interrupts_hi_lo_lo_lo_1 = {system_global_interrupts_x5_lfsrReg_70[0],
    system_global_interrupts_x5_lfsrReg_69[0],system_global_interrupts_x5_lfsrReg_68[0],
    system_global_interrupts_x5_lfsrReg_67[0],system_global_interrupts_x5_lfsrReg_66[0],
    system_global_interrupts_x5_lfsrReg_65[0],system_global_interrupts_x5_lfsrReg_64[0],
    system_global_interrupts_x5_lfsrReg_63[0]};
  wire [15:0] system_global_interrupts_hi_lo_lo_1 = {system_global_interrupts_x5_lfsrReg_78[0],
    system_global_interrupts_x5_lfsrReg_77[0],system_global_interrupts_x5_lfsrReg_76[0],
    system_global_interrupts_x5_lfsrReg_75[0],system_global_interrupts_x5_lfsrReg_74[0],
    system_global_interrupts_x5_lfsrReg_73[0],system_global_interrupts_x5_lfsrReg_72[0],
    system_global_interrupts_x5_lfsrReg_71[0],system_global_interrupts_hi_lo_lo_lo_1};
  wire [7:0] system_global_interrupts_hi_lo_hi_lo_1 = {system_global_interrupts_x5_lfsrReg_86[0],
    system_global_interrupts_x5_lfsrReg_85[0],system_global_interrupts_x5_lfsrReg_84[0],
    system_global_interrupts_x5_lfsrReg_83[0],system_global_interrupts_x5_lfsrReg_82[0],
    system_global_interrupts_x5_lfsrReg_81[0],system_global_interrupts_x5_lfsrReg_80[0],
    system_global_interrupts_x5_lfsrReg_79[0]};
  wire [31:0] system_global_interrupts_hi_lo_1 = {system_global_interrupts_x5_lfsrReg_94[0],
    system_global_interrupts_x5_lfsrReg_93[0],system_global_interrupts_x5_lfsrReg_92[0],
    system_global_interrupts_x5_lfsrReg_91[0],system_global_interrupts_x5_lfsrReg_90[0],
    system_global_interrupts_x5_lfsrReg_89[0],system_global_interrupts_x5_lfsrReg_88[0],
    system_global_interrupts_x5_lfsrReg_87[0],system_global_interrupts_hi_lo_hi_lo_1,system_global_interrupts_hi_lo_lo_1
    };
  wire [7:0] system_global_interrupts_hi_hi_lo_lo_1 = {system_global_interrupts_x5_lfsrReg_102[0],
    system_global_interrupts_x5_lfsrReg_101[0],system_global_interrupts_x5_lfsrReg_100[0],
    system_global_interrupts_x5_lfsrReg_99[0],system_global_interrupts_x5_lfsrReg_98[0],
    system_global_interrupts_x5_lfsrReg_97[0],system_global_interrupts_x5_lfsrReg_96[0],
    system_global_interrupts_x5_lfsrReg_95[0]};
  wire [15:0] system_global_interrupts_hi_hi_lo_1 = {system_global_interrupts_x5_lfsrReg_110[0],
    system_global_interrupts_x5_lfsrReg_109[0],system_global_interrupts_x5_lfsrReg_108[0],
    system_global_interrupts_x5_lfsrReg_107[0],system_global_interrupts_x5_lfsrReg_106[0],
    system_global_interrupts_x5_lfsrReg_105[0],system_global_interrupts_x5_lfsrReg_104[0],
    system_global_interrupts_x5_lfsrReg_103[0],system_global_interrupts_hi_hi_lo_lo_1};
  wire [7:0] system_global_interrupts_hi_hi_hi_lo_1 = {system_global_interrupts_x5_lfsrReg_118[0],
    system_global_interrupts_x5_lfsrReg_117[0],system_global_interrupts_x5_lfsrReg_116[0],
    system_global_interrupts_x5_lfsrReg_115[0],system_global_interrupts_x5_lfsrReg_114[0],
    system_global_interrupts_x5_lfsrReg_113[0],system_global_interrupts_x5_lfsrReg_112[0],
    system_global_interrupts_x5_lfsrReg_111[0]};
  wire [31:0] system_global_interrupts_hi_hi_1 = {system_global_interrupts_x5_lfsrReg_126[0],
    system_global_interrupts_x5_lfsrReg_125[0],system_global_interrupts_x5_lfsrReg_124[0],
    system_global_interrupts_x5_lfsrReg_123[0],system_global_interrupts_x5_lfsrReg_122[0],
    system_global_interrupts_x5_lfsrReg_121[0],system_global_interrupts_x5_lfsrReg_120[0],
    system_global_interrupts_x5_lfsrReg_119[0],system_global_interrupts_hi_hi_hi_lo_1,
    system_global_interrupts_hi_hi_lo_1};
  wire [126:0] _system_global_interrupts_T_3 = {system_global_interrupts_hi_hi_1,system_global_interrupts_hi_lo_1,
    system_global_interrupts_lo_hi_1,system_global_interrupts_lo_lo_1};
  wire [126:0] _GEN_519 = drive_interrupt_type == 32'h4 ? _system_global_interrupts_T_3 : 127'h0;
  wire [127:0] _GEN_520 = drive_interrupt_type == 32'h3 ? _system_global_interrupts_T_2 : {{1'd0}, _GEN_519};
  wire [127:0] _GEN_521 = drive_interrupt_type == 32'h2 ? 128'h2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa : _GEN_520;
  wire [127:0] _GEN_522 = drive_interrupt_type == 32'h1 ? 128'h7fffffffffffffffffffffffffffffff : _GEN_521;
  wire [127:0] _GEN_523 = drive_interrupt_type == 32'h0 ? 128'h0 : _GEN_522;
  reg [6:0] tick_value_1;
  wire  tick_1 = tick_value_1 == 7'h63;
  wire [6:0] _tick_value_T_3 = tick_value_1 + 7'h1;
  wire [31:0] drive_interrupt_type_1 = plusarg_reader_3_out;
  reg [3:0] system_local_interrupts_0_value;
  wire [3:0] _system_local_interrupts_0_wrap_value_T_1 = system_local_interrupts_0_value + 4'h1;
  wire [15:0] _system_local_interrupts_0_T_2 = 16'h1 << system_local_interrupts_0_value;
  reg [15:0] tickers_x3_lfsrReg_127;
  wire  tickers_x3_lfsrReg_hi_127 = tickers_x3_lfsrReg_127[0] ^ tickers_x3_lfsrReg_127[2] ^ tickers_x3_lfsrReg_127[3] ^
    tickers_x3_lfsrReg_127[5];
  wire [14:0] tickers_x3_lfsrReg_lo_127 = tickers_x3_lfsrReg_127[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_895 = {tickers_x3_lfsrReg_hi_127,tickers_x3_lfsrReg_lo_127};
  reg [15:0] tickers_x3_lfsrReg_128;
  wire  tickers_x3_lfsrReg_hi_128 = tickers_x3_lfsrReg_128[0] ^ tickers_x3_lfsrReg_128[2] ^ tickers_x3_lfsrReg_128[3] ^
    tickers_x3_lfsrReg_128[5];
  wire [14:0] tickers_x3_lfsrReg_lo_128 = tickers_x3_lfsrReg_128[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_902 = {tickers_x3_lfsrReg_hi_128,tickers_x3_lfsrReg_lo_128};
  reg [15:0] tickers_x3_lfsrReg_129;
  wire  tickers_x3_lfsrReg_hi_129 = tickers_x3_lfsrReg_129[0] ^ tickers_x3_lfsrReg_129[2] ^ tickers_x3_lfsrReg_129[3] ^
    tickers_x3_lfsrReg_129[5];
  wire [14:0] tickers_x3_lfsrReg_lo_129 = tickers_x3_lfsrReg_129[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_909 = {tickers_x3_lfsrReg_hi_129,tickers_x3_lfsrReg_lo_129};
  reg [15:0] tickers_x3_lfsrReg_130;
  wire  tickers_x3_lfsrReg_hi_130 = tickers_x3_lfsrReg_130[0] ^ tickers_x3_lfsrReg_130[2] ^ tickers_x3_lfsrReg_130[3] ^
    tickers_x3_lfsrReg_130[5];
  wire [14:0] tickers_x3_lfsrReg_lo_130 = tickers_x3_lfsrReg_130[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_916 = {tickers_x3_lfsrReg_hi_130,tickers_x3_lfsrReg_lo_130};
  reg [15:0] tickers_x3_lfsrReg_131;
  wire  tickers_x3_lfsrReg_hi_131 = tickers_x3_lfsrReg_131[0] ^ tickers_x3_lfsrReg_131[2] ^ tickers_x3_lfsrReg_131[3] ^
    tickers_x3_lfsrReg_131[5];
  wire [14:0] tickers_x3_lfsrReg_lo_131 = tickers_x3_lfsrReg_131[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_923 = {tickers_x3_lfsrReg_hi_131,tickers_x3_lfsrReg_lo_131};
  reg [15:0] tickers_x3_lfsrReg_132;
  wire  tickers_x3_lfsrReg_hi_132 = tickers_x3_lfsrReg_132[0] ^ tickers_x3_lfsrReg_132[2] ^ tickers_x3_lfsrReg_132[3] ^
    tickers_x3_lfsrReg_132[5];
  wire [14:0] tickers_x3_lfsrReg_lo_132 = tickers_x3_lfsrReg_132[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_930 = {tickers_x3_lfsrReg_hi_132,tickers_x3_lfsrReg_lo_132};
  reg [15:0] tickers_x3_lfsrReg_133;
  wire  tickers_x3_lfsrReg_hi_133 = tickers_x3_lfsrReg_133[0] ^ tickers_x3_lfsrReg_133[2] ^ tickers_x3_lfsrReg_133[3] ^
    tickers_x3_lfsrReg_133[5];
  wire [14:0] tickers_x3_lfsrReg_lo_133 = tickers_x3_lfsrReg_133[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_937 = {tickers_x3_lfsrReg_hi_133,tickers_x3_lfsrReg_lo_133};
  reg [15:0] tickers_x3_lfsrReg_134;
  wire  tickers_x3_lfsrReg_hi_134 = tickers_x3_lfsrReg_134[0] ^ tickers_x3_lfsrReg_134[2] ^ tickers_x3_lfsrReg_134[3] ^
    tickers_x3_lfsrReg_134[5];
  wire [14:0] tickers_x3_lfsrReg_lo_134 = tickers_x3_lfsrReg_134[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_944 = {tickers_x3_lfsrReg_hi_134,tickers_x3_lfsrReg_lo_134};
  reg [15:0] tickers_x3_lfsrReg_135;
  wire  tickers_x3_lfsrReg_hi_135 = tickers_x3_lfsrReg_135[0] ^ tickers_x3_lfsrReg_135[2] ^ tickers_x3_lfsrReg_135[3] ^
    tickers_x3_lfsrReg_135[5];
  wire [14:0] tickers_x3_lfsrReg_lo_135 = tickers_x3_lfsrReg_135[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_951 = {tickers_x3_lfsrReg_hi_135,tickers_x3_lfsrReg_lo_135};
  reg [15:0] tickers_x3_lfsrReg_136;
  wire  tickers_x3_lfsrReg_hi_136 = tickers_x3_lfsrReg_136[0] ^ tickers_x3_lfsrReg_136[2] ^ tickers_x3_lfsrReg_136[3] ^
    tickers_x3_lfsrReg_136[5];
  wire [14:0] tickers_x3_lfsrReg_lo_136 = tickers_x3_lfsrReg_136[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_958 = {tickers_x3_lfsrReg_hi_136,tickers_x3_lfsrReg_lo_136};
  reg [15:0] tickers_x3_lfsrReg_137;
  wire  tickers_x3_lfsrReg_hi_137 = tickers_x3_lfsrReg_137[0] ^ tickers_x3_lfsrReg_137[2] ^ tickers_x3_lfsrReg_137[3] ^
    tickers_x3_lfsrReg_137[5];
  wire [14:0] tickers_x3_lfsrReg_lo_137 = tickers_x3_lfsrReg_137[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_965 = {tickers_x3_lfsrReg_hi_137,tickers_x3_lfsrReg_lo_137};
  reg [15:0] tickers_x3_lfsrReg_138;
  wire  tickers_x3_lfsrReg_hi_138 = tickers_x3_lfsrReg_138[0] ^ tickers_x3_lfsrReg_138[2] ^ tickers_x3_lfsrReg_138[3] ^
    tickers_x3_lfsrReg_138[5];
  wire [14:0] tickers_x3_lfsrReg_lo_138 = tickers_x3_lfsrReg_138[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_972 = {tickers_x3_lfsrReg_hi_138,tickers_x3_lfsrReg_lo_138};
  reg [15:0] tickers_x3_lfsrReg_139;
  wire  tickers_x3_lfsrReg_hi_139 = tickers_x3_lfsrReg_139[0] ^ tickers_x3_lfsrReg_139[2] ^ tickers_x3_lfsrReg_139[3] ^
    tickers_x3_lfsrReg_139[5];
  wire [14:0] tickers_x3_lfsrReg_lo_139 = tickers_x3_lfsrReg_139[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_979 = {tickers_x3_lfsrReg_hi_139,tickers_x3_lfsrReg_lo_139};
  reg [15:0] tickers_x3_lfsrReg_140;
  wire  tickers_x3_lfsrReg_hi_140 = tickers_x3_lfsrReg_140[0] ^ tickers_x3_lfsrReg_140[2] ^ tickers_x3_lfsrReg_140[3] ^
    tickers_x3_lfsrReg_140[5];
  wire [14:0] tickers_x3_lfsrReg_lo_140 = tickers_x3_lfsrReg_140[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_986 = {tickers_x3_lfsrReg_hi_140,tickers_x3_lfsrReg_lo_140};
  reg [15:0] tickers_x3_lfsrReg_141;
  wire  tickers_x3_lfsrReg_hi_141 = tickers_x3_lfsrReg_141[0] ^ tickers_x3_lfsrReg_141[2] ^ tickers_x3_lfsrReg_141[3] ^
    tickers_x3_lfsrReg_141[5];
  wire [14:0] tickers_x3_lfsrReg_lo_141 = tickers_x3_lfsrReg_141[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_993 = {tickers_x3_lfsrReg_hi_141,tickers_x3_lfsrReg_lo_141};
  reg [15:0] tickers_x3_lfsrReg_142;
  wire  tickers_x3_lfsrReg_hi_142 = tickers_x3_lfsrReg_142[0] ^ tickers_x3_lfsrReg_142[2] ^ tickers_x3_lfsrReg_142[3] ^
    tickers_x3_lfsrReg_142[5];
  wire [14:0] tickers_x3_lfsrReg_lo_142 = tickers_x3_lfsrReg_142[15:1];
  wire [15:0] _tickers_x3_lfsrReg_T_1000 = {tickers_x3_lfsrReg_hi_142,tickers_x3_lfsrReg_lo_142};
  wire [7:0] system_local_interrupts_0_lo_1 = {tickers_x3_lfsrReg_134[0],tickers_x3_lfsrReg_133[0],
    tickers_x3_lfsrReg_132[0],tickers_x3_lfsrReg_131[0],tickers_x3_lfsrReg_130[0],tickers_x3_lfsrReg_129[0],
    tickers_x3_lfsrReg_128[0],tickers_x3_lfsrReg_127[0]};
  wire [15:0] _system_local_interrupts_0_T_3 = {tickers_x3_lfsrReg_142[0],tickers_x3_lfsrReg_141[0],
    tickers_x3_lfsrReg_140[0],tickers_x3_lfsrReg_139[0],tickers_x3_lfsrReg_138[0],tickers_x3_lfsrReg_137[0],
    tickers_x3_lfsrReg_136[0],tickers_x3_lfsrReg_135[0],system_local_interrupts_0_lo_1};
  reg [15:0] tickers_x5_lfsrReg;
  wire  tickers_x5_lfsrReg_hi = tickers_x5_lfsrReg[0] ^ tickers_x5_lfsrReg[2] ^ tickers_x5_lfsrReg[3] ^
    tickers_x5_lfsrReg[5];
  wire [14:0] tickers_x5_lfsrReg_lo = tickers_x5_lfsrReg[15:1];
  wire [15:0] _tickers_x5_lfsrReg_T_6 = {tickers_x5_lfsrReg_hi,tickers_x5_lfsrReg_lo};
  reg [15:0] tickers_x5_lfsrReg_1;
  wire  tickers_x5_lfsrReg_hi_1 = tickers_x5_lfsrReg_1[0] ^ tickers_x5_lfsrReg_1[2] ^ tickers_x5_lfsrReg_1[3] ^
    tickers_x5_lfsrReg_1[5];
  wire [14:0] tickers_x5_lfsrReg_lo_1 = tickers_x5_lfsrReg_1[15:1];
  wire [15:0] _tickers_x5_lfsrReg_T_13 = {tickers_x5_lfsrReg_hi_1,tickers_x5_lfsrReg_lo_1};
  reg [15:0] tickers_x5_lfsrReg_2;
  wire  tickers_x5_lfsrReg_hi_2 = tickers_x5_lfsrReg_2[0] ^ tickers_x5_lfsrReg_2[2] ^ tickers_x5_lfsrReg_2[3] ^
    tickers_x5_lfsrReg_2[5];
  wire [14:0] tickers_x5_lfsrReg_lo_2 = tickers_x5_lfsrReg_2[15:1];
  wire [15:0] _tickers_x5_lfsrReg_T_20 = {tickers_x5_lfsrReg_hi_2,tickers_x5_lfsrReg_lo_2};
  reg [15:0] tickers_x5_lfsrReg_3;
  wire  tickers_x5_lfsrReg_hi_3 = tickers_x5_lfsrReg_3[0] ^ tickers_x5_lfsrReg_3[2] ^ tickers_x5_lfsrReg_3[3] ^
    tickers_x5_lfsrReg_3[5];
  wire [14:0] tickers_x5_lfsrReg_lo_3 = tickers_x5_lfsrReg_3[15:1];
  wire [15:0] _tickers_x5_lfsrReg_T_27 = {tickers_x5_lfsrReg_hi_3,tickers_x5_lfsrReg_lo_3};
  reg [15:0] tickers_x5_lfsrReg_4;
  wire  tickers_x5_lfsrReg_hi_4 = tickers_x5_lfsrReg_4[0] ^ tickers_x5_lfsrReg_4[2] ^ tickers_x5_lfsrReg_4[3] ^
    tickers_x5_lfsrReg_4[5];
  wire [14:0] tickers_x5_lfsrReg_lo_4 = tickers_x5_lfsrReg_4[15:1];
  wire [15:0] _tickers_x5_lfsrReg_T_34 = {tickers_x5_lfsrReg_hi_4,tickers_x5_lfsrReg_lo_4};
  reg [15:0] tickers_x5_lfsrReg_5;
  wire  tickers_x5_lfsrReg_hi_5 = tickers_x5_lfsrReg_5[0] ^ tickers_x5_lfsrReg_5[2] ^ tickers_x5_lfsrReg_5[3] ^
    tickers_x5_lfsrReg_5[5];
  wire [14:0] tickers_x5_lfsrReg_lo_5 = tickers_x5_lfsrReg_5[15:1];
  wire [15:0] _tickers_x5_lfsrReg_T_41 = {tickers_x5_lfsrReg_hi_5,tickers_x5_lfsrReg_lo_5};
  reg [15:0] tickers_x5_lfsrReg_6;
  wire  tickers_x5_lfsrReg_hi_6 = tickers_x5_lfsrReg_6[0] ^ tickers_x5_lfsrReg_6[2] ^ tickers_x5_lfsrReg_6[3] ^
    tickers_x5_lfsrReg_6[5];
  wire [14:0] tickers_x5_lfsrReg_lo_6 = tickers_x5_lfsrReg_6[15:1];
  wire [15:0] _tickers_x5_lfsrReg_T_48 = {tickers_x5_lfsrReg_hi_6,tickers_x5_lfsrReg_lo_6};
  reg [15:0] tickers_x5_lfsrReg_7;
  wire  tickers_x5_lfsrReg_hi_7 = tickers_x5_lfsrReg_7[0] ^ tickers_x5_lfsrReg_7[2] ^ tickers_x5_lfsrReg_7[3] ^
    tickers_x5_lfsrReg_7[5];
  wire [14:0] tickers_x5_lfsrReg_lo_7 = tickers_x5_lfsrReg_7[15:1];
  wire [15:0] _tickers_x5_lfsrReg_T_55 = {tickers_x5_lfsrReg_hi_7,tickers_x5_lfsrReg_lo_7};
  reg [15:0] tickers_x5_lfsrReg_8;
  wire  tickers_x5_lfsrReg_hi_8 = tickers_x5_lfsrReg_8[0] ^ tickers_x5_lfsrReg_8[2] ^ tickers_x5_lfsrReg_8[3] ^
    tickers_x5_lfsrReg_8[5];
  wire [14:0] tickers_x5_lfsrReg_lo_8 = tickers_x5_lfsrReg_8[15:1];
  wire [15:0] _tickers_x5_lfsrReg_T_62 = {tickers_x5_lfsrReg_hi_8,tickers_x5_lfsrReg_lo_8};
  reg [15:0] tickers_x5_lfsrReg_9;
  wire  tickers_x5_lfsrReg_hi_9 = tickers_x5_lfsrReg_9[0] ^ tickers_x5_lfsrReg_9[2] ^ tickers_x5_lfsrReg_9[3] ^
    tickers_x5_lfsrReg_9[5];
  wire [14:0] tickers_x5_lfsrReg_lo_9 = tickers_x5_lfsrReg_9[15:1];
  wire [15:0] _tickers_x5_lfsrReg_T_69 = {tickers_x5_lfsrReg_hi_9,tickers_x5_lfsrReg_lo_9};
  reg [15:0] tickers_x5_lfsrReg_10;
  wire  tickers_x5_lfsrReg_hi_10 = tickers_x5_lfsrReg_10[0] ^ tickers_x5_lfsrReg_10[2] ^ tickers_x5_lfsrReg_10[3] ^
    tickers_x5_lfsrReg_10[5];
  wire [14:0] tickers_x5_lfsrReg_lo_10 = tickers_x5_lfsrReg_10[15:1];
  wire [15:0] _tickers_x5_lfsrReg_T_76 = {tickers_x5_lfsrReg_hi_10,tickers_x5_lfsrReg_lo_10};
  reg [15:0] tickers_x5_lfsrReg_11;
  wire  tickers_x5_lfsrReg_hi_11 = tickers_x5_lfsrReg_11[0] ^ tickers_x5_lfsrReg_11[2] ^ tickers_x5_lfsrReg_11[3] ^
    tickers_x5_lfsrReg_11[5];
  wire [14:0] tickers_x5_lfsrReg_lo_11 = tickers_x5_lfsrReg_11[15:1];
  wire [15:0] _tickers_x5_lfsrReg_T_83 = {tickers_x5_lfsrReg_hi_11,tickers_x5_lfsrReg_lo_11};
  reg [15:0] tickers_x5_lfsrReg_12;
  wire  tickers_x5_lfsrReg_hi_12 = tickers_x5_lfsrReg_12[0] ^ tickers_x5_lfsrReg_12[2] ^ tickers_x5_lfsrReg_12[3] ^
    tickers_x5_lfsrReg_12[5];
  wire [14:0] tickers_x5_lfsrReg_lo_12 = tickers_x5_lfsrReg_12[15:1];
  wire [15:0] _tickers_x5_lfsrReg_T_90 = {tickers_x5_lfsrReg_hi_12,tickers_x5_lfsrReg_lo_12};
  reg [15:0] tickers_x5_lfsrReg_13;
  wire  tickers_x5_lfsrReg_hi_13 = tickers_x5_lfsrReg_13[0] ^ tickers_x5_lfsrReg_13[2] ^ tickers_x5_lfsrReg_13[3] ^
    tickers_x5_lfsrReg_13[5];
  wire [14:0] tickers_x5_lfsrReg_lo_13 = tickers_x5_lfsrReg_13[15:1];
  wire [15:0] _tickers_x5_lfsrReg_T_97 = {tickers_x5_lfsrReg_hi_13,tickers_x5_lfsrReg_lo_13};
  reg [15:0] tickers_x5_lfsrReg_14;
  wire  tickers_x5_lfsrReg_hi_14 = tickers_x5_lfsrReg_14[0] ^ tickers_x5_lfsrReg_14[2] ^ tickers_x5_lfsrReg_14[3] ^
    tickers_x5_lfsrReg_14[5];
  wire [14:0] tickers_x5_lfsrReg_lo_14 = tickers_x5_lfsrReg_14[15:1];
  wire [15:0] _tickers_x5_lfsrReg_T_104 = {tickers_x5_lfsrReg_hi_14,tickers_x5_lfsrReg_lo_14};
  reg [15:0] tickers_x5_lfsrReg_15;
  wire  tickers_x5_lfsrReg_hi_15 = tickers_x5_lfsrReg_15[0] ^ tickers_x5_lfsrReg_15[2] ^ tickers_x5_lfsrReg_15[3] ^
    tickers_x5_lfsrReg_15[5];
  wire [14:0] tickers_x5_lfsrReg_lo_15 = tickers_x5_lfsrReg_15[15:1];
  wire [15:0] _tickers_x5_lfsrReg_T_111 = {tickers_x5_lfsrReg_hi_15,tickers_x5_lfsrReg_lo_15};
  wire [7:0] system_local_interrupts_0_lo_2 = {tickers_x5_lfsrReg_7[0],tickers_x5_lfsrReg_6[0],tickers_x5_lfsrReg_5[0],
    tickers_x5_lfsrReg_4[0],tickers_x5_lfsrReg_3[0],tickers_x5_lfsrReg_2[0],tickers_x5_lfsrReg_1[0],tickers_x5_lfsrReg[0
    ]};
  wire [15:0] _system_local_interrupts_0_T_4 = {tickers_x5_lfsrReg_15[0],tickers_x5_lfsrReg_14[0],tickers_x5_lfsrReg_13[
    0],tickers_x5_lfsrReg_12[0],tickers_x5_lfsrReg_11[0],tickers_x5_lfsrReg_10[0],tickers_x5_lfsrReg_9[0],
    tickers_x5_lfsrReg_8[0],system_local_interrupts_0_lo_2};
  wire [31:0] _GEN_591 = system_wfi_from_tile_0 ? dpi_drivers_0_interrupts : {{16'd0}, _system_local_interrupts_0_T_4};
  wire [31:0] _GEN_592 = drive_interrupt_type_1 == 32'h5 ? _GEN_591 : 32'h0;
  wire [31:0] _GEN_593 = drive_interrupt_type_1 == 32'h4 ? {{16'd0}, _system_local_interrupts_0_T_3} : _GEN_592;
  wire [31:0] _GEN_594 = drive_interrupt_type_1 == 32'h3 ? {{16'd0}, _system_local_interrupts_0_T_2} : _GEN_593;
  wire [31:0] _GEN_595 = drive_interrupt_type_1 == 32'h2 ? 32'haaaa : _GEN_594;
  wire [31:0] _GEN_596 = drive_interrupt_type_1 == 32'h1 ? 32'hffff : _GEN_595;
  wire [31:0] _GEN_597 = drive_interrupt_type_1 == 32'h0 ? dpi_drivers_0_interrupts : _GEN_596;
  wire  csrTraces_hartid = csrTraces_DataTap_1__0;
  SiFive_CoreIPSubsystem system (
    .clock(system_clock),
    .reset(system_reset),
    .external_source_for_core_0_clock(system_external_source_for_core_0_clock),
    .external_source_for_core_0_reset(system_external_source_for_core_0_reset),
    .halt_from_tile_0(system_halt_from_tile_0),
    .wfi_from_tile_0(system_wfi_from_tile_0),
    .cease_from_tile_0(system_cease_from_tile_0),
    .debug_from_tile_0(system_debug_from_tile_0),
    .psd_test_clock_enable(system_psd_test_clock_enable),
    .resetctrl_hartIsInReset_0(system_resetctrl_hartIsInReset_0),
    .debug_clock(system_debug_clock),
    .debug_reset(system_debug_reset),
    .debug_systemjtag_jtag_TCK(system_debug_systemjtag_jtag_TCK),
    .debug_systemjtag_jtag_TMS(system_debug_systemjtag_jtag_TMS),
    .debug_systemjtag_jtag_TDI(system_debug_systemjtag_jtag_TDI),
    .debug_systemjtag_jtag_TDO_data(system_debug_systemjtag_jtag_TDO_data),
    .debug_systemjtag_jtag_TDO_driven(system_debug_systemjtag_jtag_TDO_driven),
    .debug_systemjtag_reset(system_debug_systemjtag_reset),
    .debug_systemjtag_mfr_id(system_debug_systemjtag_mfr_id),
    .debug_systemjtag_part_number(system_debug_systemjtag_part_number),
    .debug_systemjtag_version(system_debug_systemjtag_version),
    .debug_ndreset(system_debug_ndreset),
    .debug_dmactive(system_debug_dmactive),
    .debug_dmactiveAck(system_debug_dmactiveAck),
    .reset_vector_0(system_reset_vector_0),
    .nmi_0_rnmi(system_nmi_0_rnmi),
    .nmi_0_rnmi_interrupt_vector(system_nmi_0_rnmi_interrupt_vector),
    .nmi_0_rnmi_exception_vector(system_nmi_0_rnmi_exception_vector),
    .rtc_toggle(system_rtc_toggle),
    .global_interrupts(system_global_interrupts),
    .local_interrupts_0(system_local_interrupts_0),
    .sys_port_ahb_0_hmastlock(system_sys_port_ahb_0_hmastlock),
    .sys_port_ahb_0_hready(system_sys_port_ahb_0_hready),
    .sys_port_ahb_0_htrans(system_sys_port_ahb_0_htrans),
    .sys_port_ahb_0_hsize(system_sys_port_ahb_0_hsize),
    .sys_port_ahb_0_hburst(system_sys_port_ahb_0_hburst),
    .sys_port_ahb_0_hwrite(system_sys_port_ahb_0_hwrite),
    .sys_port_ahb_0_hprot(system_sys_port_ahb_0_hprot),
    .sys_port_ahb_0_haddr(system_sys_port_ahb_0_haddr),
    .sys_port_ahb_0_hwdata(system_sys_port_ahb_0_hwdata),
    .sys_port_ahb_0_hresp(system_sys_port_ahb_0_hresp),
    .sys_port_ahb_0_hrdata(system_sys_port_ahb_0_hrdata),
    .periph_port_ahb_0_hmastlock(system_periph_port_ahb_0_hmastlock),
    .periph_port_ahb_0_hready(system_periph_port_ahb_0_hready),
    .periph_port_ahb_0_htrans(system_periph_port_ahb_0_htrans),
    .periph_port_ahb_0_hsize(system_periph_port_ahb_0_hsize),
    .periph_port_ahb_0_hburst(system_periph_port_ahb_0_hburst),
    .periph_port_ahb_0_hwrite(system_periph_port_ahb_0_hwrite),
    .periph_port_ahb_0_hprot(system_periph_port_ahb_0_hprot),
    .periph_port_ahb_0_haddr(system_periph_port_ahb_0_haddr),
    .periph_port_ahb_0_hwdata(system_periph_port_ahb_0_hwdata),
    .periph_port_ahb_0_hresp(system_periph_port_ahb_0_hresp),
    .periph_port_ahb_0_hrdata(system_periph_port_ahb_0_hrdata),
    .front_port_ahb_0_hmastlock(system_front_port_ahb_0_hmastlock),
    .front_port_ahb_0_hsel(system_front_port_ahb_0_hsel),
    .front_port_ahb_0_hready(system_front_port_ahb_0_hready),
    .front_port_ahb_0_hreadyout(system_front_port_ahb_0_hreadyout),
    .front_port_ahb_0_htrans(system_front_port_ahb_0_htrans),
    .front_port_ahb_0_hsize(system_front_port_ahb_0_hsize),
    .front_port_ahb_0_hburst(system_front_port_ahb_0_hburst),
    .front_port_ahb_0_hwrite(system_front_port_ahb_0_hwrite),
    .front_port_ahb_0_hprot(system_front_port_ahb_0_hprot),
    .front_port_ahb_0_haddr(system_front_port_ahb_0_haddr),
    .front_port_ahb_0_hwdata(system_front_port_ahb_0_hwdata),
    .front_port_ahb_0_hresp(system_front_port_ahb_0_hresp),
    .front_port_ahb_0_hrdata(system_front_port_ahb_0_hrdata)
  );
  Pow2ClockDivider func_clock (
    .clock(func_clock_clock),
    .io_clock_out(func_clock_io_clock_out)
  );
  Pow2ClockDivider_1 system_clock_divider (
    .clock(system_clock_divider_clock),
    .io_clock_out(system_clock_divider_io_clock_out)
  );
  ClockSkew #(.DELAY_RTL(0.0), .DELAY_GL(0.0)) core_clocks_skew (
    .clkin(core_clocks_skew_clkin),
    .clkout(core_clocks_skew_clkout)
  );
  system_clock_en dpiClockGate (
    .clock_in(dpiClockGate_clock_in),
    .clock_out(dpiClockGate_clock_out)
  );
  plusarg_reader #(.FORMAT("global_reset_vector=%d"), .DEFAULT(536870912), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  c_core_reset_driver c_core_reset_driver (
    .clock(c_core_reset_driver_clock),
    .out(c_core_reset_driver_out)
  );
  SiFive_DebugCompatibility_DebugCompatibility debug_compatibility (
    .clock(debug_compatibility_clock),
    .debug_outer_reset(debug_compatibility_debug_outer_reset),
    .core_resets_in_0(debug_compatibility_core_resets_in_0),
    .debug_clock(debug_compatibility_debug_clock),
    .debug_reset(debug_compatibility_debug_reset),
    .debug_dmactive(debug_compatibility_debug_dmactive),
    .debug_dmactiveAck(debug_compatibility_debug_dmactiveAck),
    .debug_resetctrl_hartIsInReset_0(debug_compatibility_debug_resetctrl_hartIsInReset_0),
    .core_resets_out_0(debug_compatibility_core_resets_out_0)
  );
  plusarg_reader #(.FORMAT("core_reset_delay=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_1 (
    .out(plusarg_reader_1_out)
  );
  CountAndDriver delayed_reset_count_and_driver (
    .clock(delayed_reset_count_and_driver_clock),
    .reset(delayed_reset_count_and_driver_reset),
    .io_default_value(delayed_reset_count_and_driver_io_default_value),
    .io_count(delayed_reset_count_and_driver_io_count),
    .io_driven_value(delayed_reset_count_and_driver_io_driven_value)
  );
  DataTap_10 coreTraces_DataTap_10 (
    ._0_clock(coreTraces_DataTap_10__0_clock),
    ._0_reset(coreTraces_DataTap_10__0_reset),
    ._0_excpt(coreTraces_DataTap_10__0_excpt),
    ._0_priv_mode(coreTraces_DataTap_10__0_priv_mode),
    ._0_hartid(coreTraces_DataTap_10__0_hartid),
    ._0_timer(coreTraces_DataTap_10__0_timer),
    ._0_valid(coreTraces_DataTap_10__0_valid),
    ._0_pc(coreTraces_DataTap_10__0_pc),
    ._0_wrdst(coreTraces_DataTap_10__0_wrdst),
    ._0_wrdata(coreTraces_DataTap_10__0_wrdata),
    ._0_wrenx(coreTraces_DataTap_10__0_wrenx),
    ._0_wrenf(coreTraces_DataTap_10__0_wrenf),
    ._0_rd0src(coreTraces_DataTap_10__0_rd0src),
    ._0_rd0val(coreTraces_DataTap_10__0_rd0val),
    ._0_rd1src(coreTraces_DataTap_10__0_rd1src),
    ._0_rd1val(coreTraces_DataTap_10__0_rd1val),
    ._0_inst(coreTraces_DataTap_10__0_inst)
  );
  DataTap_1_0 csrTraces_DataTap_1 (
    ._9(csrTraces_DataTap_1__9),
    ._8(csrTraces_DataTap_1__8),
    ._7(csrTraces_DataTap_1__7),
    ._6(csrTraces_DataTap_1__6),
    ._5(csrTraces_DataTap_1__5),
    ._4(csrTraces_DataTap_1__4),
    ._3(csrTraces_DataTap_1__3),
    ._2(csrTraces_DataTap_1__2),
    ._1(csrTraces_DataTap_1__1),
    ._0(csrTraces_DataTap_1__0)
  );
  AHBPortRAMSlave testRAM (
    .clock(testRAM_clock),
    .reset(testRAM_reset),
    .io_ahb_0_hmastlock(testRAM_io_ahb_0_hmastlock),
    .io_ahb_0_hready(testRAM_io_ahb_0_hready),
    .io_ahb_0_htrans(testRAM_io_ahb_0_htrans),
    .io_ahb_0_hsize(testRAM_io_ahb_0_hsize),
    .io_ahb_0_hburst(testRAM_io_ahb_0_hburst),
    .io_ahb_0_hwrite(testRAM_io_ahb_0_hwrite),
    .io_ahb_0_hprot(testRAM_io_ahb_0_hprot),
    .io_ahb_0_haddr(testRAM_io_ahb_0_haddr),
    .io_ahb_0_hwdata(testRAM_io_ahb_0_hwdata),
    .io_ahb_0_hresp(testRAM_io_ahb_0_hresp),
    .io_ahb_0_hrdata(testRAM_io_ahb_0_hrdata)
  );
  XSquasher #(.WIDTH(32)) system_periph_port_ahb_0_hrdata_xs (
    .valid(system_periph_port_ahb_0_hrdata_xs_valid),
    .inp(system_periph_port_ahb_0_hrdata_xs_inp),
    .outp(system_periph_port_ahb_0_hrdata_xs_outp)
  );
  XSquasher #(.WIDTH(1)) system_periph_port_ahb_0_hresp_xs (
    .valid(system_periph_port_ahb_0_hresp_xs_valid),
    .inp(system_periph_port_ahb_0_hresp_xs_inp),
    .outp(system_periph_port_ahb_0_hresp_xs_outp)
  );
  AHBPortRAMSlave_1 testRAM_1 (
    .clock(testRAM_1_clock),
    .reset(testRAM_1_reset),
    .io_ahb_0_hmastlock(testRAM_1_io_ahb_0_hmastlock),
    .io_ahb_0_hready(testRAM_1_io_ahb_0_hready),
    .io_ahb_0_htrans(testRAM_1_io_ahb_0_htrans),
    .io_ahb_0_hsize(testRAM_1_io_ahb_0_hsize),
    .io_ahb_0_hburst(testRAM_1_io_ahb_0_hburst),
    .io_ahb_0_hwrite(testRAM_1_io_ahb_0_hwrite),
    .io_ahb_0_hprot(testRAM_1_io_ahb_0_hprot),
    .io_ahb_0_haddr(testRAM_1_io_ahb_0_haddr),
    .io_ahb_0_hwdata(testRAM_1_io_ahb_0_hwdata),
    .io_ahb_0_hresp(testRAM_1_io_ahb_0_hresp),
    .io_ahb_0_hrdata(testRAM_1_io_ahb_0_hrdata)
  );
  XSquasher #(.WIDTH(32)) system_sys_port_ahb_0_hrdata_xs (
    .valid(system_sys_port_ahb_0_hrdata_xs_valid),
    .inp(system_sys_port_ahb_0_hrdata_xs_inp),
    .outp(system_sys_port_ahb_0_hrdata_xs_outp)
  );
  XSquasher #(.WIDTH(1)) system_sys_port_ahb_0_hresp_xs (
    .valid(system_sys_port_ahb_0_hresp_xs_valid),
    .inp(system_sys_port_ahb_0_hresp_xs_inp),
    .outp(system_sys_port_ahb_0_hresp_xs_outp)
  );
  WfiChecker #(.PCWIDTH(32)) wfichecker (
    .reset(wfichecker_reset),
    .clock(wfichecker_clock),
    .wfi(wfichecker_wfi),
    .csr_hartid(wfichecker_csr_hartid),
    .excpt(wfichecker_excpt),
    .bus_err_int(wfichecker_bus_err_int),
    .debug_int(wfichecker_debug_int),
    .clint_int(wfichecker_clint_int),
    .allow_wfi(wfichecker_allow_wfi),
    .debug(wfichecker_debug),
    .singleStep(wfichecker_singleStep),
    .reg_mie(wfichecker_reg_mie),
    .reg_mip(wfichecker_reg_mip),
    .inst_hartid_0(wfichecker_inst_hartid_0),
    .inst_vld_0(wfichecker_inst_vld_0),
    .pc_0(wfichecker_pc_0),
    .inst_0(wfichecker_inst_0)
  );
  core_monitor core_monitor (
    .m_0_clock(core_monitor_m_0_clock),
    .m_0_reset(core_monitor_m_0_reset),
    .m_0_excpt(core_monitor_m_0_excpt),
    .m_0_priv_mode(core_monitor_m_0_priv_mode),
    .m_0_hartid(core_monitor_m_0_hartid),
    .m_0_timer(core_monitor_m_0_timer),
    .m_0_valid(core_monitor_m_0_valid),
    .m_0_pc(core_monitor_m_0_pc),
    .m_0_wrdst(core_monitor_m_0_wrdst),
    .m_0_wrdata(core_monitor_m_0_wrdata),
    .m_0_wrenx(core_monitor_m_0_wrenx),
    .m_0_wrenf(core_monitor_m_0_wrenf),
    .m_0_rd0src(core_monitor_m_0_rd0src),
    .m_0_rd0val(core_monitor_m_0_rd0val),
    .m_0_rd1src(core_monitor_m_0_rd1src),
    .m_0_rd1val(core_monitor_m_0_rd1val),
    .m_0_inst(core_monitor_m_0_inst)
  );
  DPITestbenchHooks dpitbh (
    .clock(dpitbh_clock),
    .reset(dpitbh_reset)
  );
  plusarg_reader #(.FORMAT("drive_global_interrupt_type=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_2 (
    .out(plusarg_reader_2_out)
  );
  GlobalIntDriver dpi_driver (
    .clock(dpi_driver_clock),
    .reset(dpi_driver_reset),
    .interrupts(dpi_driver_interrupts)
  );
  plusarg_reader #(.FORMAT("drive_local_interrupt_type=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader_3 (
    .out(plusarg_reader_3_out)
  );
  NullInterruptDriver #(.ID(0), .WIDTH(32)) dpi_drivers_0 (
    .clock(dpi_drivers_0_clock),
    .reset(dpi_drivers_0_reset),
    .interrupts(dpi_drivers_0_interrupts)
  );
  assign io_success = 1'h1;
  assign system_clock = dpiClockGate_clock_out;
  assign system_reset = reset | system_debug_ndreset;
  assign system_external_source_for_core_0_clock = core_clocks_skew_clkout;
  assign system_external_source_for_core_0_reset = delayed_reset_count_and_driver_io_driven_value;
  assign system_psd_test_clock_enable = 1'h0;
  assign system_resetctrl_hartIsInReset_0 = debug_compatibility_debug_resetctrl_hartIsInReset_0;
  assign system_debug_clock = debug_compatibility_debug_clock;
  assign system_debug_reset = debug_compatibility_debug_reset;
  assign system_debug_systemjtag_jtag_TCK = 1'h1;
  assign system_debug_systemjtag_jtag_TMS = 1'h1;
  assign system_debug_systemjtag_jtag_TDI = 1'h1;
  assign system_debug_systemjtag_reset = reset;
  assign system_debug_systemjtag_mfr_id = 11'h0;
  assign system_debug_systemjtag_part_number = 16'h0;
  assign system_debug_systemjtag_version = 4'h0;
  assign system_debug_dmactiveAck = debug_compatibility_debug_dmactiveAck;
  assign system_reset_vector_0 = plusarg_reader_out;
  assign system_nmi_0_rnmi = 1'h0;
  assign system_nmi_0_rnmi_interrupt_vector = 32'h0;
  assign system_nmi_0_rnmi_exception_vector = 32'h0;
  assign system_rtc_toggle = toggle;
  assign system_global_interrupts = _GEN_523[126:0];
  assign system_local_interrupts_0 = _GEN_597[15:0];
  assign system_sys_port_ahb_0_hready = testRAM_1_io_ahb_0_hready;
  assign system_sys_port_ahb_0_hresp = system_sys_port_ahb_0_hresp_xs_outp;
  assign system_sys_port_ahb_0_hrdata = system_sys_port_ahb_0_hrdata_xs_outp;
  assign system_periph_port_ahb_0_hready = testRAM_io_ahb_0_hready;
  assign system_periph_port_ahb_0_hresp = system_periph_port_ahb_0_hresp_xs_outp;
  assign system_periph_port_ahb_0_hrdata = system_periph_port_ahb_0_hrdata_xs_outp;
  assign system_front_port_ahb_0_hmastlock = 1'h0;
  assign system_front_port_ahb_0_hsel = 1'h0;
  assign system_front_port_ahb_0_hready = 1'h0;
  assign system_front_port_ahb_0_htrans = 2'h0;
  assign system_front_port_ahb_0_hsize = 3'h0;
  assign system_front_port_ahb_0_hburst = 3'h0;
  assign system_front_port_ahb_0_hwrite = 1'h0;
  assign system_front_port_ahb_0_hprot = 4'h3;
  assign system_front_port_ahb_0_haddr = 32'h0;
  assign system_front_port_ahb_0_hwdata = 32'h0;
  assign func_clock_clock = clock;
  assign system_clock_divider_clock = func_clock_io_clock_out;
  assign core_clocks_skew_clkin = func_clock_io_clock_out;
  assign dpiClockGate_clock_in = system_clock_divider_io_clock_out;
  assign c_core_reset_driver_clock = clock;
  assign debug_compatibility_clock = system_clock;
  assign debug_compatibility_debug_outer_reset = system_debug_systemjtag_reset;
  assign debug_compatibility_core_resets_in_0 = reset | ndm_reset | c_core_reset_driver_out | system_reset;
  assign debug_compatibility_debug_dmactive = system_debug_dmactive;
  assign delayed_reset_count_and_driver_clock = clock;
  assign delayed_reset_count_and_driver_reset = reset;
  assign delayed_reset_count_and_driver_io_default_value = debug_compatibility_core_resets_out_0;
  assign delayed_reset_count_and_driver_io_count = plusarg_reader_1_out[15:0];
  assign testRAM_clock = dpiClockGate_clock_out;
  assign testRAM_reset = system_reset | reset;
  assign testRAM_io_ahb_0_hmastlock = system_periph_port_ahb_0_hmastlock;
  assign testRAM_io_ahb_0_htrans = system_periph_port_ahb_0_htrans;
  assign testRAM_io_ahb_0_hsize = system_periph_port_ahb_0_hsize;
  assign testRAM_io_ahb_0_hburst = system_periph_port_ahb_0_hburst;
  assign testRAM_io_ahb_0_hwrite = system_periph_port_ahb_0_hwrite;
  assign testRAM_io_ahb_0_hprot = system_periph_port_ahb_0_hprot;
  assign testRAM_io_ahb_0_haddr = system_periph_port_ahb_0_haddr;
  assign testRAM_io_ahb_0_hwdata = system_periph_port_ahb_0_hwdata;
  assign system_periph_port_ahb_0_hrdata_xs_valid = system_periph_port_ahb_0_hrdata_xs_io_valid_r & ~
    system_periph_port_ahb_0_hrdata_xs_io_valid_r_1 & testRAM_io_ahb_0_hready & ~testRAM_io_ahb_0_hresp;
  assign system_periph_port_ahb_0_hrdata_xs_inp = testRAM_io_ahb_0_hrdata;
  assign system_periph_port_ahb_0_hresp_xs_valid = system_periph_port_ahb_0_hresp_xs_io_valid_r;
  assign system_periph_port_ahb_0_hresp_xs_inp = testRAM_io_ahb_0_hresp;
  assign testRAM_1_clock = dpiClockGate_clock_out;
  assign testRAM_1_reset = system_reset | reset;
  assign testRAM_1_io_ahb_0_hmastlock = system_sys_port_ahb_0_hmastlock;
  assign testRAM_1_io_ahb_0_htrans = system_sys_port_ahb_0_htrans;
  assign testRAM_1_io_ahb_0_hsize = system_sys_port_ahb_0_hsize;
  assign testRAM_1_io_ahb_0_hburst = system_sys_port_ahb_0_hburst;
  assign testRAM_1_io_ahb_0_hwrite = system_sys_port_ahb_0_hwrite;
  assign testRAM_1_io_ahb_0_hprot = system_sys_port_ahb_0_hprot;
  assign testRAM_1_io_ahb_0_haddr = system_sys_port_ahb_0_haddr;
  assign testRAM_1_io_ahb_0_hwdata = system_sys_port_ahb_0_hwdata;
  assign system_sys_port_ahb_0_hrdata_xs_valid = system_sys_port_ahb_0_hrdata_xs_io_valid_r & ~
    system_sys_port_ahb_0_hrdata_xs_io_valid_r_1 & testRAM_1_io_ahb_0_hready & ~testRAM_1_io_ahb_0_hresp;
  assign system_sys_port_ahb_0_hrdata_xs_inp = testRAM_1_io_ahb_0_hrdata;
  assign system_sys_port_ahb_0_hresp_xs_valid = system_sys_port_ahb_0_hresp_xs_io_valid_r;
  assign system_sys_port_ahb_0_hresp_xs_inp = testRAM_1_io_ahb_0_hresp;
  assign wfichecker_reset = reset;
  assign wfichecker_clock = clock;
  assign wfichecker_wfi = system_wfi_from_tile_0;
  assign wfichecker_csr_hartid = {{31'd0}, csrTraces_hartid};
  assign wfichecker_excpt = csrTraces_DataTap_1__6;
  assign wfichecker_bus_err_int = 1'h0;
  assign wfichecker_debug_int = csrTraces_DataTap_1__7;
  assign wfichecker_clint_int = 1'h0;
  assign wfichecker_allow_wfi = 1'h1;
  assign wfichecker_debug = csrTraces_DataTap_1__8;
  assign wfichecker_singleStep = csrTraces_DataTap_1__9;
  assign wfichecker_reg_mie = csrTraces_DataTap_1__1;
  assign wfichecker_reg_mip = csrTraces_DataTap_1__2;
  assign wfichecker_inst_hartid_0 = coreTraces_DataTap_10__0_hartid;
  assign wfichecker_inst_vld_0 = coreTraces_DataTap_10__0_valid;
  assign wfichecker_pc_0 = coreTraces_DataTap_10__0_pc;
  assign wfichecker_inst_0 = coreTraces_DataTap_10__0_inst;
  assign core_monitor_m_0_clock = coreTraces_DataTap_10__0_clock;
  assign core_monitor_m_0_reset = coreTraces_DataTap_10__0_reset;
  assign core_monitor_m_0_excpt = coreTraces_DataTap_10__0_excpt;
  assign core_monitor_m_0_priv_mode = coreTraces_DataTap_10__0_priv_mode;
  assign core_monitor_m_0_hartid = coreTraces_DataTap_10__0_hartid;
  assign core_monitor_m_0_timer = coreTraces_DataTap_10__0_timer;
  assign core_monitor_m_0_valid = coreTraces_DataTap_10__0_valid;
  assign core_monitor_m_0_pc = coreTraces_DataTap_10__0_pc;
  assign core_monitor_m_0_wrdst = coreTraces_DataTap_10__0_wrdst;
  assign core_monitor_m_0_wrdata = coreTraces_DataTap_10__0_wrdata;
  assign core_monitor_m_0_wrenx = coreTraces_DataTap_10__0_wrenx;
  assign core_monitor_m_0_wrenf = coreTraces_DataTap_10__0_wrenf;
  assign core_monitor_m_0_rd0src = coreTraces_DataTap_10__0_rd0src;
  assign core_monitor_m_0_rd0val = coreTraces_DataTap_10__0_rd0val;
  assign core_monitor_m_0_rd1src = coreTraces_DataTap_10__0_rd1src;
  assign core_monitor_m_0_rd1val = coreTraces_DataTap_10__0_rd1val;
  assign core_monitor_m_0_inst = coreTraces_DataTap_10__0_inst;
  assign dpitbh_clock = 1'h0;
  assign dpitbh_reset = 1'h0;
  assign dpi_driver_clock = 1'h0;
  assign dpi_driver_reset = 1'h0;
  assign dpi_drivers_0_clock = 1'h0;
  assign dpi_drivers_0_reset = 1'h0;
  always @(posedge dpiClockGate_clock_out) begin
    if (reset) begin
      count <= 5'h0;
    end else begin
      count <= _count_T_1;
    end
    if (reset) begin
      toggle <= 1'h0;
    end else if (count == 5'h0) begin
      toggle <= ~toggle;
    end
    if (ram_reset) begin
      system_periph_port_ahb_0_hrdata_xs_io_valid_r <= 1'h0;
    end else if (testRAM_io_ahb_0_hready) begin
      system_periph_port_ahb_0_hrdata_xs_io_valid_r <= testRAM_io_ahb_0_htrans == 2'h2 | testRAM_io_ahb_0_htrans == 2'h3
        ;
    end
    if (ram_reset) begin
      system_periph_port_ahb_0_hrdata_xs_io_valid_r_1 <= 1'h0;
    end else if (testRAM_io_ahb_0_hready) begin
      system_periph_port_ahb_0_hrdata_xs_io_valid_r_1 <= testRAM_io_ahb_0_hwrite & (testRAM_io_ahb_0_htrans == 2'h2 |
        testRAM_io_ahb_0_htrans == 2'h3);
    end
    if (ram_reset) begin
      system_periph_port_ahb_0_hresp_xs_io_valid_r <= 1'h0;
    end else if (testRAM_io_ahb_0_hready) begin
      system_periph_port_ahb_0_hresp_xs_io_valid_r <= testRAM_io_ahb_0_htrans == 2'h2 | testRAM_io_ahb_0_htrans == 2'h3;
    end
    if (ram_reset) begin
      system_sys_port_ahb_0_hrdata_xs_io_valid_r <= 1'h0;
    end else if (testRAM_1_io_ahb_0_hready) begin
      system_sys_port_ahb_0_hrdata_xs_io_valid_r <= testRAM_1_io_ahb_0_htrans == 2'h2 | testRAM_1_io_ahb_0_htrans == 2'h3
        ;
    end
    if (ram_reset) begin
      system_sys_port_ahb_0_hrdata_xs_io_valid_r_1 <= 1'h0;
    end else if (testRAM_1_io_ahb_0_hready) begin
      system_sys_port_ahb_0_hrdata_xs_io_valid_r_1 <= testRAM_1_io_ahb_0_hwrite & (testRAM_1_io_ahb_0_htrans == 2'h2 |
        testRAM_1_io_ahb_0_htrans == 2'h3);
    end
    if (ram_reset) begin
      system_sys_port_ahb_0_hresp_xs_io_valid_r <= 1'h0;
    end else if (testRAM_1_io_ahb_0_hready) begin
      system_sys_port_ahb_0_hresp_xs_io_valid_r <= testRAM_1_io_ahb_0_htrans == 2'h2 | testRAM_1_io_ahb_0_htrans == 2'h3
        ;
    end
  end
  always @(posedge clock) begin
    if (reset) begin
      tick_value <= 7'h0;
    end else if (tick) begin
      tick_value <= 7'h0;
    end else begin
      tick_value <= _tick_value_T_1;
    end
    if (reset) begin
      system_global_interrupts_value <= 7'h0;
    end else if (tick) begin
      if (system_global_interrupts_wrap_wrap) begin
        system_global_interrupts_value <= 7'h0;
      end else begin
        system_global_interrupts_value <= _system_global_interrupts_wrap_value_T_1;
      end
    end
    if (tickers_x3_lfsrReg == 16'h0) begin
      tickers_x3_lfsrReg <= 16'h1;
    end else begin
      tickers_x3_lfsrReg <= _tickers_x3_lfsrReg_T_6;
    end
    if (tickers_x3_lfsrReg_1 == 16'h0) begin
      tickers_x3_lfsrReg_1 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_1 <= _tickers_x3_lfsrReg_T_13;
    end
    if (tickers_x3_lfsrReg_2 == 16'h0) begin
      tickers_x3_lfsrReg_2 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_2 <= _tickers_x3_lfsrReg_T_20;
    end
    if (tickers_x3_lfsrReg_3 == 16'h0) begin
      tickers_x3_lfsrReg_3 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_3 <= _tickers_x3_lfsrReg_T_27;
    end
    if (tickers_x3_lfsrReg_4 == 16'h0) begin
      tickers_x3_lfsrReg_4 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_4 <= _tickers_x3_lfsrReg_T_34;
    end
    if (tickers_x3_lfsrReg_5 == 16'h0) begin
      tickers_x3_lfsrReg_5 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_5 <= _tickers_x3_lfsrReg_T_41;
    end
    if (tickers_x3_lfsrReg_6 == 16'h0) begin
      tickers_x3_lfsrReg_6 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_6 <= _tickers_x3_lfsrReg_T_48;
    end
    if (tickers_x3_lfsrReg_7 == 16'h0) begin
      tickers_x3_lfsrReg_7 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_7 <= _tickers_x3_lfsrReg_T_55;
    end
    if (tickers_x3_lfsrReg_8 == 16'h0) begin
      tickers_x3_lfsrReg_8 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_8 <= _tickers_x3_lfsrReg_T_62;
    end
    if (tickers_x3_lfsrReg_9 == 16'h0) begin
      tickers_x3_lfsrReg_9 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_9 <= _tickers_x3_lfsrReg_T_69;
    end
    if (tickers_x3_lfsrReg_10 == 16'h0) begin
      tickers_x3_lfsrReg_10 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_10 <= _tickers_x3_lfsrReg_T_76;
    end
    if (tickers_x3_lfsrReg_11 == 16'h0) begin
      tickers_x3_lfsrReg_11 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_11 <= _tickers_x3_lfsrReg_T_83;
    end
    if (tickers_x3_lfsrReg_12 == 16'h0) begin
      tickers_x3_lfsrReg_12 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_12 <= _tickers_x3_lfsrReg_T_90;
    end
    if (tickers_x3_lfsrReg_13 == 16'h0) begin
      tickers_x3_lfsrReg_13 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_13 <= _tickers_x3_lfsrReg_T_97;
    end
    if (tickers_x3_lfsrReg_14 == 16'h0) begin
      tickers_x3_lfsrReg_14 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_14 <= _tickers_x3_lfsrReg_T_104;
    end
    if (tickers_x3_lfsrReg_15 == 16'h0) begin
      tickers_x3_lfsrReg_15 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_15 <= _tickers_x3_lfsrReg_T_111;
    end
    if (tickers_x3_lfsrReg_16 == 16'h0) begin
      tickers_x3_lfsrReg_16 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_16 <= _tickers_x3_lfsrReg_T_118;
    end
    if (tickers_x3_lfsrReg_17 == 16'h0) begin
      tickers_x3_lfsrReg_17 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_17 <= _tickers_x3_lfsrReg_T_125;
    end
    if (tickers_x3_lfsrReg_18 == 16'h0) begin
      tickers_x3_lfsrReg_18 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_18 <= _tickers_x3_lfsrReg_T_132;
    end
    if (tickers_x3_lfsrReg_19 == 16'h0) begin
      tickers_x3_lfsrReg_19 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_19 <= _tickers_x3_lfsrReg_T_139;
    end
    if (tickers_x3_lfsrReg_20 == 16'h0) begin
      tickers_x3_lfsrReg_20 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_20 <= _tickers_x3_lfsrReg_T_146;
    end
    if (tickers_x3_lfsrReg_21 == 16'h0) begin
      tickers_x3_lfsrReg_21 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_21 <= _tickers_x3_lfsrReg_T_153;
    end
    if (tickers_x3_lfsrReg_22 == 16'h0) begin
      tickers_x3_lfsrReg_22 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_22 <= _tickers_x3_lfsrReg_T_160;
    end
    if (tickers_x3_lfsrReg_23 == 16'h0) begin
      tickers_x3_lfsrReg_23 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_23 <= _tickers_x3_lfsrReg_T_167;
    end
    if (tickers_x3_lfsrReg_24 == 16'h0) begin
      tickers_x3_lfsrReg_24 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_24 <= _tickers_x3_lfsrReg_T_174;
    end
    if (tickers_x3_lfsrReg_25 == 16'h0) begin
      tickers_x3_lfsrReg_25 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_25 <= _tickers_x3_lfsrReg_T_181;
    end
    if (tickers_x3_lfsrReg_26 == 16'h0) begin
      tickers_x3_lfsrReg_26 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_26 <= _tickers_x3_lfsrReg_T_188;
    end
    if (tickers_x3_lfsrReg_27 == 16'h0) begin
      tickers_x3_lfsrReg_27 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_27 <= _tickers_x3_lfsrReg_T_195;
    end
    if (tickers_x3_lfsrReg_28 == 16'h0) begin
      tickers_x3_lfsrReg_28 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_28 <= _tickers_x3_lfsrReg_T_202;
    end
    if (tickers_x3_lfsrReg_29 == 16'h0) begin
      tickers_x3_lfsrReg_29 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_29 <= _tickers_x3_lfsrReg_T_209;
    end
    if (tickers_x3_lfsrReg_30 == 16'h0) begin
      tickers_x3_lfsrReg_30 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_30 <= _tickers_x3_lfsrReg_T_216;
    end
    if (tickers_x3_lfsrReg_31 == 16'h0) begin
      tickers_x3_lfsrReg_31 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_31 <= _tickers_x3_lfsrReg_T_223;
    end
    if (tickers_x3_lfsrReg_32 == 16'h0) begin
      tickers_x3_lfsrReg_32 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_32 <= _tickers_x3_lfsrReg_T_230;
    end
    if (tickers_x3_lfsrReg_33 == 16'h0) begin
      tickers_x3_lfsrReg_33 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_33 <= _tickers_x3_lfsrReg_T_237;
    end
    if (tickers_x3_lfsrReg_34 == 16'h0) begin
      tickers_x3_lfsrReg_34 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_34 <= _tickers_x3_lfsrReg_T_244;
    end
    if (tickers_x3_lfsrReg_35 == 16'h0) begin
      tickers_x3_lfsrReg_35 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_35 <= _tickers_x3_lfsrReg_T_251;
    end
    if (tickers_x3_lfsrReg_36 == 16'h0) begin
      tickers_x3_lfsrReg_36 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_36 <= _tickers_x3_lfsrReg_T_258;
    end
    if (tickers_x3_lfsrReg_37 == 16'h0) begin
      tickers_x3_lfsrReg_37 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_37 <= _tickers_x3_lfsrReg_T_265;
    end
    if (tickers_x3_lfsrReg_38 == 16'h0) begin
      tickers_x3_lfsrReg_38 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_38 <= _tickers_x3_lfsrReg_T_272;
    end
    if (tickers_x3_lfsrReg_39 == 16'h0) begin
      tickers_x3_lfsrReg_39 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_39 <= _tickers_x3_lfsrReg_T_279;
    end
    if (tickers_x3_lfsrReg_40 == 16'h0) begin
      tickers_x3_lfsrReg_40 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_40 <= _tickers_x3_lfsrReg_T_286;
    end
    if (tickers_x3_lfsrReg_41 == 16'h0) begin
      tickers_x3_lfsrReg_41 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_41 <= _tickers_x3_lfsrReg_T_293;
    end
    if (tickers_x3_lfsrReg_42 == 16'h0) begin
      tickers_x3_lfsrReg_42 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_42 <= _tickers_x3_lfsrReg_T_300;
    end
    if (tickers_x3_lfsrReg_43 == 16'h0) begin
      tickers_x3_lfsrReg_43 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_43 <= _tickers_x3_lfsrReg_T_307;
    end
    if (tickers_x3_lfsrReg_44 == 16'h0) begin
      tickers_x3_lfsrReg_44 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_44 <= _tickers_x3_lfsrReg_T_314;
    end
    if (tickers_x3_lfsrReg_45 == 16'h0) begin
      tickers_x3_lfsrReg_45 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_45 <= _tickers_x3_lfsrReg_T_321;
    end
    if (tickers_x3_lfsrReg_46 == 16'h0) begin
      tickers_x3_lfsrReg_46 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_46 <= _tickers_x3_lfsrReg_T_328;
    end
    if (tickers_x3_lfsrReg_47 == 16'h0) begin
      tickers_x3_lfsrReg_47 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_47 <= _tickers_x3_lfsrReg_T_335;
    end
    if (tickers_x3_lfsrReg_48 == 16'h0) begin
      tickers_x3_lfsrReg_48 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_48 <= _tickers_x3_lfsrReg_T_342;
    end
    if (tickers_x3_lfsrReg_49 == 16'h0) begin
      tickers_x3_lfsrReg_49 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_49 <= _tickers_x3_lfsrReg_T_349;
    end
    if (tickers_x3_lfsrReg_50 == 16'h0) begin
      tickers_x3_lfsrReg_50 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_50 <= _tickers_x3_lfsrReg_T_356;
    end
    if (tickers_x3_lfsrReg_51 == 16'h0) begin
      tickers_x3_lfsrReg_51 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_51 <= _tickers_x3_lfsrReg_T_363;
    end
    if (tickers_x3_lfsrReg_52 == 16'h0) begin
      tickers_x3_lfsrReg_52 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_52 <= _tickers_x3_lfsrReg_T_370;
    end
    if (tickers_x3_lfsrReg_53 == 16'h0) begin
      tickers_x3_lfsrReg_53 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_53 <= _tickers_x3_lfsrReg_T_377;
    end
    if (tickers_x3_lfsrReg_54 == 16'h0) begin
      tickers_x3_lfsrReg_54 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_54 <= _tickers_x3_lfsrReg_T_384;
    end
    if (tickers_x3_lfsrReg_55 == 16'h0) begin
      tickers_x3_lfsrReg_55 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_55 <= _tickers_x3_lfsrReg_T_391;
    end
    if (tickers_x3_lfsrReg_56 == 16'h0) begin
      tickers_x3_lfsrReg_56 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_56 <= _tickers_x3_lfsrReg_T_398;
    end
    if (tickers_x3_lfsrReg_57 == 16'h0) begin
      tickers_x3_lfsrReg_57 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_57 <= _tickers_x3_lfsrReg_T_405;
    end
    if (tickers_x3_lfsrReg_58 == 16'h0) begin
      tickers_x3_lfsrReg_58 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_58 <= _tickers_x3_lfsrReg_T_412;
    end
    if (tickers_x3_lfsrReg_59 == 16'h0) begin
      tickers_x3_lfsrReg_59 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_59 <= _tickers_x3_lfsrReg_T_419;
    end
    if (tickers_x3_lfsrReg_60 == 16'h0) begin
      tickers_x3_lfsrReg_60 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_60 <= _tickers_x3_lfsrReg_T_426;
    end
    if (tickers_x3_lfsrReg_61 == 16'h0) begin
      tickers_x3_lfsrReg_61 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_61 <= _tickers_x3_lfsrReg_T_433;
    end
    if (tickers_x3_lfsrReg_62 == 16'h0) begin
      tickers_x3_lfsrReg_62 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_62 <= _tickers_x3_lfsrReg_T_440;
    end
    if (tickers_x3_lfsrReg_63 == 16'h0) begin
      tickers_x3_lfsrReg_63 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_63 <= _tickers_x3_lfsrReg_T_447;
    end
    if (tickers_x3_lfsrReg_64 == 16'h0) begin
      tickers_x3_lfsrReg_64 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_64 <= _tickers_x3_lfsrReg_T_454;
    end
    if (tickers_x3_lfsrReg_65 == 16'h0) begin
      tickers_x3_lfsrReg_65 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_65 <= _tickers_x3_lfsrReg_T_461;
    end
    if (tickers_x3_lfsrReg_66 == 16'h0) begin
      tickers_x3_lfsrReg_66 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_66 <= _tickers_x3_lfsrReg_T_468;
    end
    if (tickers_x3_lfsrReg_67 == 16'h0) begin
      tickers_x3_lfsrReg_67 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_67 <= _tickers_x3_lfsrReg_T_475;
    end
    if (tickers_x3_lfsrReg_68 == 16'h0) begin
      tickers_x3_lfsrReg_68 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_68 <= _tickers_x3_lfsrReg_T_482;
    end
    if (tickers_x3_lfsrReg_69 == 16'h0) begin
      tickers_x3_lfsrReg_69 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_69 <= _tickers_x3_lfsrReg_T_489;
    end
    if (tickers_x3_lfsrReg_70 == 16'h0) begin
      tickers_x3_lfsrReg_70 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_70 <= _tickers_x3_lfsrReg_T_496;
    end
    if (tickers_x3_lfsrReg_71 == 16'h0) begin
      tickers_x3_lfsrReg_71 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_71 <= _tickers_x3_lfsrReg_T_503;
    end
    if (tickers_x3_lfsrReg_72 == 16'h0) begin
      tickers_x3_lfsrReg_72 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_72 <= _tickers_x3_lfsrReg_T_510;
    end
    if (tickers_x3_lfsrReg_73 == 16'h0) begin
      tickers_x3_lfsrReg_73 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_73 <= _tickers_x3_lfsrReg_T_517;
    end
    if (tickers_x3_lfsrReg_74 == 16'h0) begin
      tickers_x3_lfsrReg_74 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_74 <= _tickers_x3_lfsrReg_T_524;
    end
    if (tickers_x3_lfsrReg_75 == 16'h0) begin
      tickers_x3_lfsrReg_75 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_75 <= _tickers_x3_lfsrReg_T_531;
    end
    if (tickers_x3_lfsrReg_76 == 16'h0) begin
      tickers_x3_lfsrReg_76 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_76 <= _tickers_x3_lfsrReg_T_538;
    end
    if (tickers_x3_lfsrReg_77 == 16'h0) begin
      tickers_x3_lfsrReg_77 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_77 <= _tickers_x3_lfsrReg_T_545;
    end
    if (tickers_x3_lfsrReg_78 == 16'h0) begin
      tickers_x3_lfsrReg_78 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_78 <= _tickers_x3_lfsrReg_T_552;
    end
    if (tickers_x3_lfsrReg_79 == 16'h0) begin
      tickers_x3_lfsrReg_79 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_79 <= _tickers_x3_lfsrReg_T_559;
    end
    if (tickers_x3_lfsrReg_80 == 16'h0) begin
      tickers_x3_lfsrReg_80 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_80 <= _tickers_x3_lfsrReg_T_566;
    end
    if (tickers_x3_lfsrReg_81 == 16'h0) begin
      tickers_x3_lfsrReg_81 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_81 <= _tickers_x3_lfsrReg_T_573;
    end
    if (tickers_x3_lfsrReg_82 == 16'h0) begin
      tickers_x3_lfsrReg_82 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_82 <= _tickers_x3_lfsrReg_T_580;
    end
    if (tickers_x3_lfsrReg_83 == 16'h0) begin
      tickers_x3_lfsrReg_83 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_83 <= _tickers_x3_lfsrReg_T_587;
    end
    if (tickers_x3_lfsrReg_84 == 16'h0) begin
      tickers_x3_lfsrReg_84 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_84 <= _tickers_x3_lfsrReg_T_594;
    end
    if (tickers_x3_lfsrReg_85 == 16'h0) begin
      tickers_x3_lfsrReg_85 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_85 <= _tickers_x3_lfsrReg_T_601;
    end
    if (tickers_x3_lfsrReg_86 == 16'h0) begin
      tickers_x3_lfsrReg_86 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_86 <= _tickers_x3_lfsrReg_T_608;
    end
    if (tickers_x3_lfsrReg_87 == 16'h0) begin
      tickers_x3_lfsrReg_87 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_87 <= _tickers_x3_lfsrReg_T_615;
    end
    if (tickers_x3_lfsrReg_88 == 16'h0) begin
      tickers_x3_lfsrReg_88 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_88 <= _tickers_x3_lfsrReg_T_622;
    end
    if (tickers_x3_lfsrReg_89 == 16'h0) begin
      tickers_x3_lfsrReg_89 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_89 <= _tickers_x3_lfsrReg_T_629;
    end
    if (tickers_x3_lfsrReg_90 == 16'h0) begin
      tickers_x3_lfsrReg_90 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_90 <= _tickers_x3_lfsrReg_T_636;
    end
    if (tickers_x3_lfsrReg_91 == 16'h0) begin
      tickers_x3_lfsrReg_91 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_91 <= _tickers_x3_lfsrReg_T_643;
    end
    if (tickers_x3_lfsrReg_92 == 16'h0) begin
      tickers_x3_lfsrReg_92 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_92 <= _tickers_x3_lfsrReg_T_650;
    end
    if (tickers_x3_lfsrReg_93 == 16'h0) begin
      tickers_x3_lfsrReg_93 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_93 <= _tickers_x3_lfsrReg_T_657;
    end
    if (tickers_x3_lfsrReg_94 == 16'h0) begin
      tickers_x3_lfsrReg_94 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_94 <= _tickers_x3_lfsrReg_T_664;
    end
    if (tickers_x3_lfsrReg_95 == 16'h0) begin
      tickers_x3_lfsrReg_95 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_95 <= _tickers_x3_lfsrReg_T_671;
    end
    if (tickers_x3_lfsrReg_96 == 16'h0) begin
      tickers_x3_lfsrReg_96 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_96 <= _tickers_x3_lfsrReg_T_678;
    end
    if (tickers_x3_lfsrReg_97 == 16'h0) begin
      tickers_x3_lfsrReg_97 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_97 <= _tickers_x3_lfsrReg_T_685;
    end
    if (tickers_x3_lfsrReg_98 == 16'h0) begin
      tickers_x3_lfsrReg_98 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_98 <= _tickers_x3_lfsrReg_T_692;
    end
    if (tickers_x3_lfsrReg_99 == 16'h0) begin
      tickers_x3_lfsrReg_99 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_99 <= _tickers_x3_lfsrReg_T_699;
    end
    if (tickers_x3_lfsrReg_100 == 16'h0) begin
      tickers_x3_lfsrReg_100 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_100 <= _tickers_x3_lfsrReg_T_706;
    end
    if (tickers_x3_lfsrReg_101 == 16'h0) begin
      tickers_x3_lfsrReg_101 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_101 <= _tickers_x3_lfsrReg_T_713;
    end
    if (tickers_x3_lfsrReg_102 == 16'h0) begin
      tickers_x3_lfsrReg_102 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_102 <= _tickers_x3_lfsrReg_T_720;
    end
    if (tickers_x3_lfsrReg_103 == 16'h0) begin
      tickers_x3_lfsrReg_103 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_103 <= _tickers_x3_lfsrReg_T_727;
    end
    if (tickers_x3_lfsrReg_104 == 16'h0) begin
      tickers_x3_lfsrReg_104 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_104 <= _tickers_x3_lfsrReg_T_734;
    end
    if (tickers_x3_lfsrReg_105 == 16'h0) begin
      tickers_x3_lfsrReg_105 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_105 <= _tickers_x3_lfsrReg_T_741;
    end
    if (tickers_x3_lfsrReg_106 == 16'h0) begin
      tickers_x3_lfsrReg_106 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_106 <= _tickers_x3_lfsrReg_T_748;
    end
    if (tickers_x3_lfsrReg_107 == 16'h0) begin
      tickers_x3_lfsrReg_107 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_107 <= _tickers_x3_lfsrReg_T_755;
    end
    if (tickers_x3_lfsrReg_108 == 16'h0) begin
      tickers_x3_lfsrReg_108 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_108 <= _tickers_x3_lfsrReg_T_762;
    end
    if (tickers_x3_lfsrReg_109 == 16'h0) begin
      tickers_x3_lfsrReg_109 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_109 <= _tickers_x3_lfsrReg_T_769;
    end
    if (tickers_x3_lfsrReg_110 == 16'h0) begin
      tickers_x3_lfsrReg_110 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_110 <= _tickers_x3_lfsrReg_T_776;
    end
    if (tickers_x3_lfsrReg_111 == 16'h0) begin
      tickers_x3_lfsrReg_111 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_111 <= _tickers_x3_lfsrReg_T_783;
    end
    if (tickers_x3_lfsrReg_112 == 16'h0) begin
      tickers_x3_lfsrReg_112 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_112 <= _tickers_x3_lfsrReg_T_790;
    end
    if (tickers_x3_lfsrReg_113 == 16'h0) begin
      tickers_x3_lfsrReg_113 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_113 <= _tickers_x3_lfsrReg_T_797;
    end
    if (tickers_x3_lfsrReg_114 == 16'h0) begin
      tickers_x3_lfsrReg_114 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_114 <= _tickers_x3_lfsrReg_T_804;
    end
    if (tickers_x3_lfsrReg_115 == 16'h0) begin
      tickers_x3_lfsrReg_115 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_115 <= _tickers_x3_lfsrReg_T_811;
    end
    if (tickers_x3_lfsrReg_116 == 16'h0) begin
      tickers_x3_lfsrReg_116 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_116 <= _tickers_x3_lfsrReg_T_818;
    end
    if (tickers_x3_lfsrReg_117 == 16'h0) begin
      tickers_x3_lfsrReg_117 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_117 <= _tickers_x3_lfsrReg_T_825;
    end
    if (tickers_x3_lfsrReg_118 == 16'h0) begin
      tickers_x3_lfsrReg_118 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_118 <= _tickers_x3_lfsrReg_T_832;
    end
    if (tickers_x3_lfsrReg_119 == 16'h0) begin
      tickers_x3_lfsrReg_119 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_119 <= _tickers_x3_lfsrReg_T_839;
    end
    if (tickers_x3_lfsrReg_120 == 16'h0) begin
      tickers_x3_lfsrReg_120 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_120 <= _tickers_x3_lfsrReg_T_846;
    end
    if (tickers_x3_lfsrReg_121 == 16'h0) begin
      tickers_x3_lfsrReg_121 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_121 <= _tickers_x3_lfsrReg_T_853;
    end
    if (tickers_x3_lfsrReg_122 == 16'h0) begin
      tickers_x3_lfsrReg_122 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_122 <= _tickers_x3_lfsrReg_T_860;
    end
    if (tickers_x3_lfsrReg_123 == 16'h0) begin
      tickers_x3_lfsrReg_123 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_123 <= _tickers_x3_lfsrReg_T_867;
    end
    if (tickers_x3_lfsrReg_124 == 16'h0) begin
      tickers_x3_lfsrReg_124 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_124 <= _tickers_x3_lfsrReg_T_874;
    end
    if (tickers_x3_lfsrReg_125 == 16'h0) begin
      tickers_x3_lfsrReg_125 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_125 <= _tickers_x3_lfsrReg_T_881;
    end
    if (tickers_x3_lfsrReg_126 == 16'h0) begin
      tickers_x3_lfsrReg_126 <= 16'h1;
    end else begin
      tickers_x3_lfsrReg_126 <= _tickers_x3_lfsrReg_T_888;
    end
    if (tickers_x3_lfsrReg[0]) begin
      if (system_global_interrupts_x5_lfsrReg == 16'h0) begin
        system_global_interrupts_x5_lfsrReg <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg <= _system_global_interrupts_x5_lfsrReg_T_6;
      end
    end
    if (tickers_x3_lfsrReg_1[0]) begin
      if (system_global_interrupts_x5_lfsrReg_1 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_1 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_1 <= _system_global_interrupts_x5_lfsrReg_T_13;
      end
    end
    if (tickers_x3_lfsrReg_2[0]) begin
      if (system_global_interrupts_x5_lfsrReg_2 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_2 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_2 <= _system_global_interrupts_x5_lfsrReg_T_20;
      end
    end
    if (tickers_x3_lfsrReg_3[0]) begin
      if (system_global_interrupts_x5_lfsrReg_3 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_3 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_3 <= _system_global_interrupts_x5_lfsrReg_T_27;
      end
    end
    if (tickers_x3_lfsrReg_4[0]) begin
      if (system_global_interrupts_x5_lfsrReg_4 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_4 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_4 <= _system_global_interrupts_x5_lfsrReg_T_34;
      end
    end
    if (tickers_x3_lfsrReg_5[0]) begin
      if (system_global_interrupts_x5_lfsrReg_5 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_5 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_5 <= _system_global_interrupts_x5_lfsrReg_T_41;
      end
    end
    if (tickers_x3_lfsrReg_6[0]) begin
      if (system_global_interrupts_x5_lfsrReg_6 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_6 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_6 <= _system_global_interrupts_x5_lfsrReg_T_48;
      end
    end
    if (tickers_x3_lfsrReg_7[0]) begin
      if (system_global_interrupts_x5_lfsrReg_7 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_7 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_7 <= _system_global_interrupts_x5_lfsrReg_T_55;
      end
    end
    if (tickers_x3_lfsrReg_8[0]) begin
      if (system_global_interrupts_x5_lfsrReg_8 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_8 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_8 <= _system_global_interrupts_x5_lfsrReg_T_62;
      end
    end
    if (tickers_x3_lfsrReg_9[0]) begin
      if (system_global_interrupts_x5_lfsrReg_9 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_9 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_9 <= _system_global_interrupts_x5_lfsrReg_T_69;
      end
    end
    if (tickers_x3_lfsrReg_10[0]) begin
      if (system_global_interrupts_x5_lfsrReg_10 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_10 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_10 <= _system_global_interrupts_x5_lfsrReg_T_76;
      end
    end
    if (tickers_x3_lfsrReg_11[0]) begin
      if (system_global_interrupts_x5_lfsrReg_11 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_11 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_11 <= _system_global_interrupts_x5_lfsrReg_T_83;
      end
    end
    if (tickers_x3_lfsrReg_12[0]) begin
      if (system_global_interrupts_x5_lfsrReg_12 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_12 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_12 <= _system_global_interrupts_x5_lfsrReg_T_90;
      end
    end
    if (tickers_x3_lfsrReg_13[0]) begin
      if (system_global_interrupts_x5_lfsrReg_13 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_13 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_13 <= _system_global_interrupts_x5_lfsrReg_T_97;
      end
    end
    if (tickers_x3_lfsrReg_14[0]) begin
      if (system_global_interrupts_x5_lfsrReg_14 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_14 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_14 <= _system_global_interrupts_x5_lfsrReg_T_104;
      end
    end
    if (tickers_x3_lfsrReg_15[0]) begin
      if (system_global_interrupts_x5_lfsrReg_15 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_15 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_15 <= _system_global_interrupts_x5_lfsrReg_T_111;
      end
    end
    if (tickers_x3_lfsrReg_16[0]) begin
      if (system_global_interrupts_x5_lfsrReg_16 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_16 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_16 <= _system_global_interrupts_x5_lfsrReg_T_118;
      end
    end
    if (tickers_x3_lfsrReg_17[0]) begin
      if (system_global_interrupts_x5_lfsrReg_17 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_17 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_17 <= _system_global_interrupts_x5_lfsrReg_T_125;
      end
    end
    if (tickers_x3_lfsrReg_18[0]) begin
      if (system_global_interrupts_x5_lfsrReg_18 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_18 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_18 <= _system_global_interrupts_x5_lfsrReg_T_132;
      end
    end
    if (tickers_x3_lfsrReg_19[0]) begin
      if (system_global_interrupts_x5_lfsrReg_19 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_19 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_19 <= _system_global_interrupts_x5_lfsrReg_T_139;
      end
    end
    if (tickers_x3_lfsrReg_20[0]) begin
      if (system_global_interrupts_x5_lfsrReg_20 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_20 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_20 <= _system_global_interrupts_x5_lfsrReg_T_146;
      end
    end
    if (tickers_x3_lfsrReg_21[0]) begin
      if (system_global_interrupts_x5_lfsrReg_21 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_21 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_21 <= _system_global_interrupts_x5_lfsrReg_T_153;
      end
    end
    if (tickers_x3_lfsrReg_22[0]) begin
      if (system_global_interrupts_x5_lfsrReg_22 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_22 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_22 <= _system_global_interrupts_x5_lfsrReg_T_160;
      end
    end
    if (tickers_x3_lfsrReg_23[0]) begin
      if (system_global_interrupts_x5_lfsrReg_23 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_23 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_23 <= _system_global_interrupts_x5_lfsrReg_T_167;
      end
    end
    if (tickers_x3_lfsrReg_24[0]) begin
      if (system_global_interrupts_x5_lfsrReg_24 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_24 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_24 <= _system_global_interrupts_x5_lfsrReg_T_174;
      end
    end
    if (tickers_x3_lfsrReg_25[0]) begin
      if (system_global_interrupts_x5_lfsrReg_25 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_25 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_25 <= _system_global_interrupts_x5_lfsrReg_T_181;
      end
    end
    if (tickers_x3_lfsrReg_26[0]) begin
      if (system_global_interrupts_x5_lfsrReg_26 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_26 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_26 <= _system_global_interrupts_x5_lfsrReg_T_188;
      end
    end
    if (tickers_x3_lfsrReg_27[0]) begin
      if (system_global_interrupts_x5_lfsrReg_27 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_27 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_27 <= _system_global_interrupts_x5_lfsrReg_T_195;
      end
    end
    if (tickers_x3_lfsrReg_28[0]) begin
      if (system_global_interrupts_x5_lfsrReg_28 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_28 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_28 <= _system_global_interrupts_x5_lfsrReg_T_202;
      end
    end
    if (tickers_x3_lfsrReg_29[0]) begin
      if (system_global_interrupts_x5_lfsrReg_29 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_29 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_29 <= _system_global_interrupts_x5_lfsrReg_T_209;
      end
    end
    if (tickers_x3_lfsrReg_30[0]) begin
      if (system_global_interrupts_x5_lfsrReg_30 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_30 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_30 <= _system_global_interrupts_x5_lfsrReg_T_216;
      end
    end
    if (tickers_x3_lfsrReg_31[0]) begin
      if (system_global_interrupts_x5_lfsrReg_31 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_31 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_31 <= _system_global_interrupts_x5_lfsrReg_T_223;
      end
    end
    if (tickers_x3_lfsrReg_32[0]) begin
      if (system_global_interrupts_x5_lfsrReg_32 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_32 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_32 <= _system_global_interrupts_x5_lfsrReg_T_230;
      end
    end
    if (tickers_x3_lfsrReg_33[0]) begin
      if (system_global_interrupts_x5_lfsrReg_33 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_33 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_33 <= _system_global_interrupts_x5_lfsrReg_T_237;
      end
    end
    if (tickers_x3_lfsrReg_34[0]) begin
      if (system_global_interrupts_x5_lfsrReg_34 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_34 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_34 <= _system_global_interrupts_x5_lfsrReg_T_244;
      end
    end
    if (tickers_x3_lfsrReg_35[0]) begin
      if (system_global_interrupts_x5_lfsrReg_35 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_35 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_35 <= _system_global_interrupts_x5_lfsrReg_T_251;
      end
    end
    if (tickers_x3_lfsrReg_36[0]) begin
      if (system_global_interrupts_x5_lfsrReg_36 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_36 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_36 <= _system_global_interrupts_x5_lfsrReg_T_258;
      end
    end
    if (tickers_x3_lfsrReg_37[0]) begin
      if (system_global_interrupts_x5_lfsrReg_37 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_37 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_37 <= _system_global_interrupts_x5_lfsrReg_T_265;
      end
    end
    if (tickers_x3_lfsrReg_38[0]) begin
      if (system_global_interrupts_x5_lfsrReg_38 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_38 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_38 <= _system_global_interrupts_x5_lfsrReg_T_272;
      end
    end
    if (tickers_x3_lfsrReg_39[0]) begin
      if (system_global_interrupts_x5_lfsrReg_39 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_39 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_39 <= _system_global_interrupts_x5_lfsrReg_T_279;
      end
    end
    if (tickers_x3_lfsrReg_40[0]) begin
      if (system_global_interrupts_x5_lfsrReg_40 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_40 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_40 <= _system_global_interrupts_x5_lfsrReg_T_286;
      end
    end
    if (tickers_x3_lfsrReg_41[0]) begin
      if (system_global_interrupts_x5_lfsrReg_41 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_41 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_41 <= _system_global_interrupts_x5_lfsrReg_T_293;
      end
    end
    if (tickers_x3_lfsrReg_42[0]) begin
      if (system_global_interrupts_x5_lfsrReg_42 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_42 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_42 <= _system_global_interrupts_x5_lfsrReg_T_300;
      end
    end
    if (tickers_x3_lfsrReg_43[0]) begin
      if (system_global_interrupts_x5_lfsrReg_43 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_43 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_43 <= _system_global_interrupts_x5_lfsrReg_T_307;
      end
    end
    if (tickers_x3_lfsrReg_44[0]) begin
      if (system_global_interrupts_x5_lfsrReg_44 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_44 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_44 <= _system_global_interrupts_x5_lfsrReg_T_314;
      end
    end
    if (tickers_x3_lfsrReg_45[0]) begin
      if (system_global_interrupts_x5_lfsrReg_45 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_45 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_45 <= _system_global_interrupts_x5_lfsrReg_T_321;
      end
    end
    if (tickers_x3_lfsrReg_46[0]) begin
      if (system_global_interrupts_x5_lfsrReg_46 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_46 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_46 <= _system_global_interrupts_x5_lfsrReg_T_328;
      end
    end
    if (tickers_x3_lfsrReg_47[0]) begin
      if (system_global_interrupts_x5_lfsrReg_47 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_47 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_47 <= _system_global_interrupts_x5_lfsrReg_T_335;
      end
    end
    if (tickers_x3_lfsrReg_48[0]) begin
      if (system_global_interrupts_x5_lfsrReg_48 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_48 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_48 <= _system_global_interrupts_x5_lfsrReg_T_342;
      end
    end
    if (tickers_x3_lfsrReg_49[0]) begin
      if (system_global_interrupts_x5_lfsrReg_49 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_49 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_49 <= _system_global_interrupts_x5_lfsrReg_T_349;
      end
    end
    if (tickers_x3_lfsrReg_50[0]) begin
      if (system_global_interrupts_x5_lfsrReg_50 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_50 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_50 <= _system_global_interrupts_x5_lfsrReg_T_356;
      end
    end
    if (tickers_x3_lfsrReg_51[0]) begin
      if (system_global_interrupts_x5_lfsrReg_51 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_51 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_51 <= _system_global_interrupts_x5_lfsrReg_T_363;
      end
    end
    if (tickers_x3_lfsrReg_52[0]) begin
      if (system_global_interrupts_x5_lfsrReg_52 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_52 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_52 <= _system_global_interrupts_x5_lfsrReg_T_370;
      end
    end
    if (tickers_x3_lfsrReg_53[0]) begin
      if (system_global_interrupts_x5_lfsrReg_53 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_53 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_53 <= _system_global_interrupts_x5_lfsrReg_T_377;
      end
    end
    if (tickers_x3_lfsrReg_54[0]) begin
      if (system_global_interrupts_x5_lfsrReg_54 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_54 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_54 <= _system_global_interrupts_x5_lfsrReg_T_384;
      end
    end
    if (tickers_x3_lfsrReg_55[0]) begin
      if (system_global_interrupts_x5_lfsrReg_55 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_55 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_55 <= _system_global_interrupts_x5_lfsrReg_T_391;
      end
    end
    if (tickers_x3_lfsrReg_56[0]) begin
      if (system_global_interrupts_x5_lfsrReg_56 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_56 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_56 <= _system_global_interrupts_x5_lfsrReg_T_398;
      end
    end
    if (tickers_x3_lfsrReg_57[0]) begin
      if (system_global_interrupts_x5_lfsrReg_57 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_57 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_57 <= _system_global_interrupts_x5_lfsrReg_T_405;
      end
    end
    if (tickers_x3_lfsrReg_58[0]) begin
      if (system_global_interrupts_x5_lfsrReg_58 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_58 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_58 <= _system_global_interrupts_x5_lfsrReg_T_412;
      end
    end
    if (tickers_x3_lfsrReg_59[0]) begin
      if (system_global_interrupts_x5_lfsrReg_59 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_59 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_59 <= _system_global_interrupts_x5_lfsrReg_T_419;
      end
    end
    if (tickers_x3_lfsrReg_60[0]) begin
      if (system_global_interrupts_x5_lfsrReg_60 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_60 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_60 <= _system_global_interrupts_x5_lfsrReg_T_426;
      end
    end
    if (tickers_x3_lfsrReg_61[0]) begin
      if (system_global_interrupts_x5_lfsrReg_61 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_61 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_61 <= _system_global_interrupts_x5_lfsrReg_T_433;
      end
    end
    if (tickers_x3_lfsrReg_62[0]) begin
      if (system_global_interrupts_x5_lfsrReg_62 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_62 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_62 <= _system_global_interrupts_x5_lfsrReg_T_440;
      end
    end
    if (tickers_x3_lfsrReg_63[0]) begin
      if (system_global_interrupts_x5_lfsrReg_63 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_63 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_63 <= _system_global_interrupts_x5_lfsrReg_T_447;
      end
    end
    if (tickers_x3_lfsrReg_64[0]) begin
      if (system_global_interrupts_x5_lfsrReg_64 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_64 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_64 <= _system_global_interrupts_x5_lfsrReg_T_454;
      end
    end
    if (tickers_x3_lfsrReg_65[0]) begin
      if (system_global_interrupts_x5_lfsrReg_65 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_65 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_65 <= _system_global_interrupts_x5_lfsrReg_T_461;
      end
    end
    if (tickers_x3_lfsrReg_66[0]) begin
      if (system_global_interrupts_x5_lfsrReg_66 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_66 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_66 <= _system_global_interrupts_x5_lfsrReg_T_468;
      end
    end
    if (tickers_x3_lfsrReg_67[0]) begin
      if (system_global_interrupts_x5_lfsrReg_67 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_67 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_67 <= _system_global_interrupts_x5_lfsrReg_T_475;
      end
    end
    if (tickers_x3_lfsrReg_68[0]) begin
      if (system_global_interrupts_x5_lfsrReg_68 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_68 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_68 <= _system_global_interrupts_x5_lfsrReg_T_482;
      end
    end
    if (tickers_x3_lfsrReg_69[0]) begin
      if (system_global_interrupts_x5_lfsrReg_69 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_69 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_69 <= _system_global_interrupts_x5_lfsrReg_T_489;
      end
    end
    if (tickers_x3_lfsrReg_70[0]) begin
      if (system_global_interrupts_x5_lfsrReg_70 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_70 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_70 <= _system_global_interrupts_x5_lfsrReg_T_496;
      end
    end
    if (tickers_x3_lfsrReg_71[0]) begin
      if (system_global_interrupts_x5_lfsrReg_71 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_71 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_71 <= _system_global_interrupts_x5_lfsrReg_T_503;
      end
    end
    if (tickers_x3_lfsrReg_72[0]) begin
      if (system_global_interrupts_x5_lfsrReg_72 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_72 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_72 <= _system_global_interrupts_x5_lfsrReg_T_510;
      end
    end
    if (tickers_x3_lfsrReg_73[0]) begin
      if (system_global_interrupts_x5_lfsrReg_73 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_73 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_73 <= _system_global_interrupts_x5_lfsrReg_T_517;
      end
    end
    if (tickers_x3_lfsrReg_74[0]) begin
      if (system_global_interrupts_x5_lfsrReg_74 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_74 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_74 <= _system_global_interrupts_x5_lfsrReg_T_524;
      end
    end
    if (tickers_x3_lfsrReg_75[0]) begin
      if (system_global_interrupts_x5_lfsrReg_75 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_75 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_75 <= _system_global_interrupts_x5_lfsrReg_T_531;
      end
    end
    if (tickers_x3_lfsrReg_76[0]) begin
      if (system_global_interrupts_x5_lfsrReg_76 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_76 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_76 <= _system_global_interrupts_x5_lfsrReg_T_538;
      end
    end
    if (tickers_x3_lfsrReg_77[0]) begin
      if (system_global_interrupts_x5_lfsrReg_77 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_77 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_77 <= _system_global_interrupts_x5_lfsrReg_T_545;
      end
    end
    if (tickers_x3_lfsrReg_78[0]) begin
      if (system_global_interrupts_x5_lfsrReg_78 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_78 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_78 <= _system_global_interrupts_x5_lfsrReg_T_552;
      end
    end
    if (tickers_x3_lfsrReg_79[0]) begin
      if (system_global_interrupts_x5_lfsrReg_79 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_79 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_79 <= _system_global_interrupts_x5_lfsrReg_T_559;
      end
    end
    if (tickers_x3_lfsrReg_80[0]) begin
      if (system_global_interrupts_x5_lfsrReg_80 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_80 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_80 <= _system_global_interrupts_x5_lfsrReg_T_566;
      end
    end
    if (tickers_x3_lfsrReg_81[0]) begin
      if (system_global_interrupts_x5_lfsrReg_81 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_81 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_81 <= _system_global_interrupts_x5_lfsrReg_T_573;
      end
    end
    if (tickers_x3_lfsrReg_82[0]) begin
      if (system_global_interrupts_x5_lfsrReg_82 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_82 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_82 <= _system_global_interrupts_x5_lfsrReg_T_580;
      end
    end
    if (tickers_x3_lfsrReg_83[0]) begin
      if (system_global_interrupts_x5_lfsrReg_83 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_83 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_83 <= _system_global_interrupts_x5_lfsrReg_T_587;
      end
    end
    if (tickers_x3_lfsrReg_84[0]) begin
      if (system_global_interrupts_x5_lfsrReg_84 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_84 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_84 <= _system_global_interrupts_x5_lfsrReg_T_594;
      end
    end
    if (tickers_x3_lfsrReg_85[0]) begin
      if (system_global_interrupts_x5_lfsrReg_85 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_85 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_85 <= _system_global_interrupts_x5_lfsrReg_T_601;
      end
    end
    if (tickers_x3_lfsrReg_86[0]) begin
      if (system_global_interrupts_x5_lfsrReg_86 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_86 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_86 <= _system_global_interrupts_x5_lfsrReg_T_608;
      end
    end
    if (tickers_x3_lfsrReg_87[0]) begin
      if (system_global_interrupts_x5_lfsrReg_87 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_87 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_87 <= _system_global_interrupts_x5_lfsrReg_T_615;
      end
    end
    if (tickers_x3_lfsrReg_88[0]) begin
      if (system_global_interrupts_x5_lfsrReg_88 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_88 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_88 <= _system_global_interrupts_x5_lfsrReg_T_622;
      end
    end
    if (tickers_x3_lfsrReg_89[0]) begin
      if (system_global_interrupts_x5_lfsrReg_89 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_89 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_89 <= _system_global_interrupts_x5_lfsrReg_T_629;
      end
    end
    if (tickers_x3_lfsrReg_90[0]) begin
      if (system_global_interrupts_x5_lfsrReg_90 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_90 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_90 <= _system_global_interrupts_x5_lfsrReg_T_636;
      end
    end
    if (tickers_x3_lfsrReg_91[0]) begin
      if (system_global_interrupts_x5_lfsrReg_91 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_91 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_91 <= _system_global_interrupts_x5_lfsrReg_T_643;
      end
    end
    if (tickers_x3_lfsrReg_92[0]) begin
      if (system_global_interrupts_x5_lfsrReg_92 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_92 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_92 <= _system_global_interrupts_x5_lfsrReg_T_650;
      end
    end
    if (tickers_x3_lfsrReg_93[0]) begin
      if (system_global_interrupts_x5_lfsrReg_93 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_93 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_93 <= _system_global_interrupts_x5_lfsrReg_T_657;
      end
    end
    if (tickers_x3_lfsrReg_94[0]) begin
      if (system_global_interrupts_x5_lfsrReg_94 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_94 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_94 <= _system_global_interrupts_x5_lfsrReg_T_664;
      end
    end
    if (tickers_x3_lfsrReg_95[0]) begin
      if (system_global_interrupts_x5_lfsrReg_95 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_95 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_95 <= _system_global_interrupts_x5_lfsrReg_T_671;
      end
    end
    if (tickers_x3_lfsrReg_96[0]) begin
      if (system_global_interrupts_x5_lfsrReg_96 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_96 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_96 <= _system_global_interrupts_x5_lfsrReg_T_678;
      end
    end
    if (tickers_x3_lfsrReg_97[0]) begin
      if (system_global_interrupts_x5_lfsrReg_97 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_97 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_97 <= _system_global_interrupts_x5_lfsrReg_T_685;
      end
    end
    if (tickers_x3_lfsrReg_98[0]) begin
      if (system_global_interrupts_x5_lfsrReg_98 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_98 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_98 <= _system_global_interrupts_x5_lfsrReg_T_692;
      end
    end
    if (tickers_x3_lfsrReg_99[0]) begin
      if (system_global_interrupts_x5_lfsrReg_99 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_99 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_99 <= _system_global_interrupts_x5_lfsrReg_T_699;
      end
    end
    if (tickers_x3_lfsrReg_100[0]) begin
      if (system_global_interrupts_x5_lfsrReg_100 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_100 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_100 <= _system_global_interrupts_x5_lfsrReg_T_706;
      end
    end
    if (tickers_x3_lfsrReg_101[0]) begin
      if (system_global_interrupts_x5_lfsrReg_101 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_101 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_101 <= _system_global_interrupts_x5_lfsrReg_T_713;
      end
    end
    if (tickers_x3_lfsrReg_102[0]) begin
      if (system_global_interrupts_x5_lfsrReg_102 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_102 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_102 <= _system_global_interrupts_x5_lfsrReg_T_720;
      end
    end
    if (tickers_x3_lfsrReg_103[0]) begin
      if (system_global_interrupts_x5_lfsrReg_103 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_103 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_103 <= _system_global_interrupts_x5_lfsrReg_T_727;
      end
    end
    if (tickers_x3_lfsrReg_104[0]) begin
      if (system_global_interrupts_x5_lfsrReg_104 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_104 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_104 <= _system_global_interrupts_x5_lfsrReg_T_734;
      end
    end
    if (tickers_x3_lfsrReg_105[0]) begin
      if (system_global_interrupts_x5_lfsrReg_105 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_105 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_105 <= _system_global_interrupts_x5_lfsrReg_T_741;
      end
    end
    if (tickers_x3_lfsrReg_106[0]) begin
      if (system_global_interrupts_x5_lfsrReg_106 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_106 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_106 <= _system_global_interrupts_x5_lfsrReg_T_748;
      end
    end
    if (tickers_x3_lfsrReg_107[0]) begin
      if (system_global_interrupts_x5_lfsrReg_107 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_107 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_107 <= _system_global_interrupts_x5_lfsrReg_T_755;
      end
    end
    if (tickers_x3_lfsrReg_108[0]) begin
      if (system_global_interrupts_x5_lfsrReg_108 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_108 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_108 <= _system_global_interrupts_x5_lfsrReg_T_762;
      end
    end
    if (tickers_x3_lfsrReg_109[0]) begin
      if (system_global_interrupts_x5_lfsrReg_109 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_109 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_109 <= _system_global_interrupts_x5_lfsrReg_T_769;
      end
    end
    if (tickers_x3_lfsrReg_110[0]) begin
      if (system_global_interrupts_x5_lfsrReg_110 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_110 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_110 <= _system_global_interrupts_x5_lfsrReg_T_776;
      end
    end
    if (tickers_x3_lfsrReg_111[0]) begin
      if (system_global_interrupts_x5_lfsrReg_111 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_111 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_111 <= _system_global_interrupts_x5_lfsrReg_T_783;
      end
    end
    if (tickers_x3_lfsrReg_112[0]) begin
      if (system_global_interrupts_x5_lfsrReg_112 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_112 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_112 <= _system_global_interrupts_x5_lfsrReg_T_790;
      end
    end
    if (tickers_x3_lfsrReg_113[0]) begin
      if (system_global_interrupts_x5_lfsrReg_113 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_113 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_113 <= _system_global_interrupts_x5_lfsrReg_T_797;
      end
    end
    if (tickers_x3_lfsrReg_114[0]) begin
      if (system_global_interrupts_x5_lfsrReg_114 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_114 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_114 <= _system_global_interrupts_x5_lfsrReg_T_804;
      end
    end
    if (tickers_x3_lfsrReg_115[0]) begin
      if (system_global_interrupts_x5_lfsrReg_115 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_115 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_115 <= _system_global_interrupts_x5_lfsrReg_T_811;
      end
    end
    if (tickers_x3_lfsrReg_116[0]) begin
      if (system_global_interrupts_x5_lfsrReg_116 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_116 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_116 <= _system_global_interrupts_x5_lfsrReg_T_818;
      end
    end
    if (tickers_x3_lfsrReg_117[0]) begin
      if (system_global_interrupts_x5_lfsrReg_117 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_117 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_117 <= _system_global_interrupts_x5_lfsrReg_T_825;
      end
    end
    if (tickers_x3_lfsrReg_118[0]) begin
      if (system_global_interrupts_x5_lfsrReg_118 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_118 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_118 <= _system_global_interrupts_x5_lfsrReg_T_832;
      end
    end
    if (tickers_x3_lfsrReg_119[0]) begin
      if (system_global_interrupts_x5_lfsrReg_119 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_119 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_119 <= _system_global_interrupts_x5_lfsrReg_T_839;
      end
    end
    if (tickers_x3_lfsrReg_120[0]) begin
      if (system_global_interrupts_x5_lfsrReg_120 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_120 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_120 <= _system_global_interrupts_x5_lfsrReg_T_846;
      end
    end
    if (tickers_x3_lfsrReg_121[0]) begin
      if (system_global_interrupts_x5_lfsrReg_121 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_121 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_121 <= _system_global_interrupts_x5_lfsrReg_T_853;
      end
    end
    if (tickers_x3_lfsrReg_122[0]) begin
      if (system_global_interrupts_x5_lfsrReg_122 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_122 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_122 <= _system_global_interrupts_x5_lfsrReg_T_860;
      end
    end
    if (tickers_x3_lfsrReg_123[0]) begin
      if (system_global_interrupts_x5_lfsrReg_123 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_123 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_123 <= _system_global_interrupts_x5_lfsrReg_T_867;
      end
    end
    if (tickers_x3_lfsrReg_124[0]) begin
      if (system_global_interrupts_x5_lfsrReg_124 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_124 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_124 <= _system_global_interrupts_x5_lfsrReg_T_874;
      end
    end
    if (tickers_x3_lfsrReg_125[0]) begin
      if (system_global_interrupts_x5_lfsrReg_125 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_125 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_125 <= _system_global_interrupts_x5_lfsrReg_T_881;
      end
    end
    if (tickers_x3_lfsrReg_126[0]) begin
      if (system_global_interrupts_x5_lfsrReg_126 == 16'h0) begin
        system_global_interrupts_x5_lfsrReg_126 <= 16'h1;
      end else begin
        system_global_interrupts_x5_lfsrReg_126 <= _system_global_interrupts_x5_lfsrReg_T_888;
      end
    end
    if (reset) begin
      tick_value_1 <= 7'h0;
    end else if (tick_1) begin
      tick_value_1 <= 7'h0;
    end else begin
      tick_value_1 <= _tick_value_T_3;
    end
    if (reset) begin
      system_local_interrupts_0_value <= 4'h0;
    end else if (tick_1) begin
      system_local_interrupts_0_value <= _system_local_interrupts_0_wrap_value_T_1;
    end
    if (tick_1) begin
      if (tickers_x3_lfsrReg_127 == 16'h0) begin
        tickers_x3_lfsrReg_127 <= 16'h1;
      end else begin
        tickers_x3_lfsrReg_127 <= _tickers_x3_lfsrReg_T_895;
      end
    end
    if (tick_1) begin
      if (tickers_x3_lfsrReg_128 == 16'h0) begin
        tickers_x3_lfsrReg_128 <= 16'h1;
      end else begin
        tickers_x3_lfsrReg_128 <= _tickers_x3_lfsrReg_T_902;
      end
    end
    if (tick_1) begin
      if (tickers_x3_lfsrReg_129 == 16'h0) begin
        tickers_x3_lfsrReg_129 <= 16'h1;
      end else begin
        tickers_x3_lfsrReg_129 <= _tickers_x3_lfsrReg_T_909;
      end
    end
    if (tick_1) begin
      if (tickers_x3_lfsrReg_130 == 16'h0) begin
        tickers_x3_lfsrReg_130 <= 16'h1;
      end else begin
        tickers_x3_lfsrReg_130 <= _tickers_x3_lfsrReg_T_916;
      end
    end
    if (tick_1) begin
      if (tickers_x3_lfsrReg_131 == 16'h0) begin
        tickers_x3_lfsrReg_131 <= 16'h1;
      end else begin
        tickers_x3_lfsrReg_131 <= _tickers_x3_lfsrReg_T_923;
      end
    end
    if (tick_1) begin
      if (tickers_x3_lfsrReg_132 == 16'h0) begin
        tickers_x3_lfsrReg_132 <= 16'h1;
      end else begin
        tickers_x3_lfsrReg_132 <= _tickers_x3_lfsrReg_T_930;
      end
    end
    if (tick_1) begin
      if (tickers_x3_lfsrReg_133 == 16'h0) begin
        tickers_x3_lfsrReg_133 <= 16'h1;
      end else begin
        tickers_x3_lfsrReg_133 <= _tickers_x3_lfsrReg_T_937;
      end
    end
    if (tick_1) begin
      if (tickers_x3_lfsrReg_134 == 16'h0) begin
        tickers_x3_lfsrReg_134 <= 16'h1;
      end else begin
        tickers_x3_lfsrReg_134 <= _tickers_x3_lfsrReg_T_944;
      end
    end
    if (tick_1) begin
      if (tickers_x3_lfsrReg_135 == 16'h0) begin
        tickers_x3_lfsrReg_135 <= 16'h1;
      end else begin
        tickers_x3_lfsrReg_135 <= _tickers_x3_lfsrReg_T_951;
      end
    end
    if (tick_1) begin
      if (tickers_x3_lfsrReg_136 == 16'h0) begin
        tickers_x3_lfsrReg_136 <= 16'h1;
      end else begin
        tickers_x3_lfsrReg_136 <= _tickers_x3_lfsrReg_T_958;
      end
    end
    if (tick_1) begin
      if (tickers_x3_lfsrReg_137 == 16'h0) begin
        tickers_x3_lfsrReg_137 <= 16'h1;
      end else begin
        tickers_x3_lfsrReg_137 <= _tickers_x3_lfsrReg_T_965;
      end
    end
    if (tick_1) begin
      if (tickers_x3_lfsrReg_138 == 16'h0) begin
        tickers_x3_lfsrReg_138 <= 16'h1;
      end else begin
        tickers_x3_lfsrReg_138 <= _tickers_x3_lfsrReg_T_972;
      end
    end
    if (tick_1) begin
      if (tickers_x3_lfsrReg_139 == 16'h0) begin
        tickers_x3_lfsrReg_139 <= 16'h1;
      end else begin
        tickers_x3_lfsrReg_139 <= _tickers_x3_lfsrReg_T_979;
      end
    end
    if (tick_1) begin
      if (tickers_x3_lfsrReg_140 == 16'h0) begin
        tickers_x3_lfsrReg_140 <= 16'h1;
      end else begin
        tickers_x3_lfsrReg_140 <= _tickers_x3_lfsrReg_T_986;
      end
    end
    if (tick_1) begin
      if (tickers_x3_lfsrReg_141 == 16'h0) begin
        tickers_x3_lfsrReg_141 <= 16'h1;
      end else begin
        tickers_x3_lfsrReg_141 <= _tickers_x3_lfsrReg_T_993;
      end
    end
    if (tick_1) begin
      if (tickers_x3_lfsrReg_142 == 16'h0) begin
        tickers_x3_lfsrReg_142 <= 16'h1;
      end else begin
        tickers_x3_lfsrReg_142 <= _tickers_x3_lfsrReg_T_1000;
      end
    end
    if (tick_1) begin
      if (tickers_x5_lfsrReg == 16'h0) begin
        tickers_x5_lfsrReg <= 16'h1;
      end else begin
        tickers_x5_lfsrReg <= _tickers_x5_lfsrReg_T_6;
      end
    end
    if (tick_1) begin
      if (tickers_x5_lfsrReg_1 == 16'h0) begin
        tickers_x5_lfsrReg_1 <= 16'h1;
      end else begin
        tickers_x5_lfsrReg_1 <= _tickers_x5_lfsrReg_T_13;
      end
    end
    if (tick_1) begin
      if (tickers_x5_lfsrReg_2 == 16'h0) begin
        tickers_x5_lfsrReg_2 <= 16'h1;
      end else begin
        tickers_x5_lfsrReg_2 <= _tickers_x5_lfsrReg_T_20;
      end
    end
    if (tick_1) begin
      if (tickers_x5_lfsrReg_3 == 16'h0) begin
        tickers_x5_lfsrReg_3 <= 16'h1;
      end else begin
        tickers_x5_lfsrReg_3 <= _tickers_x5_lfsrReg_T_27;
      end
    end
    if (tick_1) begin
      if (tickers_x5_lfsrReg_4 == 16'h0) begin
        tickers_x5_lfsrReg_4 <= 16'h1;
      end else begin
        tickers_x5_lfsrReg_4 <= _tickers_x5_lfsrReg_T_34;
      end
    end
    if (tick_1) begin
      if (tickers_x5_lfsrReg_5 == 16'h0) begin
        tickers_x5_lfsrReg_5 <= 16'h1;
      end else begin
        tickers_x5_lfsrReg_5 <= _tickers_x5_lfsrReg_T_41;
      end
    end
    if (tick_1) begin
      if (tickers_x5_lfsrReg_6 == 16'h0) begin
        tickers_x5_lfsrReg_6 <= 16'h1;
      end else begin
        tickers_x5_lfsrReg_6 <= _tickers_x5_lfsrReg_T_48;
      end
    end
    if (tick_1) begin
      if (tickers_x5_lfsrReg_7 == 16'h0) begin
        tickers_x5_lfsrReg_7 <= 16'h1;
      end else begin
        tickers_x5_lfsrReg_7 <= _tickers_x5_lfsrReg_T_55;
      end
    end
    if (tick_1) begin
      if (tickers_x5_lfsrReg_8 == 16'h0) begin
        tickers_x5_lfsrReg_8 <= 16'h1;
      end else begin
        tickers_x5_lfsrReg_8 <= _tickers_x5_lfsrReg_T_62;
      end
    end
    if (tick_1) begin
      if (tickers_x5_lfsrReg_9 == 16'h0) begin
        tickers_x5_lfsrReg_9 <= 16'h1;
      end else begin
        tickers_x5_lfsrReg_9 <= _tickers_x5_lfsrReg_T_69;
      end
    end
    if (tick_1) begin
      if (tickers_x5_lfsrReg_10 == 16'h0) begin
        tickers_x5_lfsrReg_10 <= 16'h1;
      end else begin
        tickers_x5_lfsrReg_10 <= _tickers_x5_lfsrReg_T_76;
      end
    end
    if (tick_1) begin
      if (tickers_x5_lfsrReg_11 == 16'h0) begin
        tickers_x5_lfsrReg_11 <= 16'h1;
      end else begin
        tickers_x5_lfsrReg_11 <= _tickers_x5_lfsrReg_T_83;
      end
    end
    if (tick_1) begin
      if (tickers_x5_lfsrReg_12 == 16'h0) begin
        tickers_x5_lfsrReg_12 <= 16'h1;
      end else begin
        tickers_x5_lfsrReg_12 <= _tickers_x5_lfsrReg_T_90;
      end
    end
    if (tick_1) begin
      if (tickers_x5_lfsrReg_13 == 16'h0) begin
        tickers_x5_lfsrReg_13 <= 16'h1;
      end else begin
        tickers_x5_lfsrReg_13 <= _tickers_x5_lfsrReg_T_97;
      end
    end
    if (tick_1) begin
      if (tickers_x5_lfsrReg_14 == 16'h0) begin
        tickers_x5_lfsrReg_14 <= 16'h1;
      end else begin
        tickers_x5_lfsrReg_14 <= _tickers_x5_lfsrReg_T_104;
      end
    end
    if (tick_1) begin
      if (tickers_x5_lfsrReg_15 == 16'h0) begin
        tickers_x5_lfsrReg_15 <= 16'h1;
      end else begin
        tickers_x5_lfsrReg_15 <= _tickers_x5_lfsrReg_T_111;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(drive_interrupt_type == 32'h0) & ~(drive_interrupt_type == 32'h1) & ~(drive_interrupt_type == 32'h2) & ~(
          drive_interrupt_type == 32'h3) & ~(drive_interrupt_type == 32'h4) & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: DriveInterruptType.%d not supported yet\n    at Interrupts.scala:216 assert(false.B, \"DriveInterruptType.%%d not supported yet\", drive_interrupt_type)\n"
            ,drive_interrupt_type);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(drive_interrupt_type == 32'h0) & ~(drive_interrupt_type == 32'h1) & ~(drive_interrupt_type == 32'h2) & ~(
          drive_interrupt_type == 32'h3) & ~(drive_interrupt_type == 32'h4) & ~reset) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(drive_interrupt_type_1 == 32'h0) & ~(drive_interrupt_type_1 == 32'h1) & ~(drive_interrupt_type_1 == 32'h2)
           & ~(drive_interrupt_type_1 == 32'h3) & ~(drive_interrupt_type_1 == 32'h4) & ~(drive_interrupt_type_1 == 32'h5
          ) & ~reset) begin
          $fwrite(32'h80000002,
            "Assertion failed: DriveInterruptType.%d not supported yet\n    at InterruptDriver.scala:89 assert(false.B, \"DriveInterruptType.%%d not supported yet\", drive_interrupt_type)\n"
            ,drive_interrupt_type_1);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(drive_interrupt_type_1 == 32'h0) & ~(drive_interrupt_type_1 == 32'h1) & ~(drive_interrupt_type_1 == 32'h2)
           & ~(drive_interrupt_type_1 == 32'h3) & ~(drive_interrupt_type_1 == 32'h4) & ~(drive_interrupt_type_1 == 32'h5
          ) & ~reset) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  toggle = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  system_periph_port_ahb_0_hrdata_xs_io_valid_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  system_periph_port_ahb_0_hrdata_xs_io_valid_r_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  system_periph_port_ahb_0_hresp_xs_io_valid_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  system_sys_port_ahb_0_hrdata_xs_io_valid_r = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  system_sys_port_ahb_0_hrdata_xs_io_valid_r_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  system_sys_port_ahb_0_hresp_xs_io_valid_r = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  tick_value = _RAND_8[6:0];
  _RAND_9 = {1{`RANDOM}};
  system_global_interrupts_value = _RAND_9[6:0];
  _RAND_10 = {1{`RANDOM}};
  tickers_x3_lfsrReg = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  tickers_x3_lfsrReg_1 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  tickers_x3_lfsrReg_2 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  tickers_x3_lfsrReg_3 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  tickers_x3_lfsrReg_4 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  tickers_x3_lfsrReg_5 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  tickers_x3_lfsrReg_6 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  tickers_x3_lfsrReg_7 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  tickers_x3_lfsrReg_8 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  tickers_x3_lfsrReg_9 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  tickers_x3_lfsrReg_10 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  tickers_x3_lfsrReg_11 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  tickers_x3_lfsrReg_12 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  tickers_x3_lfsrReg_13 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  tickers_x3_lfsrReg_14 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  tickers_x3_lfsrReg_15 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  tickers_x3_lfsrReg_16 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  tickers_x3_lfsrReg_17 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  tickers_x3_lfsrReg_18 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  tickers_x3_lfsrReg_19 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  tickers_x3_lfsrReg_20 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  tickers_x3_lfsrReg_21 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  tickers_x3_lfsrReg_22 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  tickers_x3_lfsrReg_23 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  tickers_x3_lfsrReg_24 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  tickers_x3_lfsrReg_25 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  tickers_x3_lfsrReg_26 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  tickers_x3_lfsrReg_27 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  tickers_x3_lfsrReg_28 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  tickers_x3_lfsrReg_29 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  tickers_x3_lfsrReg_30 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  tickers_x3_lfsrReg_31 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  tickers_x3_lfsrReg_32 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  tickers_x3_lfsrReg_33 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  tickers_x3_lfsrReg_34 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  tickers_x3_lfsrReg_35 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  tickers_x3_lfsrReg_36 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  tickers_x3_lfsrReg_37 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  tickers_x3_lfsrReg_38 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  tickers_x3_lfsrReg_39 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  tickers_x3_lfsrReg_40 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  tickers_x3_lfsrReg_41 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  tickers_x3_lfsrReg_42 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  tickers_x3_lfsrReg_43 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  tickers_x3_lfsrReg_44 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  tickers_x3_lfsrReg_45 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  tickers_x3_lfsrReg_46 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  tickers_x3_lfsrReg_47 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  tickers_x3_lfsrReg_48 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  tickers_x3_lfsrReg_49 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  tickers_x3_lfsrReg_50 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  tickers_x3_lfsrReg_51 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  tickers_x3_lfsrReg_52 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  tickers_x3_lfsrReg_53 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  tickers_x3_lfsrReg_54 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  tickers_x3_lfsrReg_55 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  tickers_x3_lfsrReg_56 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  tickers_x3_lfsrReg_57 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  tickers_x3_lfsrReg_58 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  tickers_x3_lfsrReg_59 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  tickers_x3_lfsrReg_60 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  tickers_x3_lfsrReg_61 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  tickers_x3_lfsrReg_62 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  tickers_x3_lfsrReg_63 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  tickers_x3_lfsrReg_64 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  tickers_x3_lfsrReg_65 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  tickers_x3_lfsrReg_66 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  tickers_x3_lfsrReg_67 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  tickers_x3_lfsrReg_68 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  tickers_x3_lfsrReg_69 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  tickers_x3_lfsrReg_70 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  tickers_x3_lfsrReg_71 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  tickers_x3_lfsrReg_72 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  tickers_x3_lfsrReg_73 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  tickers_x3_lfsrReg_74 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  tickers_x3_lfsrReg_75 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  tickers_x3_lfsrReg_76 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  tickers_x3_lfsrReg_77 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  tickers_x3_lfsrReg_78 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  tickers_x3_lfsrReg_79 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  tickers_x3_lfsrReg_80 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  tickers_x3_lfsrReg_81 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  tickers_x3_lfsrReg_82 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  tickers_x3_lfsrReg_83 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  tickers_x3_lfsrReg_84 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  tickers_x3_lfsrReg_85 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  tickers_x3_lfsrReg_86 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  tickers_x3_lfsrReg_87 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  tickers_x3_lfsrReg_88 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  tickers_x3_lfsrReg_89 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  tickers_x3_lfsrReg_90 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  tickers_x3_lfsrReg_91 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  tickers_x3_lfsrReg_92 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  tickers_x3_lfsrReg_93 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  tickers_x3_lfsrReg_94 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  tickers_x3_lfsrReg_95 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  tickers_x3_lfsrReg_96 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  tickers_x3_lfsrReg_97 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  tickers_x3_lfsrReg_98 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  tickers_x3_lfsrReg_99 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  tickers_x3_lfsrReg_100 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  tickers_x3_lfsrReg_101 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  tickers_x3_lfsrReg_102 = _RAND_112[15:0];
  _RAND_113 = {1{`RANDOM}};
  tickers_x3_lfsrReg_103 = _RAND_113[15:0];
  _RAND_114 = {1{`RANDOM}};
  tickers_x3_lfsrReg_104 = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  tickers_x3_lfsrReg_105 = _RAND_115[15:0];
  _RAND_116 = {1{`RANDOM}};
  tickers_x3_lfsrReg_106 = _RAND_116[15:0];
  _RAND_117 = {1{`RANDOM}};
  tickers_x3_lfsrReg_107 = _RAND_117[15:0];
  _RAND_118 = {1{`RANDOM}};
  tickers_x3_lfsrReg_108 = _RAND_118[15:0];
  _RAND_119 = {1{`RANDOM}};
  tickers_x3_lfsrReg_109 = _RAND_119[15:0];
  _RAND_120 = {1{`RANDOM}};
  tickers_x3_lfsrReg_110 = _RAND_120[15:0];
  _RAND_121 = {1{`RANDOM}};
  tickers_x3_lfsrReg_111 = _RAND_121[15:0];
  _RAND_122 = {1{`RANDOM}};
  tickers_x3_lfsrReg_112 = _RAND_122[15:0];
  _RAND_123 = {1{`RANDOM}};
  tickers_x3_lfsrReg_113 = _RAND_123[15:0];
  _RAND_124 = {1{`RANDOM}};
  tickers_x3_lfsrReg_114 = _RAND_124[15:0];
  _RAND_125 = {1{`RANDOM}};
  tickers_x3_lfsrReg_115 = _RAND_125[15:0];
  _RAND_126 = {1{`RANDOM}};
  tickers_x3_lfsrReg_116 = _RAND_126[15:0];
  _RAND_127 = {1{`RANDOM}};
  tickers_x3_lfsrReg_117 = _RAND_127[15:0];
  _RAND_128 = {1{`RANDOM}};
  tickers_x3_lfsrReg_118 = _RAND_128[15:0];
  _RAND_129 = {1{`RANDOM}};
  tickers_x3_lfsrReg_119 = _RAND_129[15:0];
  _RAND_130 = {1{`RANDOM}};
  tickers_x3_lfsrReg_120 = _RAND_130[15:0];
  _RAND_131 = {1{`RANDOM}};
  tickers_x3_lfsrReg_121 = _RAND_131[15:0];
  _RAND_132 = {1{`RANDOM}};
  tickers_x3_lfsrReg_122 = _RAND_132[15:0];
  _RAND_133 = {1{`RANDOM}};
  tickers_x3_lfsrReg_123 = _RAND_133[15:0];
  _RAND_134 = {1{`RANDOM}};
  tickers_x3_lfsrReg_124 = _RAND_134[15:0];
  _RAND_135 = {1{`RANDOM}};
  tickers_x3_lfsrReg_125 = _RAND_135[15:0];
  _RAND_136 = {1{`RANDOM}};
  tickers_x3_lfsrReg_126 = _RAND_136[15:0];
  _RAND_137 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg = _RAND_137[15:0];
  _RAND_138 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_1 = _RAND_138[15:0];
  _RAND_139 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_2 = _RAND_139[15:0];
  _RAND_140 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_3 = _RAND_140[15:0];
  _RAND_141 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_4 = _RAND_141[15:0];
  _RAND_142 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_5 = _RAND_142[15:0];
  _RAND_143 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_6 = _RAND_143[15:0];
  _RAND_144 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_7 = _RAND_144[15:0];
  _RAND_145 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_8 = _RAND_145[15:0];
  _RAND_146 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_9 = _RAND_146[15:0];
  _RAND_147 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_10 = _RAND_147[15:0];
  _RAND_148 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_11 = _RAND_148[15:0];
  _RAND_149 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_12 = _RAND_149[15:0];
  _RAND_150 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_13 = _RAND_150[15:0];
  _RAND_151 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_14 = _RAND_151[15:0];
  _RAND_152 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_15 = _RAND_152[15:0];
  _RAND_153 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_16 = _RAND_153[15:0];
  _RAND_154 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_17 = _RAND_154[15:0];
  _RAND_155 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_18 = _RAND_155[15:0];
  _RAND_156 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_19 = _RAND_156[15:0];
  _RAND_157 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_20 = _RAND_157[15:0];
  _RAND_158 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_21 = _RAND_158[15:0];
  _RAND_159 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_22 = _RAND_159[15:0];
  _RAND_160 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_23 = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_24 = _RAND_161[15:0];
  _RAND_162 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_25 = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_26 = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_27 = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_28 = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_29 = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_30 = _RAND_167[15:0];
  _RAND_168 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_31 = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_32 = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_33 = _RAND_170[15:0];
  _RAND_171 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_34 = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_35 = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_36 = _RAND_173[15:0];
  _RAND_174 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_37 = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_38 = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_39 = _RAND_176[15:0];
  _RAND_177 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_40 = _RAND_177[15:0];
  _RAND_178 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_41 = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_42 = _RAND_179[15:0];
  _RAND_180 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_43 = _RAND_180[15:0];
  _RAND_181 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_44 = _RAND_181[15:0];
  _RAND_182 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_45 = _RAND_182[15:0];
  _RAND_183 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_46 = _RAND_183[15:0];
  _RAND_184 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_47 = _RAND_184[15:0];
  _RAND_185 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_48 = _RAND_185[15:0];
  _RAND_186 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_49 = _RAND_186[15:0];
  _RAND_187 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_50 = _RAND_187[15:0];
  _RAND_188 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_51 = _RAND_188[15:0];
  _RAND_189 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_52 = _RAND_189[15:0];
  _RAND_190 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_53 = _RAND_190[15:0];
  _RAND_191 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_54 = _RAND_191[15:0];
  _RAND_192 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_55 = _RAND_192[15:0];
  _RAND_193 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_56 = _RAND_193[15:0];
  _RAND_194 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_57 = _RAND_194[15:0];
  _RAND_195 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_58 = _RAND_195[15:0];
  _RAND_196 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_59 = _RAND_196[15:0];
  _RAND_197 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_60 = _RAND_197[15:0];
  _RAND_198 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_61 = _RAND_198[15:0];
  _RAND_199 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_62 = _RAND_199[15:0];
  _RAND_200 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_63 = _RAND_200[15:0];
  _RAND_201 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_64 = _RAND_201[15:0];
  _RAND_202 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_65 = _RAND_202[15:0];
  _RAND_203 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_66 = _RAND_203[15:0];
  _RAND_204 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_67 = _RAND_204[15:0];
  _RAND_205 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_68 = _RAND_205[15:0];
  _RAND_206 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_69 = _RAND_206[15:0];
  _RAND_207 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_70 = _RAND_207[15:0];
  _RAND_208 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_71 = _RAND_208[15:0];
  _RAND_209 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_72 = _RAND_209[15:0];
  _RAND_210 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_73 = _RAND_210[15:0];
  _RAND_211 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_74 = _RAND_211[15:0];
  _RAND_212 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_75 = _RAND_212[15:0];
  _RAND_213 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_76 = _RAND_213[15:0];
  _RAND_214 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_77 = _RAND_214[15:0];
  _RAND_215 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_78 = _RAND_215[15:0];
  _RAND_216 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_79 = _RAND_216[15:0];
  _RAND_217 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_80 = _RAND_217[15:0];
  _RAND_218 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_81 = _RAND_218[15:0];
  _RAND_219 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_82 = _RAND_219[15:0];
  _RAND_220 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_83 = _RAND_220[15:0];
  _RAND_221 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_84 = _RAND_221[15:0];
  _RAND_222 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_85 = _RAND_222[15:0];
  _RAND_223 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_86 = _RAND_223[15:0];
  _RAND_224 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_87 = _RAND_224[15:0];
  _RAND_225 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_88 = _RAND_225[15:0];
  _RAND_226 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_89 = _RAND_226[15:0];
  _RAND_227 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_90 = _RAND_227[15:0];
  _RAND_228 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_91 = _RAND_228[15:0];
  _RAND_229 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_92 = _RAND_229[15:0];
  _RAND_230 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_93 = _RAND_230[15:0];
  _RAND_231 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_94 = _RAND_231[15:0];
  _RAND_232 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_95 = _RAND_232[15:0];
  _RAND_233 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_96 = _RAND_233[15:0];
  _RAND_234 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_97 = _RAND_234[15:0];
  _RAND_235 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_98 = _RAND_235[15:0];
  _RAND_236 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_99 = _RAND_236[15:0];
  _RAND_237 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_100 = _RAND_237[15:0];
  _RAND_238 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_101 = _RAND_238[15:0];
  _RAND_239 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_102 = _RAND_239[15:0];
  _RAND_240 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_103 = _RAND_240[15:0];
  _RAND_241 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_104 = _RAND_241[15:0];
  _RAND_242 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_105 = _RAND_242[15:0];
  _RAND_243 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_106 = _RAND_243[15:0];
  _RAND_244 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_107 = _RAND_244[15:0];
  _RAND_245 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_108 = _RAND_245[15:0];
  _RAND_246 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_109 = _RAND_246[15:0];
  _RAND_247 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_110 = _RAND_247[15:0];
  _RAND_248 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_111 = _RAND_248[15:0];
  _RAND_249 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_112 = _RAND_249[15:0];
  _RAND_250 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_113 = _RAND_250[15:0];
  _RAND_251 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_114 = _RAND_251[15:0];
  _RAND_252 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_115 = _RAND_252[15:0];
  _RAND_253 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_116 = _RAND_253[15:0];
  _RAND_254 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_117 = _RAND_254[15:0];
  _RAND_255 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_118 = _RAND_255[15:0];
  _RAND_256 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_119 = _RAND_256[15:0];
  _RAND_257 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_120 = _RAND_257[15:0];
  _RAND_258 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_121 = _RAND_258[15:0];
  _RAND_259 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_122 = _RAND_259[15:0];
  _RAND_260 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_123 = _RAND_260[15:0];
  _RAND_261 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_124 = _RAND_261[15:0];
  _RAND_262 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_125 = _RAND_262[15:0];
  _RAND_263 = {1{`RANDOM}};
  system_global_interrupts_x5_lfsrReg_126 = _RAND_263[15:0];
  _RAND_264 = {1{`RANDOM}};
  tick_value_1 = _RAND_264[6:0];
  _RAND_265 = {1{`RANDOM}};
  system_local_interrupts_0_value = _RAND_265[3:0];
  _RAND_266 = {1{`RANDOM}};
  tickers_x3_lfsrReg_127 = _RAND_266[15:0];
  _RAND_267 = {1{`RANDOM}};
  tickers_x3_lfsrReg_128 = _RAND_267[15:0];
  _RAND_268 = {1{`RANDOM}};
  tickers_x3_lfsrReg_129 = _RAND_268[15:0];
  _RAND_269 = {1{`RANDOM}};
  tickers_x3_lfsrReg_130 = _RAND_269[15:0];
  _RAND_270 = {1{`RANDOM}};
  tickers_x3_lfsrReg_131 = _RAND_270[15:0];
  _RAND_271 = {1{`RANDOM}};
  tickers_x3_lfsrReg_132 = _RAND_271[15:0];
  _RAND_272 = {1{`RANDOM}};
  tickers_x3_lfsrReg_133 = _RAND_272[15:0];
  _RAND_273 = {1{`RANDOM}};
  tickers_x3_lfsrReg_134 = _RAND_273[15:0];
  _RAND_274 = {1{`RANDOM}};
  tickers_x3_lfsrReg_135 = _RAND_274[15:0];
  _RAND_275 = {1{`RANDOM}};
  tickers_x3_lfsrReg_136 = _RAND_275[15:0];
  _RAND_276 = {1{`RANDOM}};
  tickers_x3_lfsrReg_137 = _RAND_276[15:0];
  _RAND_277 = {1{`RANDOM}};
  tickers_x3_lfsrReg_138 = _RAND_277[15:0];
  _RAND_278 = {1{`RANDOM}};
  tickers_x3_lfsrReg_139 = _RAND_278[15:0];
  _RAND_279 = {1{`RANDOM}};
  tickers_x3_lfsrReg_140 = _RAND_279[15:0];
  _RAND_280 = {1{`RANDOM}};
  tickers_x3_lfsrReg_141 = _RAND_280[15:0];
  _RAND_281 = {1{`RANDOM}};
  tickers_x3_lfsrReg_142 = _RAND_281[15:0];
  _RAND_282 = {1{`RANDOM}};
  tickers_x5_lfsrReg = _RAND_282[15:0];
  _RAND_283 = {1{`RANDOM}};
  tickers_x5_lfsrReg_1 = _RAND_283[15:0];
  _RAND_284 = {1{`RANDOM}};
  tickers_x5_lfsrReg_2 = _RAND_284[15:0];
  _RAND_285 = {1{`RANDOM}};
  tickers_x5_lfsrReg_3 = _RAND_285[15:0];
  _RAND_286 = {1{`RANDOM}};
  tickers_x5_lfsrReg_4 = _RAND_286[15:0];
  _RAND_287 = {1{`RANDOM}};
  tickers_x5_lfsrReg_5 = _RAND_287[15:0];
  _RAND_288 = {1{`RANDOM}};
  tickers_x5_lfsrReg_6 = _RAND_288[15:0];
  _RAND_289 = {1{`RANDOM}};
  tickers_x5_lfsrReg_7 = _RAND_289[15:0];
  _RAND_290 = {1{`RANDOM}};
  tickers_x5_lfsrReg_8 = _RAND_290[15:0];
  _RAND_291 = {1{`RANDOM}};
  tickers_x5_lfsrReg_9 = _RAND_291[15:0];
  _RAND_292 = {1{`RANDOM}};
  tickers_x5_lfsrReg_10 = _RAND_292[15:0];
  _RAND_293 = {1{`RANDOM}};
  tickers_x5_lfsrReg_11 = _RAND_293[15:0];
  _RAND_294 = {1{`RANDOM}};
  tickers_x5_lfsrReg_12 = _RAND_294[15:0];
  _RAND_295 = {1{`RANDOM}};
  tickers_x5_lfsrReg_13 = _RAND_295[15:0];
  _RAND_296 = {1{`RANDOM}};
  tickers_x5_lfsrReg_14 = _RAND_296[15:0];
  _RAND_297 = {1{`RANDOM}};
  tickers_x5_lfsrReg_15 = _RAND_297[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
