//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_12(
  input  [31:0] _EVAL,
  input         _EVAL_0,
  output        _EVAL_1,
  input  [31:0] _EVAL_2,
  input  [3:0]  _EVAL_3,
  input  [3:0]  _EVAL_4,
  output [31:0] _EVAL_5,
  output [2:0]  _EVAL_6,
  output        _EVAL_7,
  output        _EVAL_8,
  output [31:0] _EVAL_9,
  output [3:0]  _EVAL_10,
  output        _EVAL_11,
  input  [3:0]  _EVAL_12,
  input  [2:0]  _EVAL_13,
  input         _EVAL_14,
  output [31:0] _EVAL_15,
  input  [3:0]  _EVAL_16,
  output [2:0]  _EVAL_17,
  input         _EVAL_18,
  input         _EVAL_19,
  output [3:0]  _EVAL_20,
  input         _EVAL_21,
  input  [2:0]  _EVAL_22,
  output [3:0]  _EVAL_23,
  input  [3:0]  _EVAL_24,
  output [2:0]  _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  output [3:0]  _EVAL_28,
  output        _EVAL_29,
  input         _EVAL_30,
  output        _EVAL_31,
  output [3:0]  _EVAL_32,
  input         _EVAL_33,
  output [1:0]  _EVAL_34,
  output        _EVAL_35,
  input  [1:0]  _EVAL_36,
  input         _EVAL_37,
  output [3:0]  _EVAL_38,
  output [1:0]  _EVAL_39,
  output [2:0]  _EVAL_40,
  output        _EVAL_41,
  output        _EVAL_42,
  input         _EVAL_43,
  input  [1:0]  _EVAL_44,
  input  [31:0] _EVAL_45,
  input         _EVAL_46,
  input  [2:0]  _EVAL_47,
  input         _EVAL_48,
  input  [2:0]  _EVAL_49,
  input  [3:0]  _EVAL_50,
  input         _EVAL_51,
  output [3:0]  _EVAL_52,
  output        _EVAL_53,
  output        _EVAL_54,
  output [1:0]  _EVAL_55,
  input  [3:0]  _EVAL_56,
  input         _EVAL_57,
  input         _EVAL_58,
  output        _EVAL_59,
  input  [2:0]  _EVAL_60,
  input  [31:0] _EVAL_61,
  input  [1:0]  _EVAL_62,
  input         _EVAL_63,
  input         _EVAL_64,
  output        _EVAL_65,
  input         _EVAL_66,
  output [31:0] _EVAL_67,
  input  [3:0]  _EVAL_68,
  input  [31:0] _EVAL_69,
  output [1:0]  _EVAL_70,
  output        _EVAL_71,
  output        _EVAL_72
);
  wire [3:0] rsink__EVAL;
  wire [31:0] rsink__EVAL_0;
  wire [1:0] rsink__EVAL_1;
  wire  rsink__EVAL_2;
  wire [1:0] rsink__EVAL_3;
  wire  rsink__EVAL_4;
  wire  rsink__EVAL_5;
  wire [2:0] rsink__EVAL_6;
  wire [3:0] rsink__EVAL_7;
  wire [3:0] rsink__EVAL_8;
  wire [3:0] rsink__EVAL_9;
  wire [3:0] rsink__EVAL_10;
  wire  rsink__EVAL_11;
  wire [2:0] rsink__EVAL_12;
  wire  rsink__EVAL_13;
  wire [3:0] rsink__EVAL_14;
  wire  rsink__EVAL_15;
  wire  rsink__EVAL_16;
  wire  rsink__EVAL_17;
  wire  rsink__EVAL_18;
  wire [3:0] rsink__EVAL_19;
  wire  rsink__EVAL_20;
  wire  rsink__EVAL_21;
  wire [3:0] rsink__EVAL_22;
  wire  rsink__EVAL_23;
  wire  rsink__EVAL_24;
  wire [2:0] rsink__EVAL_25;
  wire  rsink__EVAL_26;
  wire [3:0] rsink__EVAL_27;
  wire [31:0] rsink__EVAL_28;
  wire [2:0] rsink__EVAL_29;
  wire [31:0] rsink__EVAL_30;
  wire  rsink__EVAL_31;
  wire [1:0] rsink__EVAL_32;
  wire [31:0] rsink__EVAL_33;
  wire  rsink__EVAL_34;
  wire [3:0] rsink__EVAL_35;
  wire  rsink__EVAL_36;
  wire  rsink__EVAL_37;
  wire  rsink__EVAL_38;
  wire  rsink__EVAL_39;
  wire [3:0] rsink__EVAL_40;
  wire  rsink__EVAL_41;
  wire [2:0] rsink__EVAL_42;
  wire [31:0] rsink__EVAL_43;
  wire [3:0] rsink__EVAL_44;
  wire  rsink__EVAL_45;
  wire [31:0] rsink__EVAL_46;
  wire [1:0] rsink__EVAL_47;
  wire [2:0] rsink__EVAL_48;
  wire [3:0] rsink__EVAL_49;
  wire  rsink__EVAL_50;
  wire [3:0] rsink__EVAL_51;
  wire [2:0] rsink__EVAL_52;
  wire [3:0] rsink__EVAL_53;
  wire  rsink__EVAL_54;
  wire [2:0] rsink__EVAL_55;
  wire  rsink__EVAL_56;
  wire [1:0] rsink__EVAL_57;
  wire  rsink__EVAL_58;
  wire  rsink__EVAL_59;
  wire  rsink__EVAL_60;
  wire [2:0] rsink__EVAL_61;
  wire [1:0] rsink__EVAL_62;
  wire  rsink__EVAL_63;
  wire [31:0] rsink__EVAL_64;
  wire  rsink__EVAL_65;
  wire [1:0] rsink__EVAL_66;
  wire  rsink__EVAL_67;
  wire  rsink__EVAL_68;
  wire  rsink__EVAL_69;
  wire  rsink__EVAL_70;
  wire [31:0] rsink__EVAL_71;
  wire [31:0] rsink__EVAL_72;
  _EVAL_11 rsink (
    ._EVAL(rsink__EVAL),
    ._EVAL_0(rsink__EVAL_0),
    ._EVAL_1(rsink__EVAL_1),
    ._EVAL_2(rsink__EVAL_2),
    ._EVAL_3(rsink__EVAL_3),
    ._EVAL_4(rsink__EVAL_4),
    ._EVAL_5(rsink__EVAL_5),
    ._EVAL_6(rsink__EVAL_6),
    ._EVAL_7(rsink__EVAL_7),
    ._EVAL_8(rsink__EVAL_8),
    ._EVAL_9(rsink__EVAL_9),
    ._EVAL_10(rsink__EVAL_10),
    ._EVAL_11(rsink__EVAL_11),
    ._EVAL_12(rsink__EVAL_12),
    ._EVAL_13(rsink__EVAL_13),
    ._EVAL_14(rsink__EVAL_14),
    ._EVAL_15(rsink__EVAL_15),
    ._EVAL_16(rsink__EVAL_16),
    ._EVAL_17(rsink__EVAL_17),
    ._EVAL_18(rsink__EVAL_18),
    ._EVAL_19(rsink__EVAL_19),
    ._EVAL_20(rsink__EVAL_20),
    ._EVAL_21(rsink__EVAL_21),
    ._EVAL_22(rsink__EVAL_22),
    ._EVAL_23(rsink__EVAL_23),
    ._EVAL_24(rsink__EVAL_24),
    ._EVAL_25(rsink__EVAL_25),
    ._EVAL_26(rsink__EVAL_26),
    ._EVAL_27(rsink__EVAL_27),
    ._EVAL_28(rsink__EVAL_28),
    ._EVAL_29(rsink__EVAL_29),
    ._EVAL_30(rsink__EVAL_30),
    ._EVAL_31(rsink__EVAL_31),
    ._EVAL_32(rsink__EVAL_32),
    ._EVAL_33(rsink__EVAL_33),
    ._EVAL_34(rsink__EVAL_34),
    ._EVAL_35(rsink__EVAL_35),
    ._EVAL_36(rsink__EVAL_36),
    ._EVAL_37(rsink__EVAL_37),
    ._EVAL_38(rsink__EVAL_38),
    ._EVAL_39(rsink__EVAL_39),
    ._EVAL_40(rsink__EVAL_40),
    ._EVAL_41(rsink__EVAL_41),
    ._EVAL_42(rsink__EVAL_42),
    ._EVAL_43(rsink__EVAL_43),
    ._EVAL_44(rsink__EVAL_44),
    ._EVAL_45(rsink__EVAL_45),
    ._EVAL_46(rsink__EVAL_46),
    ._EVAL_47(rsink__EVAL_47),
    ._EVAL_48(rsink__EVAL_48),
    ._EVAL_49(rsink__EVAL_49),
    ._EVAL_50(rsink__EVAL_50),
    ._EVAL_51(rsink__EVAL_51),
    ._EVAL_52(rsink__EVAL_52),
    ._EVAL_53(rsink__EVAL_53),
    ._EVAL_54(rsink__EVAL_54),
    ._EVAL_55(rsink__EVAL_55),
    ._EVAL_56(rsink__EVAL_56),
    ._EVAL_57(rsink__EVAL_57),
    ._EVAL_58(rsink__EVAL_58),
    ._EVAL_59(rsink__EVAL_59),
    ._EVAL_60(rsink__EVAL_60),
    ._EVAL_61(rsink__EVAL_61),
    ._EVAL_62(rsink__EVAL_62),
    ._EVAL_63(rsink__EVAL_63),
    ._EVAL_64(rsink__EVAL_64),
    ._EVAL_65(rsink__EVAL_65),
    ._EVAL_66(rsink__EVAL_66),
    ._EVAL_67(rsink__EVAL_67),
    ._EVAL_68(rsink__EVAL_68),
    ._EVAL_69(rsink__EVAL_69),
    ._EVAL_70(rsink__EVAL_70),
    ._EVAL_71(rsink__EVAL_71),
    ._EVAL_72(rsink__EVAL_72)
  );
  assign rsink__EVAL_66 = _EVAL_36;
  assign _EVAL_59 = rsink__EVAL_70;
  assign _EVAL_28 = rsink__EVAL_44;
  assign _EVAL_52 = rsink__EVAL_49;
  assign rsink__EVAL_51 = _EVAL_16;
  assign rsink__EVAL_23 = _EVAL_64;
  assign rsink__EVAL_7 = _EVAL_68;
  assign rsink__EVAL_4 = _EVAL_48;
  assign rsink__EVAL_72 = _EVAL_61;
  assign _EVAL_53 = rsink__EVAL_5;
  assign rsink__EVAL_36 = _EVAL_27;
  assign rsink__EVAL_60 = _EVAL_66;
  assign _EVAL_42 = rsink__EVAL_34;
  assign _EVAL_38 = rsink__EVAL_10;
  assign _EVAL_55 = rsink__EVAL_57;
  assign _EVAL_72 = rsink__EVAL_58;
  assign rsink__EVAL_11 = _EVAL_26;
  assign rsink__EVAL_28 = _EVAL_45;
  assign _EVAL_29 = rsink__EVAL_21;
  assign rsink__EVAL_26 = _EVAL_58;
  assign _EVAL_39 = rsink__EVAL_1;
  assign _EVAL_31 = rsink__EVAL_45;
  assign _EVAL_65 = rsink__EVAL_56;
  assign rsink__EVAL_42 = _EVAL_47;
  assign _EVAL_23 = rsink__EVAL_22;
  assign rsink__EVAL_53 = _EVAL_4;
  assign _EVAL_8 = rsink__EVAL_38;
  assign rsink__EVAL_63 = _EVAL_33;
  assign rsink__EVAL_59 = _EVAL_14;
  assign _EVAL_1 = rsink__EVAL_67;
  assign _EVAL_54 = rsink__EVAL_2;
  assign rsink__EVAL_48 = _EVAL_22;
  assign rsink__EVAL_65 = _EVAL_63;
  assign _EVAL_71 = rsink__EVAL_69;
  assign rsink__EVAL_47 = _EVAL_62;
  assign rsink__EVAL_33 = _EVAL_69;
  assign _EVAL_40 = rsink__EVAL_12;
  assign _EVAL_20 = rsink__EVAL_14;
  assign rsink__EVAL_31 = _EVAL_46;
  assign _EVAL_11 = rsink__EVAL_17;
  assign rsink__EVAL = _EVAL_50;
  assign rsink__EVAL_9 = _EVAL_24;
  assign rsink__EVAL_71 = _EVAL;
  assign rsink__EVAL_37 = _EVAL_30;
  assign rsink__EVAL_18 = _EVAL_21;
  assign _EVAL_70 = rsink__EVAL_32;
  assign rsink__EVAL_13 = _EVAL_18;
  assign _EVAL_15 = rsink__EVAL_30;
  assign rsink__EVAL_54 = _EVAL_57;
  assign _EVAL_10 = rsink__EVAL_8;
  assign rsink__EVAL_0 = _EVAL_2;
  assign rsink__EVAL_40 = _EVAL_56;
  assign rsink__EVAL_16 = _EVAL_37;
  assign _EVAL_7 = rsink__EVAL_20;
  assign rsink__EVAL_15 = _EVAL_51;
  assign rsink__EVAL_50 = _EVAL_43;
  assign _EVAL_34 = rsink__EVAL_62;
  assign _EVAL_17 = rsink__EVAL_52;
  assign _EVAL_67 = rsink__EVAL_43;
  assign _EVAL_35 = rsink__EVAL_68;
  assign rsink__EVAL_55 = _EVAL_60;
  assign _EVAL_6 = rsink__EVAL_29;
  assign rsink__EVAL_61 = _EVAL_49;
  assign rsink__EVAL_39 = _EVAL_19;
  assign rsink__EVAL_25 = _EVAL_13;
  assign _EVAL_41 = rsink__EVAL_24;
  assign rsink__EVAL_35 = _EVAL_3;
  assign rsink__EVAL_19 = _EVAL_12;
  assign _EVAL_5 = rsink__EVAL_64;
  assign _EVAL_32 = rsink__EVAL_27;
  assign _EVAL_9 = rsink__EVAL_46;
  assign rsink__EVAL_3 = _EVAL_44;
  assign _EVAL_25 = rsink__EVAL_6;
  assign rsink__EVAL_41 = _EVAL_0;
endmodule
