//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_199(
  output        _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  input         _EVAL_2,
  input         _EVAL_3,
  input  [15:0] _EVAL_4,
  input         _EVAL_5,
  input  [10:0] _EVAL_6,
  input         _EVAL_7,
  input  [3:0]  _EVAL_8
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg  _EVAL_9;
  wire  _EVAL_10;
  reg  _EVAL_12;
  wire  _EVAL_13;
  wire  _EVAL_15;
  wire  _EVAL_17;
  reg  _EVAL_18;
  reg  _EVAL_19;
  reg  _EVAL_20;
  wire  _EVAL_25;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_35;
  reg  _EVAL_36;
  wire  _EVAL_38;
  wire  _EVAL_39;
  reg  _EVAL_40;
  wire  _EVAL_41;
  reg  _EVAL_42;
  reg  _EVAL_43;
  reg  _EVAL_44;
  reg  _EVAL_45;
  wire [31:0] _EVAL_47;
  reg  _EVAL_48;
  reg  _EVAL_50;
  reg  _EVAL_51;
  reg  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_56;
  reg  _EVAL_57;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  reg  _EVAL_63;
  wire  _EVAL_65;
  reg  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_69;
  reg  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  reg  _EVAL_73;
  reg  _EVAL_74;
  reg  _EVAL_76;
  reg  _EVAL_78;
  reg  _EVAL_80;
  wire  _EVAL_81;
  reg  _EVAL_82;
  reg  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  reg  _EVAL_94;
  wire  _EVAL_95;
  reg  _EVAL_97;
  wire  _EVAL_106;
  wire  _EVAL_108;
  reg  _EVAL_110;
  wire  _EVAL_111;
  reg  _EVAL_112;
  wire  _EVAL_115;
  reg  _EVAL_116;
  reg  _EVAL_117;
  assign _EVAL_108 = _EVAL_47[23];
  assign _EVAL_111 = _EVAL_47[13];
  assign _EVAL_88 = _EVAL_47[30];
  assign _EVAL_25 = _EVAL_47[16];
  assign _EVAL_17 = _EVAL_47[0];
  assign _EVAL_67 = _EVAL_47[25];
  assign _EVAL_13 = _EVAL_47[3];
  assign _EVAL_38 = _EVAL_47[7];
  assign _EVAL_47 = {_EVAL_8,_EVAL_4,_EVAL_6,1'h1};
  assign _EVAL_53 = _EVAL_47[28];
  assign _EVAL_28 = _EVAL_47[15];
  assign _EVAL_56 = _EVAL_47[4];
  assign _EVAL = _EVAL_51;
  assign _EVAL_62 = _EVAL_47[11];
  assign _EVAL_60 = _EVAL_47[5];
  assign _EVAL_95 = _EVAL_47[26];
  assign _EVAL_72 = _EVAL_47[27];
  assign _EVAL_65 = _EVAL_47[1];
  assign _EVAL_115 = _EVAL_47[17];
  assign _EVAL_41 = _EVAL_47[20];
  assign _EVAL_90 = _EVAL_47[31];
  assign _EVAL_10 = _EVAL_47[8];
  assign _EVAL_15 = _EVAL_47[10];
  assign _EVAL_85 = _EVAL_47[21];
  assign _EVAL_61 = _EVAL_47[24];
  assign _EVAL_54 = _EVAL_47[12];
  assign _EVAL_29 = _EVAL_47[19];
  assign _EVAL_106 = _EVAL_47[9];
  assign _EVAL_89 = _EVAL_47[14];
  assign _EVAL_39 = _EVAL_47[6];
  assign _EVAL_71 = _EVAL_47[22];
  assign _EVAL_35 = _EVAL_47[18];
  assign _EVAL_81 = _EVAL_47[29];
  assign _EVAL_69 = _EVAL_47[2];
  always @(posedge _EVAL_5) begin
    if (_EVAL_2) begin
      _EVAL_9 <= _EVAL_115;
    end else if (_EVAL_1) begin
      _EVAL_9 <= _EVAL_82;
    end
    if (_EVAL_2) begin
      _EVAL_12 <= _EVAL_53;
    end else if (_EVAL_1) begin
      _EVAL_12 <= _EVAL_94;
    end
    if (_EVAL_2) begin
      _EVAL_18 <= _EVAL_71;
    end else if (_EVAL_1) begin
      _EVAL_18 <= _EVAL_80;
    end
    if (_EVAL_2) begin
      _EVAL_19 <= _EVAL_95;
    end else if (_EVAL_1) begin
      _EVAL_19 <= _EVAL_50;
    end
    if (_EVAL_2) begin
      _EVAL_20 <= _EVAL_38;
    end else if (_EVAL_1) begin
      _EVAL_20 <= _EVAL_36;
    end
    if (_EVAL_2) begin
      _EVAL_36 <= _EVAL_10;
    end else if (_EVAL_1) begin
      _EVAL_36 <= _EVAL_57;
    end
    if (_EVAL_2) begin
      _EVAL_40 <= _EVAL_90;
    end else if (_EVAL_1) begin
      _EVAL_40 <= _EVAL_3;
    end
    if (_EVAL_2) begin
      _EVAL_42 <= _EVAL_61;
    end else if (_EVAL_1) begin
      _EVAL_42 <= _EVAL_45;
    end
    if (_EVAL_2) begin
      _EVAL_43 <= _EVAL_29;
    end else if (_EVAL_1) begin
      _EVAL_43 <= _EVAL_112;
    end
    if (_EVAL_2) begin
      _EVAL_44 <= _EVAL_65;
    end else if (_EVAL_1) begin
      _EVAL_44 <= _EVAL_84;
    end
    if (_EVAL_2) begin
      _EVAL_45 <= _EVAL_67;
    end else if (_EVAL_1) begin
      _EVAL_45 <= _EVAL_19;
    end
    if (_EVAL_2) begin
      _EVAL_48 <= _EVAL_39;
    end else if (_EVAL_1) begin
      _EVAL_48 <= _EVAL_20;
    end
    if (_EVAL_2) begin
      _EVAL_50 <= _EVAL_72;
    end else if (_EVAL_1) begin
      _EVAL_50 <= _EVAL_12;
    end
    if (_EVAL_2) begin
      _EVAL_51 <= _EVAL_17;
    end else if (_EVAL_1) begin
      _EVAL_51 <= _EVAL_44;
    end
    if (_EVAL_2) begin
      _EVAL_52 <= _EVAL_88;
    end else if (_EVAL_1) begin
      _EVAL_52 <= _EVAL_40;
    end
    if (_EVAL_2) begin
      _EVAL_57 <= _EVAL_106;
    end else if (_EVAL_1) begin
      _EVAL_57 <= _EVAL_110;
    end
    if (_EVAL_2) begin
      _EVAL_63 <= _EVAL_25;
    end else if (_EVAL_1) begin
      _EVAL_63 <= _EVAL_9;
    end
    if (_EVAL_2) begin
      _EVAL_66 <= _EVAL_56;
    end else if (_EVAL_1) begin
      _EVAL_66 <= _EVAL_116;
    end
    if (_EVAL_2) begin
      _EVAL_70 <= _EVAL_13;
    end else if (_EVAL_1) begin
      _EVAL_70 <= _EVAL_66;
    end
    if (_EVAL_2) begin
      _EVAL_73 <= _EVAL_62;
    end else if (_EVAL_1) begin
      _EVAL_73 <= _EVAL_76;
    end
    if (_EVAL_2) begin
      _EVAL_74 <= _EVAL_89;
    end else if (_EVAL_1) begin
      _EVAL_74 <= _EVAL_97;
    end
    if (_EVAL_2) begin
      _EVAL_76 <= _EVAL_54;
    end else if (_EVAL_1) begin
      _EVAL_76 <= _EVAL_117;
    end
    if (_EVAL_2) begin
      _EVAL_78 <= _EVAL_85;
    end else if (_EVAL_1) begin
      _EVAL_78 <= _EVAL_18;
    end
    if (_EVAL_2) begin
      _EVAL_80 <= _EVAL_108;
    end else if (_EVAL_1) begin
      _EVAL_80 <= _EVAL_42;
    end
    if (_EVAL_2) begin
      _EVAL_82 <= _EVAL_35;
    end else if (_EVAL_1) begin
      _EVAL_82 <= _EVAL_43;
    end
    if (_EVAL_2) begin
      _EVAL_84 <= _EVAL_69;
    end else if (_EVAL_1) begin
      _EVAL_84 <= _EVAL_70;
    end
    if (_EVAL_2) begin
      _EVAL_94 <= _EVAL_81;
    end else if (_EVAL_1) begin
      _EVAL_94 <= _EVAL_52;
    end
    if (_EVAL_2) begin
      _EVAL_97 <= _EVAL_28;
    end else if (_EVAL_1) begin
      _EVAL_97 <= _EVAL_63;
    end
    if (_EVAL_2) begin
      _EVAL_110 <= _EVAL_15;
    end else if (_EVAL_1) begin
      _EVAL_110 <= _EVAL_73;
    end
    if (_EVAL_2) begin
      _EVAL_112 <= _EVAL_41;
    end else if (_EVAL_1) begin
      _EVAL_112 <= _EVAL_78;
    end
    if (_EVAL_2) begin
      _EVAL_116 <= _EVAL_60;
    end else if (_EVAL_1) begin
      _EVAL_116 <= _EVAL_48;
    end
    if (_EVAL_2) begin
      _EVAL_117 <= _EVAL_111;
    end else if (_EVAL_1) begin
      _EVAL_117 <= _EVAL_74;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_9 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_12 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_18 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_19 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_20 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_36 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_40 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_42 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_43 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_44 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_45 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_48 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_50 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_51 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_52 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_57 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_63 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _EVAL_66 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _EVAL_70 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  _EVAL_73 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  _EVAL_74 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _EVAL_76 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  _EVAL_78 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  _EVAL_80 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  _EVAL_82 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  _EVAL_84 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  _EVAL_94 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  _EVAL_97 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  _EVAL_110 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  _EVAL_112 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  _EVAL_116 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  _EVAL_117 = _RAND_31[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
