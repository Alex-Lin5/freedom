//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_19(
  output [4:0]  _EVAL,
  input  [30:0] _EVAL_0,
  input  [2:0]  _EVAL_1,
  input  [2:0]  _EVAL_2,
  input  [31:0] _EVAL_3,
  output [31:0] _EVAL_4,
  output        _EVAL_5,
  output [2:0]  _EVAL_6,
  output        _EVAL_7,
  output [30:0] _EVAL_8,
  output [2:0]  _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [4:0]  _EVAL_13,
  input  [31:0] _EVAL_14,
  output [2:0]  _EVAL_15,
  output [2:0]  _EVAL_16,
  input         _EVAL_17,
  output        _EVAL_18,
  input  [4:0]  _EVAL_19,
  output        _EVAL_20,
  input         _EVAL_21,
  input         _EVAL_22,
  input         _EVAL_23,
  output        _EVAL_24,
  input  [3:0]  _EVAL_25,
  input         _EVAL_26,
  output        _EVAL_27,
  output [1:0]  _EVAL_28,
  output        _EVAL_29,
  input         _EVAL_30,
  input  [2:0]  _EVAL_31,
  input         _EVAL_32,
  input         _EVAL_33,
  input         _EVAL_34,
  output        _EVAL_35,
  output        _EVAL_36,
  output [4:0]  _EVAL_37,
  output        _EVAL_38,
  input         _EVAL_39,
  input  [1:0]  _EVAL_40,
  input  [2:0]  _EVAL_41,
  output [2:0]  _EVAL_42,
  output [31:0] _EVAL_43,
  output [3:0]  _EVAL_44,
  input         _EVAL_45,
  input         _EVAL_46,
  output        _EVAL_47,
  output        _EVAL_48
);
  wire [30:0] bundleOut_0_a_q__EVAL;
  wire  bundleOut_0_a_q__EVAL_0;
  wire [2:0] bundleOut_0_a_q__EVAL_1;
  wire  bundleOut_0_a_q__EVAL_2;
  wire  bundleOut_0_a_q__EVAL_3;
  wire  bundleOut_0_a_q__EVAL_4;
  wire  bundleOut_0_a_q__EVAL_5;
  wire [31:0] bundleOut_0_a_q__EVAL_6;
  wire  bundleOut_0_a_q__EVAL_7;
  wire [2:0] bundleOut_0_a_q__EVAL_8;
  wire  bundleOut_0_a_q__EVAL_9;
  wire [4:0] bundleOut_0_a_q__EVAL_10;
  wire  bundleOut_0_a_q__EVAL_11;
  wire  bundleOut_0_a_q__EVAL_12;
  wire [3:0] bundleOut_0_a_q__EVAL_13;
  wire [30:0] bundleOut_0_a_q__EVAL_14;
  wire  bundleOut_0_a_q__EVAL_15;
  wire [2:0] bundleOut_0_a_q__EVAL_16;
  wire [31:0] bundleOut_0_a_q__EVAL_17;
  wire [3:0] bundleOut_0_a_q__EVAL_18;
  wire  bundleOut_0_a_q__EVAL_19;
  wire [2:0] bundleOut_0_a_q__EVAL_20;
  wire  bundleOut_0_a_q__EVAL_21;
  wire  bundleOut_0_a_q__EVAL_22;
  wire  bundleOut_0_a_q__EVAL_23;
  wire [2:0] bundleOut_0_a_q__EVAL_24;
  wire [4:0] bundleOut_0_a_q__EVAL_25;
  wire  bundleOut_0_a_q__EVAL_26;
  wire  bundleOut_0_a_q__EVAL_27;
  wire [2:0] bundleOut_0_a_q__EVAL_28;
  wire [31:0] bundleIn_0_d_q__EVAL;
  wire  bundleIn_0_d_q__EVAL_0;
  wire  bundleIn_0_d_q__EVAL_1;
  wire  bundleIn_0_d_q__EVAL_2;
  wire [2:0] bundleIn_0_d_q__EVAL_3;
  wire [4:0] bundleIn_0_d_q__EVAL_4;
  wire  bundleIn_0_d_q__EVAL_5;
  wire  bundleIn_0_d_q__EVAL_6;
  wire  bundleIn_0_d_q__EVAL_7;
  wire  bundleIn_0_d_q__EVAL_8;
  wire [31:0] bundleIn_0_d_q__EVAL_9;
  wire [1:0] bundleIn_0_d_q__EVAL_10;
  wire  bundleIn_0_d_q__EVAL_11;
  wire  bundleIn_0_d_q__EVAL_12;
  wire  bundleIn_0_d_q__EVAL_13;
  wire [2:0] bundleIn_0_d_q__EVAL_14;
  wire [2:0] bundleIn_0_d_q__EVAL_15;
  wire [2:0] bundleIn_0_d_q__EVAL_16;
  wire [4:0] bundleIn_0_d_q__EVAL_17;
  wire  bundleIn_0_d_q__EVAL_18;
  wire  bundleIn_0_d_q__EVAL_19;
  wire [1:0] bundleIn_0_d_q__EVAL_20;
  _EVAL_17 bundleOut_0_a_q (
    ._EVAL(bundleOut_0_a_q__EVAL),
    ._EVAL_0(bundleOut_0_a_q__EVAL_0),
    ._EVAL_1(bundleOut_0_a_q__EVAL_1),
    ._EVAL_2(bundleOut_0_a_q__EVAL_2),
    ._EVAL_3(bundleOut_0_a_q__EVAL_3),
    ._EVAL_4(bundleOut_0_a_q__EVAL_4),
    ._EVAL_5(bundleOut_0_a_q__EVAL_5),
    ._EVAL_6(bundleOut_0_a_q__EVAL_6),
    ._EVAL_7(bundleOut_0_a_q__EVAL_7),
    ._EVAL_8(bundleOut_0_a_q__EVAL_8),
    ._EVAL_9(bundleOut_0_a_q__EVAL_9),
    ._EVAL_10(bundleOut_0_a_q__EVAL_10),
    ._EVAL_11(bundleOut_0_a_q__EVAL_11),
    ._EVAL_12(bundleOut_0_a_q__EVAL_12),
    ._EVAL_13(bundleOut_0_a_q__EVAL_13),
    ._EVAL_14(bundleOut_0_a_q__EVAL_14),
    ._EVAL_15(bundleOut_0_a_q__EVAL_15),
    ._EVAL_16(bundleOut_0_a_q__EVAL_16),
    ._EVAL_17(bundleOut_0_a_q__EVAL_17),
    ._EVAL_18(bundleOut_0_a_q__EVAL_18),
    ._EVAL_19(bundleOut_0_a_q__EVAL_19),
    ._EVAL_20(bundleOut_0_a_q__EVAL_20),
    ._EVAL_21(bundleOut_0_a_q__EVAL_21),
    ._EVAL_22(bundleOut_0_a_q__EVAL_22),
    ._EVAL_23(bundleOut_0_a_q__EVAL_23),
    ._EVAL_24(bundleOut_0_a_q__EVAL_24),
    ._EVAL_25(bundleOut_0_a_q__EVAL_25),
    ._EVAL_26(bundleOut_0_a_q__EVAL_26),
    ._EVAL_27(bundleOut_0_a_q__EVAL_27),
    ._EVAL_28(bundleOut_0_a_q__EVAL_28)
  );
  _EVAL_18 bundleIn_0_d_q (
    ._EVAL(bundleIn_0_d_q__EVAL),
    ._EVAL_0(bundleIn_0_d_q__EVAL_0),
    ._EVAL_1(bundleIn_0_d_q__EVAL_1),
    ._EVAL_2(bundleIn_0_d_q__EVAL_2),
    ._EVAL_3(bundleIn_0_d_q__EVAL_3),
    ._EVAL_4(bundleIn_0_d_q__EVAL_4),
    ._EVAL_5(bundleIn_0_d_q__EVAL_5),
    ._EVAL_6(bundleIn_0_d_q__EVAL_6),
    ._EVAL_7(bundleIn_0_d_q__EVAL_7),
    ._EVAL_8(bundleIn_0_d_q__EVAL_8),
    ._EVAL_9(bundleIn_0_d_q__EVAL_9),
    ._EVAL_10(bundleIn_0_d_q__EVAL_10),
    ._EVAL_11(bundleIn_0_d_q__EVAL_11),
    ._EVAL_12(bundleIn_0_d_q__EVAL_12),
    ._EVAL_13(bundleIn_0_d_q__EVAL_13),
    ._EVAL_14(bundleIn_0_d_q__EVAL_14),
    ._EVAL_15(bundleIn_0_d_q__EVAL_15),
    ._EVAL_16(bundleIn_0_d_q__EVAL_16),
    ._EVAL_17(bundleIn_0_d_q__EVAL_17),
    ._EVAL_18(bundleIn_0_d_q__EVAL_18),
    ._EVAL_19(bundleIn_0_d_q__EVAL_19),
    ._EVAL_20(bundleIn_0_d_q__EVAL_20)
  );
  assign bundleOut_0_a_q__EVAL_22 = _EVAL_23;
  assign bundleIn_0_d_q__EVAL_4 = _EVAL_13;
  assign _EVAL_4 = bundleOut_0_a_q__EVAL_6;
  assign _EVAL_43 = bundleIn_0_d_q__EVAL_9;
  assign _EVAL_8 = bundleOut_0_a_q__EVAL_14;
  assign _EVAL_6 = bundleIn_0_d_q__EVAL_16;
  assign _EVAL_9 = bundleIn_0_d_q__EVAL_3;
  assign _EVAL_35 = bundleOut_0_a_q__EVAL_27;
  assign bundleOut_0_a_q__EVAL_19 = _EVAL_45;
  assign _EVAL = bundleIn_0_d_q__EVAL_17;
  assign _EVAL_28 = bundleIn_0_d_q__EVAL_20;
  assign bundleOut_0_a_q__EVAL_1 = _EVAL_2;
  assign bundleOut_0_a_q__EVAL_5 = _EVAL_32;
  assign bundleOut_0_a_q__EVAL_11 = _EVAL_46;
  assign bundleOut_0_a_q__EVAL_12 = _EVAL_10;
  assign bundleIn_0_d_q__EVAL = _EVAL_14;
  assign bundleIn_0_d_q__EVAL_0 = _EVAL_34;
  assign bundleOut_0_a_q__EVAL_18 = _EVAL_25;
  assign bundleOut_0_a_q__EVAL_20 = _EVAL_1;
  assign _EVAL_15 = bundleOut_0_a_q__EVAL_16;
  assign bundleOut_0_a_q__EVAL_23 = _EVAL_22;
  assign bundleOut_0_a_q__EVAL_17 = _EVAL_3;
  assign bundleOut_0_a_q__EVAL_0 = _EVAL_21;
  assign bundleIn_0_d_q__EVAL_12 = _EVAL_30;
  assign _EVAL_16 = bundleOut_0_a_q__EVAL_24;
  assign _EVAL_7 = bundleIn_0_d_q__EVAL_7;
  assign bundleOut_0_a_q__EVAL_7 = _EVAL_11;
  assign _EVAL_36 = bundleIn_0_d_q__EVAL_19;
  assign _EVAL_5 = bundleOut_0_a_q__EVAL_9;
  assign bundleOut_0_a_q__EVAL_10 = _EVAL_19;
  assign bundleIn_0_d_q__EVAL_15 = _EVAL_12;
  assign bundleOut_0_a_q__EVAL_3 = _EVAL_39;
  assign _EVAL_44 = bundleOut_0_a_q__EVAL_13;
  assign bundleOut_0_a_q__EVAL_28 = _EVAL_41;
  assign _EVAL_20 = bundleIn_0_d_q__EVAL_13;
  assign bundleIn_0_d_q__EVAL_5 = _EVAL_22;
  assign bundleIn_0_d_q__EVAL_10 = _EVAL_40;
  assign bundleIn_0_d_q__EVAL_2 = _EVAL_17;
  assign bundleIn_0_d_q__EVAL_1 = _EVAL_46;
  assign bundleIn_0_d_q__EVAL_14 = _EVAL_31;
  assign bundleOut_0_a_q__EVAL = _EVAL_0;
  assign _EVAL_48 = bundleOut_0_a_q__EVAL_21;
  assign _EVAL_42 = bundleOut_0_a_q__EVAL_8;
  assign _EVAL_47 = bundleIn_0_d_q__EVAL_11;
  assign _EVAL_27 = bundleIn_0_d_q__EVAL_8;
  assign _EVAL_37 = bundleOut_0_a_q__EVAL_25;
  assign _EVAL_29 = bundleOut_0_a_q__EVAL_15;
  assign bundleIn_0_d_q__EVAL_6 = _EVAL_26;
  assign _EVAL_38 = bundleOut_0_a_q__EVAL_4;
  assign _EVAL_18 = bundleOut_0_a_q__EVAL_26;
  assign bundleIn_0_d_q__EVAL_18 = _EVAL_33;
  assign _EVAL_24 = bundleOut_0_a_q__EVAL_2;
endmodule
