//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_43_assert(
  input  [3:0]  _EVAL,
  input  [4:0]  _EVAL_0,
  input  [2:0]  _EVAL_1,
  input  [2:0]  _EVAL_2,
  input         _EVAL_3,
  input  [4:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  input  [3:0]  _EVAL_7,
  input  [2:0]  _EVAL_8,
  input         _EVAL_9,
  input  [1:0]  _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input  [3:0]  _EVAL_13,
  input         _EVAL_14,
  input  [31:0] _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire  _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire [32:0] _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire [32:0] _EVAL_34;
  wire  _EVAL_35;
  wire [31:0] _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  reg [5:0] _EVAL_39;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire [1:0] _EVAL_45;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  reg [1:0] _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire [17:0] _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire [17:0] _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire [31:0] _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire [22:0] _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire [5:0] _EVAL_94;
  wire  _EVAL_95;
  reg [5:0] _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire [32:0] _EVAL_99;
  reg [5:0] _EVAL_100;
  wire  _EVAL_101;
  wire [1:0] _EVAL_102;
  wire [31:0] _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire [31:0] _EVAL_112;
  wire  _EVAL_113;
  wire [32:0] _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire [17:0] _EVAL_122;
  wire  _EVAL_123;
  wire [31:0] _EVAL_124;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  reg [4:0] _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire [17:0] _EVAL_132;
  wire  _EVAL_133;
  wire [3:0] _EVAL_134;
  wire [32:0] _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  reg [3:0] _EVAL_138;
  wire  _EVAL_139;
  wire [32:0] _EVAL_140;
  wire  _EVAL_141;
  wire [17:0] _EVAL_142;
  wire  _EVAL_143;
  wire [7:0] _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire [5:0] _EVAL_149;
  wire [32:0] _EVAL_150;
  wire  _EVAL_151;
  wire [32:0] _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  reg [2:0] _EVAL_158;
  wire  _EVAL_160;
  wire [31:0] _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire [32:0] _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire [32:0] _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire [32:0] _EVAL_186;
  wire  _EVAL_187;
  wire [32:0] _EVAL_188;
  wire [3:0] _EVAL_189;
  wire [6:0] _EVAL_190;
  wire [31:0] _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  reg [31:0] _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire [7:0] _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire [7:0] _EVAL_211;
  wire [32:0] _EVAL_212;
  wire [31:0] _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire [17:0] _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire [1:0] _EVAL_219;
  wire  _EVAL_220;
  wire [3:0] _EVAL_221;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire [2:0] _EVAL_225;
  wire [6:0] _EVAL_226;
  wire [22:0] _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire [31:0] _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  wire [32:0] _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire [5:0] _EVAL_244;
  wire [17:0] _EVAL_245;
  wire [32:0] _EVAL_246;
  wire  _EVAL_247;
  reg [2:0] _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire [32:0] _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire [31:0] _EVAL_265;
  wire  _EVAL_266;
  wire [32:0] _EVAL_267;
  wire [31:0] _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  reg  _EVAL_273;
  wire  _EVAL_274;
  wire [32:0] _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  reg  _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire [32:0] _EVAL_283;
  wire  _EVAL_284;
  wire [32:0] _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire [31:0] _EVAL_291;
  wire  _EVAL_292;
  reg [17:0] _EVAL_293;
  wire  _EVAL_294;
  wire  _EVAL_295;
  reg [3:0] _EVAL_296;
  wire  _EVAL_297;
  reg [4:0] _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire [6:0] _EVAL_301;
  wire [17:0] _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_307;
  wire  _EVAL_308;
  wire [31:0] plusarg_reader_out;
  wire [1:0] _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire  _EVAL_314;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_317;
  wire  _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_320;
  wire  _EVAL_321;
  wire  _EVAL_322;
  wire [3:0] _EVAL_323;
  wire  _EVAL_324;
  reg [2:0] _EVAL_325;
  wire  _EVAL_326;
  wire  _EVAL_327;
  wire  _EVAL_328;
  wire  _EVAL_329;
  wire  _EVAL_330;
  wire  _EVAL_331;
  wire  _EVAL_332;
  wire  _EVAL_333;
  wire  _EVAL_334;
  wire [6:0] _EVAL_335;
  wire  _EVAL_336;
  wire  _EVAL_337;
  wire  _EVAL_338;
  wire  _EVAL_339;
  wire  _EVAL_340;
  wire  _EVAL_341;
  wire  _EVAL_342;
  wire  _EVAL_343;
  wire [2:0] _EVAL_344;
  wire  _EVAL_345;
  wire  _EVAL_346;
  wire  _EVAL_347;
  wire  _EVAL_348;
  wire  _EVAL_349;
  reg [31:0] _EVAL_350;
  wire [5:0] _EVAL_351;
  wire [5:0] _EVAL_352;
  wire  _EVAL_353;
  wire [7:0] _EVAL_354;
  wire  _EVAL_355;
  wire [32:0] _EVAL_356;
  wire  _EVAL_357;
  wire  _EVAL_358;
  wire [5:0] _EVAL_359;
  wire  _EVAL_360;
  wire  _EVAL_361;
  reg [5:0] _EVAL_362;
  wire [32:0] _EVAL_363;
  wire [31:0] _EVAL_364;
  wire  _EVAL_365;
  wire  _EVAL_366;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_311 = _EVAL_0[4:3];
  assign _EVAL_124 = _EVAL_15 & _EVAL_236;
  assign _EVAL_104 = _EVAL_18 & _EVAL_44;
  assign _EVAL_264 = _EVAL_51 & _EVAL_332;
  assign _EVAL_180 = _EVAL_318 & _EVAL_88;
  assign _EVAL_213 = 32'h1 << _EVAL_0;
  assign _EVAL_219 = _EVAL_4[4:3];
  assign _EVAL_155 = _EVAL_124 == 32'h0;
  assign _EVAL_150 = {1'b0,$signed(_EVAL_15)};
  assign _EVAL_166 = {1'b0,$signed(_EVAL_112)};
  assign _EVAL_331 = _EVAL == _EVAL_138;
  assign _EVAL_86 = _EVAL_0 == 5'h10;
  assign _EVAL_141 = _EVAL_206 & _EVAL_168;
  assign _EVAL_329 = _EVAL_239 | _EVAL_6;
  assign _EVAL_246 = $signed(_EVAL_356) & -33'sh400000;
  assign _EVAL_123 = _EVAL_8 == 3'h5;
  assign _EVAL_109 = ~_EVAL_126;
  assign _EVAL_156 = _EVAL_4 == 5'h11;
  assign _EVAL_36 = _EVAL_15 ^ 32'h20000000;
  assign _EVAL_102 = 2'h1 << _EVAL_257;
  assign _EVAL_177 = _EVAL_8 == 3'h4;
  assign _EVAL_49 = _EVAL >= 4'h2;
  assign _EVAL_319 = ~_EVAL_151;
  assign _EVAL_115 = $signed(_EVAL_212) == 33'sh0;
  assign _EVAL_151 = _EVAL_2[2];
  assign _EVAL_75 = ~_EVAL_6;
  assign _EVAL_307 = _EVAL_247 | _EVAL_6;
  assign _EVAL_230 = _EVAL_18 & _EVAL_249;
  assign _EVAL_95 = _EVAL_167 | _EVAL_348;
  assign _EVAL_143 = _EVAL_269 | _EVAL_26;
  assign _EVAL_317 = _EVAL_49 | _EVAL_6;
  assign _EVAL_184 = ~_EVAL_179;
  assign _EVAL_245 = _EVAL_293 >> _EVAL_0;
  assign _EVAL_139 = _EVAL_2 == 3'h6;
  assign _EVAL_243 = ~_EVAL_324;
  assign _EVAL_66 = _EVAL_12 & _EVAL_177;
  assign _EVAL_207 = ~_EVAL_127;
  assign _EVAL_281 = _EVAL_142[0];
  assign _EVAL_54 = ~_EVAL_176;
  assign _EVAL_22 = _EVAL_12 & _EVAL_123;
  assign _EVAL_256 = _EVAL_17 == _EVAL_273;
  assign _EVAL_218 = _EVAL_101 | _EVAL_6;
  assign _EVAL_98 = _EVAL_326 | _EVAL_6;
  assign _EVAL_274 = _EVAL_2 == 3'h5;
  assign _EVAL_165 = _EVAL_318 & _EVAL_119;
  assign _EVAL_237 = _EVAL_2 == _EVAL_248;
  assign _EVAL_241 = ~_EVAL_288;
  assign _EVAL_135 = $signed(_EVAL_166) & -33'sh4000;
  assign _EVAL_206 = _EVAL_45[0];
  assign _EVAL_223 = ~_EVAL_17;
  assign _EVAL_27 = _EVAL_2 == 3'h2;
  assign _EVAL_32 = _EVAL_1 <= 3'h1;
  assign _EVAL_301 = _EVAL_362 - 6'h1;
  assign _EVAL_286 = ~_EVAL_98;
  assign _EVAL_252 = _EVAL_199 | _EVAL_131;
  assign _EVAL_302 = _EVAL_364[17:0];
  assign _EVAL_236 = {{24'd0}, _EVAL_354};
  assign _EVAL_76 = _EVAL_12 & _EVAL_147;
  assign _EVAL_282 = ~_EVAL_194;
  assign _EVAL_271 = _EVAL_277 & _EVAL_328;
  assign _EVAL_35 = 4'h2 == _EVAL;
  assign _EVAL_314 = _EVAL_107 | _EVAL_250;
  assign _EVAL_363 = _EVAL_267;
  assign _EVAL_92 = ~_EVAL_153;
  assign _EVAL_112 = _EVAL_15 ^ 32'h1800000;
  assign _EVAL_345 = ~_EVAL_307;
  assign _EVAL_334 = _EVAL_349 | _EVAL_264;
  assign _EVAL_289 = _EVAL_7 == _EVAL_323;
  assign _EVAL_68 = _EVAL_2 == 3'h1;
  assign _EVAL_266 = _EVAL_145 | _EVAL_6;
  assign _EVAL_231 = _EVAL_10 <= 2'h2;
  assign _EVAL_215 = ~_EVAL_90;
  assign _EVAL_80 = _EVAL_341 ? _EVAL_213 : 32'h0;
  assign _EVAL_261 = _EVAL_152;
  assign _EVAL_321 = _EVAL_4 == 5'h10;
  assign _EVAL_106 = ~_EVAL_276;
  assign _EVAL_147 = _EVAL_8 == 3'h0;
  assign _EVAL_216 = _EVAL_70 & _EVAL_122;
  assign _EVAL_119 = _EVAL_15[0];
  assign _EVAL_48 = _EVAL_1 <= 3'h2;
  assign _EVAL_308 = _EVAL_156 | _EVAL_321;
  assign _EVAL_338 = ~_EVAL_193;
  assign _EVAL_337 = _EVAL_13 >= 4'h2;
  assign _EVAL_214 = _EVAL_1 <= 3'h4;
  assign _EVAL_239 = _EVAL_10 == _EVAL_50;
  assign _EVAL_172 = ~_EVAL_313;
  assign _EVAL_84 = _EVAL_49 | _EVAL_187;
  assign _EVAL_209 = ~_EVAL_366;
  assign _EVAL_347 = $signed(_EVAL_363) == 33'sh0;
  assign _EVAL_33 = _EVAL_157 | _EVAL_6;
  assign _EVAL_169 = ~_EVAL_71;
  assign _EVAL_297 = _EVAL_26 & _EVAL_194;
  assign _EVAL_232 = _EVAL_0 == 5'h11;
  assign _EVAL_85 = _EVAL_223 | _EVAL_9;
  assign _EVAL_114 = {1'b0,$signed(_EVAL_291)};
  assign _EVAL_340 = _EVAL_219 == 2'h0;
  assign _EVAL_154 = _EVAL_224 | _EVAL_6;
  assign _EVAL_174 = _EVAL_238 | _EVAL_6;
  assign _EVAL_67 = _EVAL_18 & _EVAL_274;
  assign _EVAL_128 = 4'h6 == _EVAL;
  assign _EVAL_247 = _EVAL_1 != 3'h0;
  assign _EVAL_222 = _EVAL_53 | _EVAL_294;
  assign _EVAL_168 = _EVAL_116 & _EVAL_119;
  assign _EVAL_90 = _EVAL_245[0];
  assign _EVAL_242 = _EVAL_189 == 4'h0;
  assign _EVAL_57 = _EVAL_16 == _EVAL_279;
  assign _EVAL_280 = _EVAL_51 & _EVAL_95;
  assign _EVAL_234 = _EVAL_350 < plusarg_reader_out;
  assign _EVAL_194 = _EVAL_362 == 6'h0;
  assign _EVAL_196 = _EVAL_311 == 2'h0;
  assign _EVAL_186 = $signed(_EVAL_285) & -33'sh2000;
  assign _EVAL_56 = ~_EVAL_203;
  assign _EVAL_360 = _EVAL_199 & _EVAL_278;
  assign _EVAL_29 = _EVAL_60 | _EVAL_333;
  assign _EVAL_146 = _EVAL_28 | _EVAL_254;
  assign _EVAL_28 = $signed(_EVAL_261) == 33'sh0;
  assign _EVAL_182 = _EVAL_12 & _EVAL_64;
  assign _EVAL_295 = ~_EVAL_357;
  assign _EVAL_164 = _EVAL_334 | _EVAL_6;
  assign _EVAL_224 = _EVAL_134 == 4'h0;
  assign _EVAL_342 = _EVAL_215 | _EVAL_6;
  assign _EVAL_153 = _EVAL_231 | _EVAL_6;
  assign _EVAL_324 = _EVAL_48 | _EVAL_6;
  assign _EVAL_111 = _EVAL_12 & _EVAL_208;
  assign _EVAL_31 = ~_EVAL_229;
  assign _EVAL_37 = _EVAL_272 | _EVAL_6;
  assign _EVAL_131 = _EVAL_128 & _EVAL_77;
  assign _EVAL_170 = ~_EVAL_154;
  assign _EVAL_357 = _EVAL_120 | _EVAL_6;
  assign _EVAL_26 = _EVAL_3 & _EVAL_12;
  assign _EVAL_294 = plusarg_reader_out == 32'h0;
  assign _EVAL_24 = _EVAL_32 | _EVAL_6;
  assign _EVAL_217 = ~_EVAL_327;
  assign _EVAL_226 = _EVAL_39 - 6'h1;
  assign _EVAL_59 = _EVAL_80[17:0];
  assign _EVAL_126 = _EVAL_305 | _EVAL_6;
  assign _EVAL_205 = ~_EVAL_173;
  assign _EVAL_30 = _EVAL_35 & _EVAL_348;
  assign _EVAL_120 = _EVAL_1 == 3'h0;
  assign _EVAL_335 = _EVAL_100 - 6'h1;
  assign _EVAL_326 = _EVAL_13 == _EVAL_296;
  assign _EVAL_221 = ~_EVAL_323;
  assign _EVAL_181 = _EVAL_344 <= 3'h6;
  assign _EVAL_332 = $signed(_EVAL_25) == 33'sh0;
  assign _EVAL_161 = _EVAL_15 ^ 32'hc000000;
  assign _EVAL_292 = _EVAL_4 == 5'h8;
  assign _EVAL_91 = _EVAL_361 & _EVAL_86;
  assign _EVAL_341 = _EVAL_269 & _EVAL_65;
  assign _EVAL_132 = _EVAL_59 | _EVAL_293;
  assign _EVAL_225 = _EVAL_0[2:0];
  assign _EVAL_278 = _EVAL_349 | _EVAL_280;
  assign _EVAL_88 = ~_EVAL_119;
  assign _EVAL_113 = ~_EVAL_270;
  assign _EVAL_52 = _EVAL_18 & _EVAL_27;
  assign _EVAL_152 = $signed(_EVAL_150) & -33'sh5000;
  assign _EVAL_200 = _EVAL_349 | _EVAL_175;
  assign _EVAL_330 = ~_EVAL_174;
  assign _EVAL_211 = ~_EVAL_201;
  assign _EVAL_227 = 23'hff << _EVAL;
  assign _EVAL_315 = _EVAL_214 | _EVAL_6;
  assign _EVAL_107 = _EVAL_49 | _EVAL_183;
  assign _EVAL_55 = _EVAL <= 4'h8;
  assign _EVAL_58 = _EVAL_232 | _EVAL_86;
  assign _EVAL_220 = _EVAL_12 & _EVAL_127;
  assign _EVAL_351 = _EVAL_226[5:0];
  assign _EVAL_201 = _EVAL_89[7:0];
  assign _EVAL_101 = _EVAL_10 != 2'h2;
  assign _EVAL_21 = _EVAL_18 & _EVAL_139;
  assign _EVAL_188 = _EVAL_135;
  assign _EVAL_361 = _EVAL <= 4'hb;
  assign _EVAL_73 = _EVAL_360 | _EVAL_6;
  assign _EVAL_105 = _EVAL_26 & _EVAL_118;
  assign _EVAL_257 = _EVAL[0];
  assign _EVAL_60 = _EVAL_146 | _EVAL_347;
  assign _EVAL_187 = _EVAL_136 & _EVAL_318;
  assign _EVAL_167 = _EVAL_29 | _EVAL_332;
  assign _EVAL_117 = _EVAL_237 | _EVAL_6;
  assign _EVAL_198 = _EVAL_242 | _EVAL_6;
  assign _EVAL_64 = _EVAL_8 == 3'h2;
  assign _EVAL_333 = $signed(_EVAL_240) == 33'sh0;
  assign _EVAL_364 = _EVAL_299 ? _EVAL_191 : 32'h0;
  assign _EVAL_44 = _EVAL_2 == 3'h3;
  assign _EVAL_260 = _EVAL_10 == 2'h0;
  assign _EVAL_38 = _EVAL_18 & _EVAL_162;
  assign _EVAL_353 = _EVAL_35 & _EVAL_259;
  assign _EVAL_118 = _EVAL_96 == 6'h0;
  assign _EVAL_77 = _EVAL_0 == 5'h8;
  assign _EVAL_69 = ~_EVAL_185;
  assign _EVAL_299 = _EVAL_105 & _EVAL_207;
  assign _EVAL_290 = ~_EVAL_121;
  assign _EVAL_25 = _EVAL_186;
  assign _EVAL_71 = _EVAL_63 | _EVAL_6;
  assign _EVAL_272 = _EVAL_222 | _EVAL_234;
  assign _EVAL_134 = _EVAL_7 & _EVAL_221;
  assign _EVAL_61 = ~_EVAL_20;
  assign _EVAL_259 = _EVAL_196 & _EVAL_78;
  assign _EVAL_62 = ~_EVAL_37;
  assign _EVAL_176 = _EVAL_281 | _EVAL_6;
  assign _EVAL_94 = _EVAL_211[7:2];
  assign _EVAL_20 = _EVAL_223 | _EVAL_6;
  assign _EVAL_34 = $signed(_EVAL_275) & -33'sh1000;
  assign _EVAL_108 = _EVAL_116 & _EVAL_88;
  assign _EVAL_144 = _EVAL_227[7:0];
  assign _EVAL_254 = $signed(_EVAL_188) == 33'sh0;
  assign _EVAL_327 = _EVAL_200 | _EVAL_6;
  assign _EVAL_238 = ~_EVAL_9;
  assign _EVAL_291 = _EVAL_15 ^ 32'h2000000;
  assign _EVAL_72 = _EVAL_337 | _EVAL_6;
  assign _EVAL_270 = _EVAL_322 | _EVAL_6;
  assign _EVAL_148 = _EVAL_18 & _EVAL_338;
  assign _EVAL_203 = _EVAL_81 | _EVAL_6;
  assign _EVAL_212 = _EVAL_34;
  assign _EVAL_346 = _EVAL_58 | _EVAL_259;
  assign _EVAL_199 = _EVAL_271 | _EVAL_91;
  assign _EVAL_110 = _EVAL_1 <= 3'h3;
  assign _EVAL_284 = _EVAL_18 & _EVAL_68;
  assign _EVAL_19 = _EVAL_308 | _EVAL_339;
  assign _EVAL_178 = |_EVAL_293;
  assign _EVAL_316 = _EVAL_206 & _EVAL_180;
  assign _EVAL_43 = ~_EVAL_117;
  assign _EVAL_359 = _EVAL_335[5:0];
  assign _EVAL_63 = _EVAL_1 == _EVAL_158;
  assign _EVAL_283 = $signed(_EVAL_99) & -33'sh4000;
  assign _EVAL_303 = _EVAL_346 | _EVAL_77;
  assign _EVAL_197 = _EVAL_206 & _EVAL_165;
  assign _EVAL_192 = ~_EVAL_315;
  assign _EVAL_258 = _EVAL_57 | _EVAL_6;
  assign _EVAL_149 = _EVAL_354[7:2];
  assign _EVAL_358 = ~_EVAL_218;
  assign _EVAL_322 = _EVAL_8 <= 3'h6;
  assign _EVAL_204 = _EVAL_278 | _EVAL_6;
  assign _EVAL_339 = _EVAL_340 & _EVAL_181;
  assign _EVAL_312 = ~_EVAL_304;
  assign _EVAL_189 = ~_EVAL_7;
  assign _EVAL_202 = _EVAL_2 == 3'h7;
  assign _EVAL_277 = _EVAL <= 4'h2;
  assign _EVAL_228 = ~_EVAL_24;
  assign _EVAL_250 = _EVAL_206 & _EVAL_108;
  assign _EVAL_116 = ~_EVAL_318;
  assign _EVAL_93 = _EVAL_0 == _EVAL_298;
  assign _EVAL_175 = _EVAL_51 & _EVAL_251;
  assign _EVAL_79 = _EVAL_233 | _EVAL_30;
  assign _EVAL_305 = _EVAL_353 & _EVAL_79;
  assign _EVAL_288 = _EVAL_289 | _EVAL_6;
  assign _EVAL_179 = _EVAL_93 | _EVAL_6;
  assign _EVAL_285 = {1'b0,$signed(_EVAL_36)};
  assign _EVAL_130 = _EVAL_84 | _EVAL_316;
  assign _EVAL_185 = _EVAL_42 | _EVAL_6;
  assign _EVAL_103 = _EVAL_140[31:0];
  assign _EVAL_162 = _EVAL_2 == 3'h0;
  assign _EVAL_323 = {_EVAL_336,_EVAL_130,_EVAL_87,_EVAL_314};
  assign _EVAL_99 = {1'b0,$signed(_EVAL_268)};
  assign _EVAL_355 = ~_EVAL_73;
  assign _EVAL_133 = _EVAL_8[0];
  assign _EVAL_263 = _EVAL_18 & _EVAL_202;
  assign _EVAL_87 = _EVAL_107 | _EVAL_141;
  assign _EVAL_136 = _EVAL_45[1];
  assign _EVAL_251 = _EVAL_29 | _EVAL_348;
  assign _EVAL_89 = 23'hff << _EVAL_13;
  assign _EVAL_51 = _EVAL <= 4'h6;
  assign _EVAL_23 = ~_EVAL_164;
  assign _EVAL_45 = _EVAL_102 | 2'h1;
  assign _EVAL_313 = _EVAL_260 | _EVAL_6;
  assign _EVAL_171 = _EVAL_283;
  assign _EVAL_183 = _EVAL_136 & _EVAL_116;
  assign _EVAL_269 = _EVAL_11 & _EVAL_18;
  assign _EVAL_142 = _EVAL_132 >> _EVAL_4;
  assign _EVAL_127 = _EVAL_8 == 3'h6;
  assign _EVAL_276 = _EVAL_85 | _EVAL_6;
  assign _EVAL_365 = _EVAL_12 & _EVAL_282;
  assign _EVAL_354 = ~_EVAL_144;
  assign _EVAL_193 = _EVAL_100 == 6'h0;
  assign _EVAL_262 = ~_EVAL_33;
  assign _EVAL_122 = ~_EVAL_302;
  assign _EVAL_275 = {1'b0,$signed(_EVAL_265)};
  assign _EVAL_42 = _EVAL_19 | _EVAL_292;
  assign _EVAL_336 = _EVAL_84 | _EVAL_197;
  assign _EVAL_140 = _EVAL_350 + 32'h1;
  assign _EVAL_348 = $signed(_EVAL_171) == 33'sh0;
  assign _EVAL_173 = _EVAL_110 | _EVAL_6;
  assign _EVAL_160 = ~_EVAL_163;
  assign _EVAL_352 = _EVAL_190[5:0];
  assign _EVAL_235 = ~_EVAL_266;
  assign _EVAL_349 = _EVAL_55 & _EVAL_115;
  assign _EVAL_356 = {1'b0,$signed(_EVAL_161)};
  assign _EVAL_65 = _EVAL_39 == 6'h0;
  assign _EVAL_255 = _EVAL_269 & _EVAL_193;
  assign _EVAL_320 = ~_EVAL_14;
  assign _EVAL_137 = ~_EVAL_72;
  assign _EVAL_343 = ~_EVAL_198;
  assign _EVAL_163 = _EVAL_331 | _EVAL_6;
  assign _EVAL_145 = _EVAL_15 == _EVAL_195;
  assign _EVAL_53 = ~_EVAL_178;
  assign _EVAL_268 = _EVAL_15 ^ 32'h80000000;
  assign _EVAL_70 = _EVAL_293 | _EVAL_59;
  assign _EVAL_267 = $signed(_EVAL_114) & -33'sh10000;
  assign _EVAL_287 = _EVAL_155 | _EVAL_6;
  assign _EVAL_47 = ~_EVAL_317;
  assign _EVAL_304 = _EVAL_303 | _EVAL_6;
  assign _EVAL_208 = _EVAL_8 == 3'h1;
  assign _EVAL_249 = _EVAL_2 == 3'h4;
  assign _EVAL_78 = _EVAL_225 <= 3'h6;
  assign _EVAL_240 = _EVAL_246;
  assign _EVAL_253 = ~_EVAL_258;
  assign _EVAL_81 = _EVAL_8 == _EVAL_325;
  assign _EVAL_300 = ~_EVAL_329;
  assign _EVAL_244 = _EVAL_301[5:0];
  assign _EVAL_233 = _EVAL_277 & _EVAL_115;
  assign _EVAL_191 = 32'h1 << _EVAL_4;
  assign _EVAL_265 = _EVAL_15 ^ 32'h3000;
  assign _EVAL_190 = _EVAL_96 - 6'h1;
  assign _EVAL_83 = ~_EVAL_287;
  assign _EVAL_328 = _EVAL_232 | _EVAL_259;
  assign _EVAL_344 = _EVAL_4[2:0];
  assign _EVAL_157 = _EVAL_4 == _EVAL_129;
  assign _EVAL_121 = _EVAL_320 | _EVAL_6;
  assign _EVAL_229 = _EVAL_252 | _EVAL_6;
  assign _EVAL_366 = _EVAL_256 | _EVAL_6;
  assign _EVAL_97 = ~_EVAL_204;
  assign _EVAL_41 = ~_EVAL_342;
  assign _EVAL_318 = _EVAL_15[1];
  always @(posedge _EVAL_5) begin
    if (_EVAL_6) begin
      _EVAL_39 <= 6'h0;
    end else if (_EVAL_269) begin
      if (_EVAL_65) begin
        if (_EVAL_319) begin
          _EVAL_39 <= _EVAL_149;
        end else begin
          _EVAL_39 <= 6'h0;
        end
      end else begin
        _EVAL_39 <= _EVAL_351;
      end
    end
    if (_EVAL_297) begin
      _EVAL_50 <= _EVAL_10;
    end
    if (_EVAL_6) begin
      _EVAL_96 <= 6'h0;
    end else if (_EVAL_26) begin
      if (_EVAL_118) begin
        if (_EVAL_133) begin
          _EVAL_96 <= _EVAL_94;
        end else begin
          _EVAL_96 <= 6'h0;
        end
      end else begin
        _EVAL_96 <= _EVAL_352;
      end
    end
    if (_EVAL_6) begin
      _EVAL_100 <= 6'h0;
    end else if (_EVAL_269) begin
      if (_EVAL_193) begin
        if (_EVAL_319) begin
          _EVAL_100 <= _EVAL_149;
        end else begin
          _EVAL_100 <= 6'h0;
        end
      end else begin
        _EVAL_100 <= _EVAL_359;
      end
    end
    if (_EVAL_297) begin
      _EVAL_129 <= _EVAL_4;
    end
    if (_EVAL_255) begin
      _EVAL_138 <= _EVAL;
    end
    if (_EVAL_255) begin
      _EVAL_158 <= _EVAL_1;
    end
    if (_EVAL_255) begin
      _EVAL_195 <= _EVAL_15;
    end
    if (_EVAL_255) begin
      _EVAL_248 <= _EVAL_2;
    end
    if (_EVAL_297) begin
      _EVAL_273 <= _EVAL_17;
    end
    if (_EVAL_297) begin
      _EVAL_279 <= _EVAL_16;
    end
    if (_EVAL_6) begin
      _EVAL_293 <= 18'h0;
    end else begin
      _EVAL_293 <= _EVAL_216;
    end
    if (_EVAL_297) begin
      _EVAL_296 <= _EVAL_13;
    end
    if (_EVAL_255) begin
      _EVAL_298 <= _EVAL_0;
    end
    if (_EVAL_297) begin
      _EVAL_325 <= _EVAL_8;
    end
    if (_EVAL_6) begin
      _EVAL_350 <= 32'h0;
    end else if (_EVAL_143) begin
      _EVAL_350 <= 32'h0;
    end else begin
      _EVAL_350 <= _EVAL_103;
    end
    if (_EVAL_6) begin
      _EVAL_362 <= 6'h0;
    end else if (_EVAL_26) begin
      if (_EVAL_194) begin
        if (_EVAL_133) begin
          _EVAL_362 <= _EVAL_94;
        end else begin
          _EVAL_362 <= 6'h0;
        end
      end else begin
        _EVAL_362 <= _EVAL_244;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_300) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f36715f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5c11f1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_235) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_358) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3f6b67a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_253) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c45d15f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(144d3671)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_61) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd11a5d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70d71475)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_228) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc39cf25)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_330) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0eea111)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2178656)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_286) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b85b216)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_341 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(539d57c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_286) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ba33b54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c68677)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bac49b5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_330) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96f8d36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c02dfb4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_62) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f5402de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_62) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61113991)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_184) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb4dabad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8679806b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11c3fdd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_205) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbef639a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d3252fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5bb123d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_235) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67136739)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_12 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19170e96)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_330) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1dcc2daa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_12 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99756db3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_192) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9542730)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_341 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_358) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_355) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_169) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d48272)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_299 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(197db3d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e5e7d7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bbbd4638)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(877ce92a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8f59948)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a14925b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_31) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_330) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_358) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76209f63)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(327ad5b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_109) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_137) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3cb5bb31)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8dad8378)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_106) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a14925b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(720e3aab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bb5ca69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_343) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_23) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85c30015)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_92) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a64bfbf6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_217) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88ea01f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_243) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_31) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e1f4f7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_343) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f37c4934)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20900a40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3106f0d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_355) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1c123e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f5cf68f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_172) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(519578c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_217) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7a4d1fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_343) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e204b9d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_228) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13f34650)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_192) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_172) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6c11525)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_343) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_330) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6aa35856)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_295) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8192c660)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_92) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a4df57a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a043f288)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3444c489)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_243) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca0f5cda)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_358) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c7f7dfa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_137) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_69) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1b8884e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34c5eb3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_330) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4075fce7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5d0d660)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_76 & _EVAL_330) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3e49092)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e63cafe9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_345) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(262e2a8a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_111 & _EVAL_106) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c459cce3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_97) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_300) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b17b74c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ae7365b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a5e5ddd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a5260ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_97) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7ee962b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe611b07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_230 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_66 & _EVAL_69) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ba52862)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_312) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c95b9703)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eab85a60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_253) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a107253)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_330) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_184) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba9f60b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd630046)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_365 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4fda11b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_169) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_205) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_75) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a1efc12)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64547168)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ccd75c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_263 & _EVAL_345) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_22 & _EVAL_75) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80379e92)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_220 & _EVAL_61) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efa6cc29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_38 & _EVAL_312) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_148 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(450f4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_67 & _EVAL_23) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_21 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_109) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3cdda38d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_39 = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_50 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_96 = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_100 = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_129 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_138 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_158 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_195 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_248 = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_273 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_279 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_293 = _RAND_11[17:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_296 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_298 = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_325 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_350 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_362 = _RAND_16[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
