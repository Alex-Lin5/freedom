//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_52(
  output [2:0]  _EVAL,
  input  [2:0]  _EVAL_0,
  output        _EVAL_1,
  input  [4:0]  _EVAL_2,
  output [1:0]  _EVAL_3,
  input         _EVAL_4,
  input  [4:0]  _EVAL_5,
  input  [3:0]  _EVAL_6,
  output        _EVAL_7,
  input         _EVAL_8,
  input  [31:0] _EVAL_9,
  output [31:0] _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  output [2:0]  _EVAL_13,
  output [2:0]  _EVAL_14,
  output        _EVAL_15,
  input         _EVAL_16,
  output        _EVAL_17,
  input  [2:0]  _EVAL_18,
  output        _EVAL_19,
  output        _EVAL_20,
  output        _EVAL_21,
  output [3:0]  _EVAL_22,
  output [31:0] _EVAL_23,
  input         _EVAL_24,
  input  [31:0] _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  input  [1:0]  _EVAL_28,
  output [4:0]  _EVAL_29,
  output [3:0]  _EVAL_30,
  input         _EVAL_31,
  output [3:0]  _EVAL_32,
  input         _EVAL_33,
  input         _EVAL_34,
  input         _EVAL_35,
  input  [31:0] _EVAL_36,
  output [4:0]  _EVAL_37,
  output        _EVAL_38,
  output        _EVAL_39,
  input         _EVAL_40,
  output [31:0] _EVAL_41,
  output        _EVAL_42,
  output        _EVAL_43,
  input         _EVAL_44,
  input  [3:0]  _EVAL_45,
  input  [3:0]  _EVAL_46,
  output        _EVAL_47,
  input         _EVAL_48
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire [3:0] _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire [2:0] _EVAL_60;
  wire [1:0] _EVAL_61;
  reg [2:0] _EVAL_62;
  wire [7:0] _EVAL_63;
  wire [22:0] _EVAL_64;
  wire [2:0] _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire [1:0] _EVAL_68;
  wire [3:0] _EVAL_69;
  wire  _EVAL_70;
  wire [5:0] _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire [1:0] _EVAL_77;
  wire [3:0] _EVAL_79;
  reg  _EVAL_80;
  wire [3:0] _EVAL_81;
  wire [3:0] _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire [5:0] _EVAL_85;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire [4:0] _EVAL_89;
  wire  _EVAL_90;
  wire [3:0] _EVAL_91;
  wire [32:0] _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_96;
  reg [3:0] _EVAL_97;
  wire [3:0] _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire [7:0] _EVAL_101;
  wire  _EVAL_103;
  wire [31:0] _EVAL_104;
  wire [1:0] _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire [3:0] _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  reg [3:0] _EVAL_112;
  wire  _EVAL_113;
  wire [5:0] _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire [1:0] _EVAL_117;
  wire  _EVAL_118;
  wire [31:0] _EVAL_119;
  wire [3:0] _EVAL_120;
  wire [32:0] _EVAL_121;
  wire  _EVAL_122;
  wire [32:0] _EVAL_123;
  wire [1:0] _EVAL_124;
  wire [3:0] _EVAL_126;
  wire [3:0] _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  reg  _EVAL_133;
  wire [32:0] _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire [4:0] _EVAL_139;
  wire  _EVAL_140;
  reg [4:0] _EVAL_141;
  wire  _EVAL_142;
  reg  _EVAL_143;
  wire [1:0] _EVAL_144;
  wire  _EVAL_145;
  wire [31:0] _EVAL_146;
  wire [3:0] _EVAL_147;
  wire  _EVAL_149;
  wire [3:0] _EVAL_150;
  wire [3:0] _EVAL_151;
  reg  _EVAL_152;
  wire [1:0] _EVAL_153;
  wire [31:0] _EVAL_154;
  wire [7:0] _EVAL_155;
  wire [5:0] _EVAL_156;
  wire  _EVAL_157;
  wire [3:0] _EVAL_158;
  wire [4:0] _EVAL_159;
  wire [3:0] _EVAL_160;
  reg [1:0] _EVAL_161;
  wire  _EVAL_162;
  wire [3:0] _EVAL_163;
  wire  _EVAL_164;
  wire [3:0] _EVAL_165;
  wire [1:0] _EVAL_166;
  wire  _EVAL_167;
  reg  _EVAL_168;
  wire  _EVAL_169;
  wire [3:0] _EVAL_170;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire [31:0] _EVAL_174;
  wire [7:0] _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire [7:0] _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_188;
  wire [31:0] _EVAL_189;
  wire  _EVAL_190;
  reg [31:0] _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire [3:0] _EVAL_195;
  wire  _EVAL_197;
  wire [1:0] _EVAL_199;
  wire  _EVAL_200;
  wire [4:0] _EVAL_201;
  wire  _EVAL_202;
  wire [1:0] _EVAL_203;
  wire  _EVAL_204;
  wire [31:0] _EVAL_205;
  reg [31:0] _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  reg  _EVAL_209;
  wire [1:0] _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire [3:0] _EVAL_213;
  reg [5:0] _EVAL_214;
  wire [3:0] _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire [32:0] _EVAL_222;
  wire  _EVAL_223;
  wire [7:0] _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire [1:0] _EVAL_230;
  wire  _EVAL_231;
  wire [31:0] _EVAL_232;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire [6:0] _EVAL_237;
  reg [5:0] _EVAL_238;
  wire [3:0] _EVAL_239;
  wire [32:0] _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire [7:0] _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire [1:0] _EVAL_247;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire [3:0] _EVAL_252;
  wire [3:0] _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire [3:0] _EVAL_256;
  wire  _EVAL_257;
  reg [3:0] _EVAL_258;
  wire  _EVAL_259;
  wire [3:0] _EVAL_260;
  wire [1:0] _EVAL_261;
  wire [1:0] _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire [3:0] _EVAL_265;
  wire  _EVAL_266;
  wire [3:0] _EVAL_267;
  wire  _EVAL_268;
  wire [31:0] _EVAL_269;
  reg  _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire [3:0] _EVAL_277;
  wire [1:0] _EVAL_278;
  wire  _EVAL_279;
  wire  _EVAL_280;
  wire [3:0] _EVAL_281;
  wire  _EVAL_282;
  wire [3:0] _EVAL_283;
  wire  _EVAL_285;
  wire [3:0] _EVAL_286;
  wire [3:0] _EVAL_288;
  wire [1:0] _EVAL_289;
  wire [5:0] _EVAL_290;
  wire [7:0] _EVAL_291;
  wire [3:0] _EVAL_292;
  wire [3:0] _EVAL_293;
  wire [7:0] _EVAL_294;
  wire [1:0] _EVAL_295;
  wire [31:0] _EVAL_296;
  wire [3:0] _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire [7:0] _EVAL_300;
  wire [1:0] _EVAL_301;
  wire [3:0] _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire [2:0] _EVAL_306;
  wire [3:0] _EVAL_309;
  wire  _EVAL_310;
  wire [3:0] _EVAL_311;
  wire  _EVAL_313;
  wire  _EVAL_314;
  wire [1:0] _EVAL_316;
  wire [1:0] _EVAL_317;
  wire  _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_320;
  wire [3:0] _EVAL_321;
  wire  _EVAL_322;
  wire [31:0] _EVAL_323;
  wire  _EVAL_324;
  wire  _EVAL_325;
  wire [3:0] _EVAL_327;
  wire  _EVAL_328;
  wire  _EVAL_329;
  wire [7:0] _EVAL_330;
  wire  _EVAL_331;
  wire  _EVAL_332;
  wire  _EVAL_333;
  wire [3:0] _EVAL_335;
  wire [3:0] _EVAL_336;
  wire [1:0] _EVAL_337;
  wire  _EVAL_338;
  wire  _EVAL_339;
  wire  _EVAL_340;
  wire [2:0] _EVAL_341;
  wire  _EVAL_342;
  wire [5:0] _EVAL_343;
  wire  _EVAL_344;
  wire [7:0] _EVAL_345;
  wire [7:0] _EVAL_346;
  wire [3:0] _EVAL_347;
  wire  _EVAL_348;
  wire [3:0] _EVAL_349;
  wire [1:0] _EVAL_350;
  wire  _EVAL_351;
  wire  _EVAL_352;
  wire  _EVAL_353;
  wire [7:0] _EVAL_354;
  wire [1:0] _EVAL_355;
  wire  _EVAL_356;
  wire  _EVAL_357;
  wire  _EVAL_358;
  wire  _EVAL_359;
  wire [1:0] _EVAL_360;
  wire [1:0] _EVAL_362;
  wire  _EVAL_363;
  wire  _EVAL_364;
  wire  _EVAL_365;
  wire  _EVAL_366;
  wire  _EVAL_367;
  wire [4:0] _EVAL_368;
  wire  _EVAL_369;
  wire [1:0] _EVAL_370;
  wire [15:0] _EVAL_371;
  wire  _EVAL_372;
  wire  _EVAL_373;
  wire [7:0] _EVAL_374;
  wire  _EVAL_375;
  wire [2:0] _EVAL_376;
  wire  _EVAL_378;
  wire  _EVAL_379;
  wire  _EVAL_380;
  wire  _EVAL_382;
  wire [3:0] _EVAL_383;
  wire  _EVAL_384;
  wire  _EVAL_386;
  wire  _EVAL_387;
  wire  _EVAL_388;
  wire [4:0] _EVAL_389;
  wire [3:0] _EVAL_390;
  wire  _EVAL_391;
  wire [2:0] _EVAL_393;
  wire  _EVAL_394;
  wire  _EVAL_395;
  wire [7:0] _EVAL_396;
  wire  _EVAL_397;
  wire  _EVAL_398;
  wire  _EVAL_399;
  wire  _EVAL_400;
  wire [3:0] _EVAL_401;
  wire  _EVAL_402;
  wire [31:0] _EVAL_403;
  wire  _EVAL_404;
  wire  _EVAL_405;
  wire  _EVAL_406;
  wire [31:0] _EVAL_407;
  wire [1:0] _EVAL_408;
  wire  _EVAL_409;
  wire  _EVAL_410;
  wire [1:0] _EVAL_411;
  wire [3:0] _EVAL_413;
  wire [31:0] _EVAL_414;
  wire  _EVAL_415;
  reg  _EVAL_416;
  wire  _EVAL_417;
  wire  _EVAL_418;
  wire [7:0] _EVAL_419;
  wire [1:0] _EVAL_420;
  wire [22:0] _EVAL_421;
  wire [3:0] _EVAL_422;
  wire [1:0] _EVAL_423;
  wire  _EVAL_424;
  wire  _EVAL_425;
  wire [1:0] _EVAL_426;
  wire  _EVAL_427;
  wire  _EVAL_428;
  wire  _EVAL_429;
  wire  _EVAL_430;
  wire [6:0] _EVAL_431;
  wire  _EVAL_432;
  wire  _EVAL_433;
  wire  _EVAL_434;
  wire  _EVAL_435;
  wire [1:0] _EVAL_436;
  wire [31:0] _EVAL_437;
  wire [1:0] _EVAL_438;
  wire  _EVAL_439;
  wire  _EVAL_440;
  reg [2:0] _EVAL_441;
  wire  _EVAL_442;
  wire [3:0] _EVAL_443;
  wire [1:0] _EVAL_444;
  wire [1:0] _EVAL_445;
  wire  _EVAL_446;
  wire  _EVAL_447;
  wire  _EVAL_448;
  wire  _EVAL_449;
  wire  _EVAL_450;
  wire [31:0] _EVAL_451;
  wire  _EVAL_452;
  wire [1:0] _EVAL_453;
  wire [7:0] _EVAL_454;
  wire [3:0] _EVAL_455;
  wire [1:0] _EVAL_456;
  wire [31:0] _EVAL_457;
  wire [5:0] _EVAL_458;
  wire [31:0] _EVAL_459;
  wire [1:0] _EVAL_460;
  wire  _EVAL_461;
  reg [31:0] _EVAL_462;
  wire [31:0] _EVAL_463;
  wire  _EVAL_464;
  wire [1:0] _EVAL_465;
  wire  _EVAL_466;
  wire  _EVAL_467;
  wire  _EVAL_468;
  wire  _EVAL_470;
  wire  _EVAL_471;
  wire [3:0] _EVAL_472;
  wire [32:0] _EVAL_474;
  wire  _EVAL_475;
  wire  _EVAL_477;
  wire  _EVAL_478;
  wire  _EVAL_479;
  wire [1:0] _EVAL_480;
  wire  _EVAL_481;
  wire  _EVAL_482;
  reg  _EVAL_483;
  wire [1:0] _EVAL_485;
  wire [1:0] _EVAL_486;
  wire  _EVAL_487;
  wire  _EVAL_488;
  wire [3:0] _EVAL_489;
  wire [3:0] _EVAL_490;
  wire  _EVAL_492;
  wire  _EVAL_493;
  wire  _EVAL_494;
  wire [31:0] _EVAL_495;
  wire  _EVAL_496;
  wire  _EVAL_497;
  assign _EVAL_230 = {_EVAL_464,_EVAL_282};
  assign _EVAL_496 = _EVAL_462[5];
  assign _EVAL_373 = _EVAL_462[6];
  assign _EVAL_103 = _EVAL_191[5];
  assign _EVAL_74 = _EVAL_206[0];
  assign _EVAL_82 = _EVAL_97 >> _EVAL_426;
  assign _EVAL_466 = $signed(_EVAL_474) == 33'sh0;
  assign _EVAL_262 = {_EVAL_391,_EVAL_415};
  assign _EVAL_321 = _EVAL_97 >> _EVAL_465;
  assign _EVAL_259 = _EVAL_462[10];
  assign _EVAL_57 = _EVAL_97 >> _EVAL_370;
  assign _EVAL_434 = _EVAL_191[30];
  assign _EVAL_303 = _EVAL_462[25];
  assign _EVAL_70 = _EVAL_18 == 3'h0;
  assign _EVAL_232 = _EVAL_191 & _EVAL_403;
  assign _EVAL_281 = _EVAL_147 | _EVAL_195;
  assign _EVAL_10 = _EVAL_495 | _EVAL_437;
  assign _EVAL_345 = _EVAL_404 ? 8'hff : 8'h0;
  assign _EVAL_75 = _EVAL_462[13];
  assign _EVAL_193 = _EVAL_238 == 6'h0;
  assign _EVAL_442 = _EVAL_189[31];
  assign _EVAL = _EVAL_424 ? _EVAL_376 : 3'h0;
  assign _EVAL_87 = _EVAL_285 & _EVAL_145;
  assign _EVAL_175 = _EVAL_400 ? 8'hff : 8'h0;
  assign _EVAL_453 = {_EVAL_340,_EVAL_475};
  assign _EVAL_446 = _EVAL_191[8];
  assign _EVAL_460 = {_EVAL_435,_EVAL_164};
  assign _EVAL_474 = _EVAL_121;
  assign _EVAL_351 = _EVAL_249 | _EVAL_279;
  assign _EVAL_244 = ~_EVAL_346;
  assign _EVAL_207 = _EVAL_462[31];
  assign _EVAL_269 = {_EVAL_63,_EVAL_396,_EVAL_101,_EVAL_291};
  assign _EVAL_382 = _EVAL_347[0];
  assign _EVAL_66 = _EVAL_191[24];
  assign _EVAL_417 = _EVAL_161 == 2'h0;
  assign _EVAL_145 = _EVAL_492 & _EVAL_109;
  assign _EVAL_118 = _EVAL_253[0];
  assign _EVAL_286 = _EVAL_97 >> _EVAL_68;
  assign _EVAL_60 = {_EVAL_456, 1'h0};
  assign _EVAL_355 = _EVAL_54 ? _EVAL_362 : _EVAL_161;
  assign _EVAL_127 = {{1'd0}, _EVAL_341};
  assign _EVAL_38 = _EVAL_59 | _EVAL_72;
  assign _EVAL_478 = _EVAL_191[26];
  assign _EVAL_197 = _EVAL_34 | _EVAL_397;
  assign _EVAL_472 = ~_EVAL_158;
  assign _EVAL_457 = {_EVAL_382,_EVAL_225,_EVAL_305,_EVAL_122,_EVAL_52,_EVAL_241,_EVAL_217,_EVAL_328,_EVAL_419,_EVAL_371
    };
  assign _EVAL_162 = _EVAL_45 <= 4'h2;
  assign _EVAL_190 = _EVAL_462[28];
  assign _EVAL_289 = {_EVAL_325,_EVAL_488};
  assign _EVAL_14 = _EVAL_424 ? _EVAL_393 : 3'h0;
  assign _EVAL_497 = _EVAL_104[31];
  assign _EVAL_65 = {{1'd0}, _EVAL_485};
  assign _EVAL_256 = _EVAL_443 | _EVAL_349;
  assign _EVAL_117 = _EVAL_278 | 2'h1;
  assign _EVAL_139 = _EVAL_242 ? _EVAL_141 : 5'h0;
  assign _EVAL_467 = _EVAL_494 & _EVAL_384;
  assign _EVAL_285 = _EVAL_117[0];
  assign _EVAL_408 = _EVAL_306[1:0];
  assign _EVAL_186 = _EVAL_286[0];
  assign _EVAL_438 = ~_EVAL_247;
  assign _EVAL_379 = _EVAL_251 ? _EVAL_351 : _EVAL_487;
  assign _EVAL_369 = _EVAL_81[0];
  assign _EVAL_306 = {_EVAL_317, 1'h0};
  assign _EVAL_151 = _EVAL_97 >> _EVAL_423;
  assign _EVAL_246 = _EVAL_161 == 2'h3;
  assign _EVAL_452 = _EVAL_424 & _EVAL_48;
  assign _EVAL_47 = _EVAL_372 | _EVAL_452;
  assign _EVAL_229 = _EVAL_438[1];
  assign _EVAL_401 = _EVAL_97 >> _EVAL_203;
  assign _EVAL_389 = _EVAL_424 ? _EVAL_2 : 5'h0;
  assign _EVAL_394 = $signed(_EVAL_93) == 33'sh0;
  assign _EVAL_413 = _EVAL_97 >> _EVAL_261;
  assign _EVAL_468 = _EVAL_386 ? _EVAL_304 : _EVAL_236;
  assign _EVAL_386 = _EVAL_442 == _EVAL_497;
  assign _EVAL_426 = {_EVAL_402,_EVAL_190};
  assign _EVAL_189 = _EVAL_232 | _EVAL_146;
  assign _EVAL_90 = _EVAL_281[0];
  assign _EVAL_493 = _EVAL_62[0];
  assign _EVAL_309 = ~_EVAL_112;
  assign _EVAL_481 = _EVAL_462[14];
  assign _EVAL_444 = {_EVAL_130,_EVAL_353};
  assign _EVAL_52 = _EVAL_336[0];
  assign _EVAL_439 = _EVAL_441[0];
  assign _EVAL_240 = {1'b0,$signed(_EVAL_174)};
  assign _EVAL_212 = _EVAL_197 & _EVAL_35;
  assign _EVAL_155 = _EVAL_50 ? 8'hff : 8'h0;
  assign _EVAL_319 = 3'h3 == _EVAL_65;
  assign _EVAL_111 = _EVAL_191[6];
  assign _EVAL_77 = {_EVAL_448,_EVAL_481};
  assign _EVAL_114 = _EVAL_244[7:2];
  assign _EVAL_418 = _EVAL_12[2];
  assign _EVAL_407 = _EVAL_424 ? _EVAL_9 : 32'h0;
  assign _EVAL_106 = 3'h1 == _EVAL_65;
  assign _EVAL_372 = _EVAL_242 & _EVAL_152;
  assign _EVAL_436 = _EVAL_461 ? _EVAL_350 : _EVAL_355;
  assign _EVAL_195 = _EVAL_85[3:0];
  assign _EVAL_310 = _EVAL_462[24];
  assign _EVAL_251 = _EVAL_12 == 3'h3;
  assign _EVAL_101 = _EVAL_194 ? 8'hff : 8'h0;
  assign _EVAL_338 = _EVAL_335[0];
  assign _EVAL_402 = _EVAL_191[28];
  assign _EVAL_221 = 3'h0 == _EVAL_65;
  assign _EVAL_76 = _EVAL_401[0];
  assign _EVAL_243 = _EVAL_183 ? _EVAL_229 : _EVAL_483;
  assign _EVAL_368 = {_EVAL_163, 1'h0};
  assign _EVAL_325 = _EVAL_191[4];
  assign _EVAL_433 = _EVAL_490[0];
  assign _EVAL_219 = _EVAL_191[10];
  assign _EVAL_313 = _EVAL_422[0];
  assign _EVAL_91 = {_EVAL_149,_EVAL_84,_EVAL_181,_EVAL_378};
  assign _EVAL_218 = ~_EVAL_418;
  assign _EVAL_181 = _EVAL_280 | _EVAL_116;
  assign _EVAL_486 = {_EVAL_200,_EVAL_207};
  assign _EVAL_421 = 23'hff << _EVAL_6;
  assign _EVAL_72 = _EVAL_424 & _EVAL_33;
  assign _EVAL_147 = _EVAL_163 | _EVAL_213;
  assign _EVAL_288 = _EVAL_97 >> _EVAL_360;
  assign _EVAL_487 = _EVAL_430 ? _EVAL_351 : 1'h1;
  assign _EVAL_210 = {_EVAL_219,_EVAL_259};
  assign _EVAL_177 = _EVAL_462[29];
  assign _EVAL_414 = _EVAL_275 ? _EVAL_191 : _EVAL_462;
  assign _EVAL_445 = {_EVAL_432,_EVAL_202};
  assign _EVAL_293 = _EVAL_239 & _EVAL_472;
  assign _EVAL_342 = _EVAL_191[16];
  assign _EVAL_261 = {_EVAL_172,_EVAL_234};
  assign _EVAL_204 = _EVAL_191[29];
  assign _EVAL_94 = _EVAL_40 & _EVAL_243;
  assign _EVAL_135 = _EVAL_266 | _EVAL_380;
  assign _EVAL_146 = {_EVAL_178,_EVAL_454,_EVAL_155,_EVAL_175};
  assign _EVAL_431 = _EVAL_238 - 6'h1;
  assign _EVAL_290 = _EVAL_354[7:2];
  assign _EVAL_425 = _EVAL_191[19];
  assign _EVAL_344 = _EVAL_191[22];
  assign _EVAL_166 = {_EVAL_342,_EVAL_409};
  assign _EVAL_375 = _EVAL_108[0];
  assign _EVAL_250 = _EVAL_143 | _EVAL_11;
  assign _EVAL_435 = _EVAL_191[23];
  assign _EVAL_390 = _EVAL_97 >> _EVAL_289;
  assign _EVAL_383 = _EVAL_159[3:0];
  assign _EVAL_58 = _EVAL_242 & _EVAL_83;
  assign _EVAL_98 = _EVAL_97 >> _EVAL_420;
  assign _EVAL_264 = _EVAL_483 & _EVAL_329;
  assign _EVAL_299 = _EVAL_191[15];
  assign _EVAL_337 = {_EVAL_110,_EVAL_128};
  assign _EVAL_297 = _EVAL_97 >> _EVAL_445;
  assign _EVAL_356 = _EVAL_170[0];
  assign _EVAL_252 = _EVAL_97 >> _EVAL_444;
  assign _EVAL_384 = _EVAL_161 != 2'h0;
  assign _EVAL_395 = _EVAL_492 & _EVAL_74;
  assign _EVAL_179 = _EVAL_242 & _EVAL_133;
  assign _EVAL_400 = _EVAL_256[0];
  assign _EVAL_239 = {_EVAL_207,_EVAL_164,_EVAL_228,_EVAL_475};
  assign _EVAL_397 = _EVAL_107 & _EVAL_467;
  assign _EVAL_280 = _EVAL_266 | _EVAL_157;
  assign _EVAL_23 = _EVAL_142 ? _EVAL_462 : _EVAL_25;
  assign _EVAL_427 = _EVAL_191[12];
  assign _EVAL_282 = _EVAL_462[20];
  assign _EVAL_296 = _EVAL_36 ^ 32'h2000;
  assign _EVAL_254 = _EVAL_209 | _EVAL_11;
  assign _EVAL_30 = _EVAL_327 | _EVAL_120;
  assign _EVAL_137 = _EVAL_100 | _EVAL_329;
  assign _EVAL_458 = {_EVAL_443, 2'h0};
  assign _EVAL_121 = $signed(_EVAL_123) & 33'shab002000;
  assign _EVAL_185 = _EVAL_455[0];
  assign _EVAL_160 = _EVAL_97 >> _EVAL_262;
  assign _EVAL_93 = _EVAL_222;
  assign _EVAL_228 = _EVAL_462[15];
  assign _EVAL_495 = _EVAL_242 ? _EVAL_206 : 32'h0;
  assign _EVAL_302 = _EVAL_97 >> _EVAL_166;
  assign _EVAL_156 = _EVAL_431[5:0];
  assign _EVAL_410 = _EVAL_246 | _EVAL_100;
  assign _EVAL_318 = _EVAL_252[0];
  assign _EVAL_432 = _EVAL_191[0];
  assign _EVAL_255 = _EVAL_467 & _EVAL_449;
  assign _EVAL_223 = _EVAL_160[0];
  assign _EVAL_327 = _EVAL_242 ? _EVAL_258 : 4'h0;
  assign _EVAL_398 = _EVAL_462[11];
  assign _EVAL_380 = _EVAL_348 & _EVAL_492;
  assign _EVAL_353 = _EVAL_462[18];
  assign _EVAL_128 = _EVAL_462[17];
  assign _EVAL_260 = _EVAL_97 >> _EVAL_77;
  assign _EVAL_378 = _EVAL_280 | _EVAL_73;
  assign _EVAL_454 = _EVAL_406 ? 8'hff : 8'h0;
  assign _EVAL_64 = 23'hff << _EVAL_45;
  assign _EVAL_271 = _EVAL_191[27];
  assign _EVAL_317 = {_EVAL_329,_EVAL_100};
  assign _EVAL_123 = {1'b0,$signed(_EVAL_296)};
  assign _EVAL_279 = _EVAL_274 & _EVAL_394;
  assign _EVAL_107 = _EVAL_193 & _EVAL_449;
  assign _EVAL_63 = _EVAL_333 ? 8'hff : 8'h0;
  assign _EVAL_348 = _EVAL_117[1];
  assign _EVAL_349 = _EVAL_458[3:0];
  assign _EVAL_88 = _EVAL_62[1];
  assign _EVAL_17 = _EVAL_447 | _EVAL_450;
  assign _EVAL_192 = _EVAL_285 & _EVAL_395;
  assign _EVAL_158 = _EVAL_309 | _EVAL_127;
  assign _EVAL_424 = _EVAL_183 ? _EVAL_227 : _EVAL_483;
  assign _EVAL_1 = _EVAL_179 | _EVAL_429;
  assign _EVAL_265 = _EVAL_97 >> _EVAL_124;
  assign _EVAL_263 = _EVAL_462[26];
  assign _EVAL_374 = _EVAL_358 ? 8'hff : 8'h0;
  assign _EVAL_32 = _EVAL_6;
  assign _EVAL_100 = _EVAL_161 == 2'h2;
  assign _EVAL_130 = _EVAL_191[18];
  assign _EVAL_358 = _EVAL_112[1];
  assign _EVAL_391 = _EVAL_191[21];
  assign _EVAL_332 = _EVAL_424 & _EVAL_27;
  assign _EVAL_42 = _EVAL_183 ? _EVAL_137 : _EVAL_220;
  assign _EVAL_300 = _EVAL_421[7:0];
  assign _EVAL_149 = _EVAL_135 | _EVAL_192;
  assign _EVAL_388 = _EVAL_462[27];
  assign _EVAL_464 = _EVAL_191[20];
  assign _EVAL_331 = _EVAL_462[1];
  assign _EVAL_488 = _EVAL_462[4];
  assign _EVAL_470 = _EVAL_438[0];
  assign _EVAL_81 = _EVAL_97 >> _EVAL_230;
  assign _EVAL_316 = {_EVAL_434,_EVAL_184};
  assign _EVAL_339 = _EVAL_191[2];
  assign _EVAL_202 = _EVAL_462[0];
  assign _EVAL_341 = _EVAL_112[3:1];
  assign _EVAL_352 = _EVAL_212 & _EVAL_193;
  assign _EVAL_494 = _EVAL_141 == _EVAL_5;
  assign _EVAL_366 = _EVAL_302[0];
  assign _EVAL_163 = _EVAL_201[3:0];
  assign _EVAL_437 = _EVAL_424 ? _EVAL_36 : 32'h0;
  assign _EVAL_278 = 2'h1 << _EVAL_298;
  assign _EVAL_447 = _EVAL_242 & _EVAL_80;
  assign _EVAL_415 = _EVAL_462[21];
  assign _EVAL_96 = ~_EVAL_397;
  assign _EVAL_294 = _EVAL_357 ? 8'hff : 8'h0;
  assign _EVAL_283 = _EVAL_424 ? _EVAL_46 : 4'h0;
  assign _EVAL_237 = _EVAL_214 - _EVAL_343;
  assign _EVAL_222 = $signed(_EVAL_240) & 33'shab000000;
  assign _EVAL_159 = {_EVAL_277, 1'h0};
  assign _EVAL_247 = _EVAL_60[1:0];
  assign _EVAL_461 = _EVAL_365 & _EVAL_100;
  assign _EVAL_154 = _EVAL_242 ? _EVAL_119 : 32'h0;
  assign _EVAL_142 = _EVAL_322 & _EVAL_467;
  assign _EVAL_479 = _EVAL_270 & _EVAL_100;
  assign _EVAL_477 = ~_EVAL_410;
  assign _EVAL_56 = _EVAL_462[22];
  assign _EVAL_291 = _EVAL_90 ? 8'hff : 8'h0;
  assign _EVAL_231 = _EVAL_390[0];
  assign _EVAL_475 = _EVAL_462[7];
  assign _EVAL_172 = _EVAL_191[9];
  assign _EVAL_41 = _EVAL_154 | _EVAL_407;
  assign _EVAL_119 = _EVAL_439 ? _EVAL_457 : _EVAL_459;
  assign _EVAL_440 = _EVAL_99 & _EVAL_109;
  assign _EVAL_205 = ~_EVAL_104;
  assign _EVAL_73 = _EVAL_285 & _EVAL_440;
  assign _EVAL_443 = _EVAL_383 | _EVAL_267;
  assign _EVAL_249 = _EVAL_162 & _EVAL_466;
  assign _EVAL_323 = _EVAL_182 ? _EVAL_104 : _EVAL_205;
  assign _EVAL_105 = {_EVAL_271,_EVAL_388};
  assign _EVAL_322 = _EVAL_193 & _EVAL_70;
  assign _EVAL_203 = {_EVAL_208,_EVAL_398};
  assign _EVAL_217 = _EVAL_489[0];
  assign _EVAL_157 = _EVAL_348 & _EVAL_99;
  assign _EVAL_430 = _EVAL_12 == 3'h2;
  assign _EVAL_465 = {_EVAL_425,_EVAL_405};
  assign _EVAL_85 = {_EVAL_147, 2'h0};
  assign _EVAL_22 = _EVAL_150 | _EVAL_283;
  assign _EVAL_357 = _EVAL_112[0];
  assign _EVAL_55 = _EVAL_256[3];
  assign _EVAL_266 = _EVAL_258 >= 4'h2;
  assign _EVAL_234 = _EVAL_462[9];
  assign _EVAL_53 = _EVAL_477 & _EVAL_176;
  assign _EVAL_182 = _EVAL_62[2];
  assign _EVAL_350 = _EVAL_100 ? 2'h1 : _EVAL_355;
  assign _EVAL_320 = _EVAL_462[12];
  assign _EVAL_367 = _EVAL_462[2];
  assign _EVAL_3 = _EVAL_28;
  assign _EVAL_144 = {_EVAL_339,_EVAL_367};
  assign _EVAL_406 = _EVAL_256[2];
  assign _EVAL_311 = _EVAL_97 >> _EVAL_61;
  assign _EVAL_324 = _EVAL_288[0];
  assign _EVAL_15 = _EVAL_34 | _EVAL_397;
  assign _EVAL_492 = _EVAL_206[1];
  assign _EVAL_19 = _EVAL_58 | _EVAL_332;
  assign _EVAL_7 = _EVAL_35 & _EVAL_96;
  assign _EVAL_21 = _EVAL_24;
  assign _EVAL_301 = {_EVAL_204,_EVAL_177};
  assign _EVAL_132 = _EVAL_321[0];
  assign _EVAL_236 = _EVAL_88 == _EVAL_442;
  assign _EVAL_411 = {_EVAL_359,_EVAL_169};
  assign _EVAL_365 = _EVAL_40 & _EVAL_257;
  assign _EVAL_485 = _EVAL_0[1:0];
  assign _EVAL_277 = _EVAL_292 & _EVAL_472;
  assign _EVAL_122 = _EVAL_82[0];
  assign _EVAL_165 = _EVAL_97 >> _EVAL_301;
  assign _EVAL_220 = _EVAL_479 | _EVAL_264;
  assign _EVAL_340 = _EVAL_191[7];
  assign _EVAL_140 = _EVAL_413[0];
  assign _EVAL_153 = {_EVAL_446,_EVAL_51};
  assign _EVAL_138 = _EVAL_260[0];
  assign _EVAL_363 = _EVAL_112[2];
  assign _EVAL_482 = _EVAL_183 ? _EVAL_137 : _EVAL_220;
  assign _EVAL_314 = _EVAL_470 & _EVAL_100;
  assign _EVAL_61 = {_EVAL_111,_EVAL_373};
  assign _EVAL_108 = _EVAL_97 >> _EVAL_337;
  assign _EVAL_404 = _EVAL_112[3];
  assign _EVAL_336 = _EVAL_97 >> _EVAL_105;
  assign _EVAL_456 = _EVAL_317 | _EVAL_408;
  assign _EVAL_39 = _EVAL_94 & _EVAL_53;
  assign _EVAL_360 = {_EVAL_427,_EVAL_320};
  assign _EVAL_20 = _EVAL_142 ? _EVAL_254 : _EVAL_31;
  assign _EVAL_370 = {_EVAL_428,_EVAL_75};
  assign _EVAL_13 = _EVAL_142 ? 3'h1 : _EVAL_18;
  assign _EVAL_170 = _EVAL_97 >> _EVAL_411;
  assign _EVAL_54 = _EVAL_173 & _EVAL_131;
  assign _EVAL_245 = _EVAL_99 & _EVAL_74;
  assign _EVAL_126 = _EVAL_97 >> _EVAL_453;
  assign _EVAL_224 = _EVAL_363 ? 8'hff : 8'h0;
  assign _EVAL_268 = _EVAL_151[0];
  assign _EVAL_329 = _EVAL_4 & _EVAL_53;
  assign _EVAL_194 = _EVAL_281[1];
  assign _EVAL_89 = {_EVAL_383, 1'h0};
  assign _EVAL_201 = {_EVAL_293, 1'h0};
  assign _EVAL_275 = _EVAL_493 == _EVAL_468;
  assign _EVAL_115 = _EVAL_191[25];
  assign _EVAL_347 = _EVAL_97 >> _EVAL_486;
  assign _EVAL_354 = ~_EVAL_300;
  assign _EVAL_428 = _EVAL_191[13];
  assign _EVAL_173 = _EVAL_94 & _EVAL_329;
  assign _EVAL_134 = _EVAL_189 + _EVAL_323;
  assign _EVAL_176 = _EVAL_379 | _EVAL_417;
  assign _EVAL_178 = _EVAL_55 ? 8'hff : 8'h0;
  assign _EVAL_208 = _EVAL_191[11];
  assign _EVAL_448 = _EVAL_191[14];
  assign _EVAL_83 = _EVAL_416 | _EVAL_209;
  assign _EVAL_333 = _EVAL_281[3];
  assign _EVAL_364 = _EVAL_451[31];
  assign _EVAL_37 = _EVAL_5;
  assign _EVAL_346 = _EVAL_64[7:0];
  assign _EVAL_480 = {_EVAL_115,_EVAL_303};
  assign _EVAL_68 = {_EVAL_299,_EVAL_228};
  assign _EVAL_124 = {_EVAL_66,_EVAL_310};
  assign _EVAL_51 = _EVAL_462[8];
  assign _EVAL_257 = _EVAL_183 ? _EVAL_470 : _EVAL_270;
  assign _EVAL_305 = _EVAL_165[0];
  assign _EVAL_199 = {_EVAL_471,_EVAL_331};
  assign _EVAL_463 = _EVAL_462 & _EVAL_403;
  assign _EVAL_188 = _EVAL_183 & _EVAL_40;
  assign _EVAL_376 = _EVAL_131 ? 3'h4 : _EVAL_12;
  assign _EVAL_403 = {_EVAL_345,_EVAL_224,_EVAL_374,_EVAL_294};
  assign _EVAL_69 = _EVAL_97 >> _EVAL_316;
  assign _EVAL_409 = _EVAL_462[16];
  assign _EVAL_131 = ~_EVAL_379;
  assign _EVAL_359 = _EVAL_191[3];
  assign _EVAL_459 = _EVAL_182 ? _EVAL_451 : _EVAL_414;
  assign _EVAL_274 = 4'h2 == _EVAL_45;
  assign _EVAL_343 = {{5'd0}, _EVAL_167};
  assign _EVAL_292 = {_EVAL_200,_EVAL_435,_EVAL_299,_EVAL_340};
  assign _EVAL_110 = _EVAL_191[17];
  assign _EVAL_330 = {_EVAL_399,_EVAL_235,_EVAL_185,_EVAL_231,_EVAL_356,_EVAL_338,_EVAL_118,_EVAL_211};
  assign _EVAL_200 = _EVAL_191[31];
  assign _EVAL_29 = _EVAL_139 | _EVAL_389;
  assign _EVAL_429 = _EVAL_424 & _EVAL_16;
  assign _EVAL_396 = _EVAL_67 ? 8'hff : 8'h0;
  assign _EVAL_43 = _EVAL_142 ? _EVAL_250 : _EVAL_11;
  assign _EVAL_393 = _EVAL_131 ? 3'h0 : _EVAL_0;
  assign _EVAL_184 = _EVAL_462[30];
  assign _EVAL_211 = _EVAL_297[0];
  assign _EVAL_489 = _EVAL_97 >> _EVAL_480;
  assign _EVAL_328 = _EVAL_265[0];
  assign _EVAL_490 = _EVAL_97 >> _EVAL_210;
  assign _EVAL_405 = _EVAL_462[19];
  assign _EVAL_362 = _EVAL_417 ? 2'h3 : _EVAL_161;
  assign _EVAL_71 = _EVAL_237[5:0];
  assign _EVAL_183 = _EVAL_214 == 6'h0;
  assign _EVAL_104 = _EVAL_463 | _EVAL_269;
  assign _EVAL_169 = _EVAL_462[3];
  assign _EVAL_174 = _EVAL_36 ^ 32'h80000000;
  assign _EVAL_99 = ~_EVAL_492;
  assign _EVAL_120 = _EVAL_424 ? _EVAL_45 : 4'h0;
  assign _EVAL_298 = _EVAL_258[0];
  assign _EVAL_164 = _EVAL_462[23];
  assign _EVAL_79 = _EVAL_97 >> _EVAL_460;
  assign _EVAL_399 = _EVAL_126[0];
  assign _EVAL_150 = _EVAL_242 ? _EVAL_91 : 4'h0;
  assign _EVAL_113 = _EVAL_79[0];
  assign _EVAL_371 = {_EVAL_186,_EVAL_138,_EVAL_248,_EVAL_324,_EVAL_76,_EVAL_433,_EVAL_140,_EVAL_313,_EVAL_330};
  assign _EVAL_167 = _EVAL_40 & _EVAL_482;
  assign _EVAL_59 = _EVAL_242 & _EVAL_168;
  assign _EVAL_419 = {_EVAL_113,_EVAL_268,_EVAL_223,_EVAL_369,_EVAL_132,_EVAL_318,_EVAL_375,_EVAL_366};
  assign _EVAL_253 = _EVAL_97 >> _EVAL_199;
  assign _EVAL_50 = _EVAL_256[1];
  assign _EVAL_242 = _EVAL_183 ? _EVAL_314 : _EVAL_270;
  assign _EVAL_455 = _EVAL_97 >> _EVAL_295;
  assign _EVAL_267 = _EVAL_89[3:0];
  assign _EVAL_451 = _EVAL_134[31:0];
  assign _EVAL_449 = _EVAL_18 == 3'h1;
  assign _EVAL_335 = _EVAL_97 >> _EVAL_144;
  assign _EVAL_213 = _EVAL_368[3:0];
  assign _EVAL_422 = _EVAL_97 >> _EVAL_153;
  assign _EVAL_116 = _EVAL_285 & _EVAL_245;
  assign _EVAL_295 = {_EVAL_103,_EVAL_496};
  assign _EVAL_109 = ~_EVAL_74;
  assign _EVAL_227 = _EVAL_229 & _EVAL_329;
  assign _EVAL_387 = _EVAL_18[0];
  assign _EVAL_420 = {_EVAL_478,_EVAL_263};
  assign _EVAL_248 = _EVAL_57[0];
  assign _EVAL_225 = _EVAL_69[0];
  assign _EVAL_423 = {_EVAL_344,_EVAL_56};
  assign _EVAL_216 = _EVAL_106 ? 4'he : 4'h8;
  assign _EVAL_84 = _EVAL_135 | _EVAL_87;
  assign _EVAL_241 = _EVAL_98[0];
  assign _EVAL_450 = _EVAL_424 & _EVAL_26;
  assign _EVAL_67 = _EVAL_281[2];
  assign _EVAL_235 = _EVAL_311[0];
  assign _EVAL_304 = ~_EVAL_364;
  assign _EVAL_471 = _EVAL_191[1];
  always @(posedge _EVAL_8) begin
    if (_EVAL_54) begin
      if (_EVAL_417) begin
        _EVAL_62 <= _EVAL_0;
      end
    end
    if (_EVAL_54) begin
      if (_EVAL_417) begin
        _EVAL_80 <= _EVAL_26;
      end
    end
    if (_EVAL_54) begin
      if (_EVAL_417) begin
        if (_EVAL_319) begin
          _EVAL_97 <= 4'hc;
        end else if (_EVAL_221) begin
          _EVAL_97 <= 4'h6;
        end else begin
          _EVAL_97 <= _EVAL_216;
        end
      end
    end
    if (_EVAL_54) begin
      if (_EVAL_417) begin
        _EVAL_112 <= _EVAL_46;
      end
    end
    if (_EVAL_54) begin
      if (_EVAL_417) begin
        _EVAL_133 <= _EVAL_16;
      end
    end
    if (_EVAL_54) begin
      if (_EVAL_417) begin
        _EVAL_141 <= _EVAL_2;
      end
    end
    if (_EVAL_352) begin
      if (_EVAL_255) begin
        _EVAL_143 <= _EVAL_11;
      end
    end
    if (_EVAL_54) begin
      if (_EVAL_417) begin
        _EVAL_152 <= _EVAL_48;
      end
    end
    if (_EVAL_44) begin
      _EVAL_161 <= 2'h0;
    end else if (_EVAL_352) begin
      if (_EVAL_467) begin
        if (_EVAL_449) begin
          _EVAL_161 <= 2'h2;
        end else begin
          _EVAL_161 <= 2'h0;
        end
      end else begin
        _EVAL_161 <= _EVAL_436;
      end
    end else begin
      _EVAL_161 <= _EVAL_436;
    end
    if (_EVAL_54) begin
      if (_EVAL_417) begin
        _EVAL_168 <= _EVAL_33;
      end
    end
    if (_EVAL_54) begin
      if (_EVAL_417) begin
        _EVAL_191 <= _EVAL_9;
      end
    end
    if (_EVAL_54) begin
      if (_EVAL_417) begin
        _EVAL_206 <= _EVAL_36;
      end
    end
    if (_EVAL_352) begin
      if (_EVAL_255) begin
        _EVAL_209 <= _EVAL_31;
      end
    end
    if (_EVAL_44) begin
      _EVAL_214 <= 6'h0;
    end else if (_EVAL_188) begin
      if (_EVAL_227) begin
        if (_EVAL_218) begin
          _EVAL_214 <= _EVAL_114;
        end else begin
          _EVAL_214 <= 6'h0;
        end
      end else begin
        _EVAL_214 <= 6'h0;
      end
    end else begin
      _EVAL_214 <= _EVAL_71;
    end
    if (_EVAL_44) begin
      _EVAL_238 <= 6'h0;
    end else if (_EVAL_212) begin
      if (_EVAL_193) begin
        if (_EVAL_387) begin
          _EVAL_238 <= _EVAL_290;
        end else begin
          _EVAL_238 <= 6'h0;
        end
      end else begin
        _EVAL_238 <= _EVAL_156;
      end
    end
    if (_EVAL_54) begin
      if (_EVAL_417) begin
        _EVAL_258 <= _EVAL_45;
      end
    end
    if (_EVAL_44) begin
      _EVAL_270 <= 1'h0;
    end else if (_EVAL_183) begin
      _EVAL_270 <= _EVAL_314;
    end
    if (_EVAL_54) begin
      if (_EVAL_417) begin
        _EVAL_416 <= _EVAL_27;
      end
    end
    if (_EVAL_54) begin
      if (_EVAL_417) begin
        _EVAL_441 <= _EVAL_12;
      end
    end
    if (_EVAL_352) begin
      if (_EVAL_255) begin
        _EVAL_462 <= _EVAL_25;
      end
    end
    if (_EVAL_44) begin
      _EVAL_483 <= 1'h0;
    end else if (_EVAL_183) begin
      _EVAL_483 <= _EVAL_227;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_62 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_80 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_97 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_112 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_133 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_141 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_143 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_152 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_161 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_168 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_191 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_206 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_209 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_214 = _RAND_13[5:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_238 = _RAND_14[5:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_258 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_270 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _EVAL_416 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _EVAL_441 = _RAND_18[2:0];
  _RAND_19 = {1{`RANDOM}};
  _EVAL_462 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  _EVAL_483 = _RAND_20[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
