//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_127_assert(
  input         _EVAL_83,
  input         _EVAL_85,
  input         _EVAL_102,
  input         _EVAL_121,
  input  [2:0]  _EVAL_134,
  input  [11:0] _EVAL_151,
  input         _EVAL_204,
  input         _EVAL_230,
  input         _EVAL_419,
  input         _EVAL_470,
  input         _EVAL_525,
  input  [31:0] _EVAL_531,
  input         _EVAL_663,
  input         _EVAL_687,
  input         _EVAL_701,
  input         _EVAL_802,
  input         _EVAL_881,
  input         _EVAL_882,
  input         _EVAL_909,
  input         _EVAL_913,
  input         _EVAL_954,
  input         _EVAL_973,
  input         _EVAL_999,
  input         _EVAL_1019,
  input         _EVAL_1031,
  input         _EVAL_1039,
  input         _EVAL_1041,
  input         _EVAL_1080,
  input         _EVAL_1084,
  input         _EVAL_1119,
  input         _EVAL_1136,
  input         _EVAL_1147,
  input         _EVAL_1172,
  input         _EVAL_1311,
  input         _EVAL_1323,
  input         _EVAL_1480,
  input         _EVAL_1485,
  input         _EVAL_1487,
  input         _EVAL_1526,
  input         _EVAL_1567,
  input         _EVAL_1586,
  input         _EVAL_1647,
  input         _EVAL_1702,
  input         _EVAL_1722,
  input         _EVAL_1731,
  input         _EVAL_1839,
  input         _EVAL_1912,
  input         _EVAL_1930,
  input         _EVAL_1962,
  input         _EVAL_2041,
  input         _EVAL_2063,
  input         _EVAL_2064,
  input         _EVAL_2067,
  input         _EVAL_2069,
  input         _EVAL_2087,
  input         _EVAL_2192,
  input         _EVAL_2246,
  input         _EVAL_2279,
  input         _EVAL_2291,
  input         _EVAL_2306,
  input         _EVAL_2338,
  input         _EVAL_2343,
  input         _EVAL_2359,
  input         _EVAL_2371,
  input         _EVAL_2393,
  input         _EVAL_2398,
  input         _EVAL_2447,
  input         _EVAL_2466,
  input         _EVAL_2505,
  input         _EVAL_2530
);
  wire  _EVAL_193;
  wire  _EVAL_198;
  wire  _EVAL_203;
  wire  _EVAL_206;
  wire  _EVAL_211;
  wire  _EVAL_219;
  wire  _EVAL_224;
  wire  _EVAL_226;
  wire  _EVAL_229;
  wire  _EVAL_247;
  wire  _EVAL_252;
  wire  _EVAL_255;
  wire  _EVAL_259;
  wire  _EVAL_261;
  wire  _EVAL_264;
  wire  _EVAL_266;
  wire  _EVAL_269;
  wire  _EVAL_272;
  wire  _EVAL_276;
  wire  _EVAL_285;
  wire  _EVAL_290;
  wire  _EVAL_292;
  wire  _EVAL_294;
  wire  _EVAL_296;
  wire  _EVAL_301;
  wire  _EVAL_309;
  wire  _EVAL_328;
  wire  _EVAL_331;
  wire  _EVAL_335;
  wire  _EVAL_339;
  wire  _EVAL_340;
  wire  _EVAL_341;
  wire  _EVAL_344;
  wire  _EVAL_347;
  wire  _EVAL_352;
  wire  _EVAL_371;
  wire  _EVAL_374;
  wire  _EVAL_376;
  wire  _EVAL_399;
  wire  _EVAL_406;
  wire  _EVAL_411;
  wire  _EVAL_415;
  wire  _EVAL_425;
  wire  _EVAL_433;
  wire  _EVAL_435;
  wire  _EVAL_453;
  wire  _EVAL_458;
  wire  _EVAL_464;
  wire  _EVAL_467;
  wire  _EVAL_475;
  wire  _EVAL_478;
  wire  _EVAL_479;
  wire  _EVAL_489;
  wire  _EVAL_496;
  wire  _EVAL_510;
  wire  _EVAL_518;
  wire  _EVAL_520;
  wire  _EVAL_522;
  wire  _EVAL_526;
  wire  _EVAL_538;
  wire  _EVAL_544;
  wire  _EVAL_557;
  wire  _EVAL_574;
  wire  _EVAL_578;
  wire  _EVAL_583;
  wire  _EVAL_586;
  wire  _EVAL_588;
  wire  _EVAL_603;
  wire  _EVAL_605;
  wire  _EVAL_609;
  wire  _EVAL_613;
  wire  _EVAL_633;
  wire  _EVAL_636;
  wire  _EVAL_643;
  wire  _EVAL_644;
  wire  _EVAL_645;
  wire  _EVAL_648;
  wire  _EVAL_656;
  wire  _EVAL_664;
  wire  _EVAL_669;
  wire  _EVAL_677;
  wire  _EVAL_678;
  wire  _EVAL_680;
  wire  _EVAL_693;
  wire  _EVAL_698;
  wire  _EVAL_716;
  wire  _EVAL_719;
  wire  _EVAL_738;
  wire  _EVAL_742;
  wire  _EVAL_746;
  wire  _EVAL_749;
  wire  _EVAL_750;
  wire  _EVAL_751;
  wire  _EVAL_752;
  wire  _EVAL_758;
  wire  _EVAL_761;
  wire  _EVAL_762;
  wire  _EVAL_764;
  wire  _EVAL_766;
  wire  _EVAL_774;
  wire  _EVAL_777;
  wire  _EVAL_785;
  wire  _EVAL_786;
  wire  _EVAL_789;
  wire  _EVAL_794;
  wire  _EVAL_806;
  wire  _EVAL_808;
  wire  _EVAL_812;
  wire  _EVAL_813;
  wire  _EVAL_814;
  wire  _EVAL_822;
  wire  _EVAL_826;
  wire  _EVAL_827;
  wire  _EVAL_829;
  wire  _EVAL_838;
  wire  _EVAL_839;
  wire  _EVAL_841;
  wire  _EVAL_864;
  wire  _EVAL_868;
  wire  _EVAL_884;
  wire  _EVAL_886;
  wire  _EVAL_887;
  wire  _EVAL_900;
  wire  _EVAL_908;
  wire  _EVAL_923;
  wire  _EVAL_940;
  wire  _EVAL_944;
  wire  _EVAL_946;
  wire  _EVAL_948;
  wire  _EVAL_950;
  wire  _EVAL_953;
  wire  _EVAL_961;
  wire  _EVAL_976;
  wire  _EVAL_977;
  wire  _EVAL_978;
  wire  _EVAL_979;
  wire  _EVAL_982;
  wire  _EVAL_984;
  wire  _EVAL_987;
  wire  _EVAL_988;
  wire  _EVAL_992;
  wire  _EVAL_994;
  wire  _EVAL_998;
  wire  _EVAL_1004;
  wire  _EVAL_1008;
  wire  _EVAL_1011;
  wire  _EVAL_1020;
  wire  _EVAL_1021;
  wire  _EVAL_1026;
  wire  _EVAL_1044;
  wire  _EVAL_1054;
  wire  _EVAL_1055;
  wire  _EVAL_1061;
  wire  _EVAL_1071;
  wire  _EVAL_1078;
  wire  _EVAL_1087;
  wire  _EVAL_1089;
  wire  _EVAL_1093;
  wire  _EVAL_1098;
  wire  _EVAL_1101;
  wire  _EVAL_1104;
  wire  _EVAL_1106;
  wire  _EVAL_1108;
  wire  _EVAL_1115;
  wire  _EVAL_1127;
  wire  _EVAL_1134;
  wire  _EVAL_1138;
  wire  _EVAL_1148;
  wire  _EVAL_1152;
  wire  _EVAL_1154;
  wire  _EVAL_1156;
  wire  _EVAL_1158;
  wire  _EVAL_1162;
  wire  _EVAL_1165;
  wire  _EVAL_1166;
  wire  _EVAL_1173;
  wire  _EVAL_1176;
  wire  _EVAL_1184;
  wire  _EVAL_1185;
  wire  _EVAL_1188;
  wire  _EVAL_1197;
  wire  _EVAL_1199;
  wire  _EVAL_1205;
  wire  _EVAL_1207;
  wire  _EVAL_1224;
  wire  _EVAL_1225;
  wire  _EVAL_1226;
  wire  _EVAL_1232;
  wire  _EVAL_1234;
  wire  _EVAL_1236;
  wire  _EVAL_1237;
  wire  _EVAL_1241;
  wire  _EVAL_1242;
  wire  _EVAL_1243;
  wire  _EVAL_1247;
  wire  _EVAL_1253;
  wire  _EVAL_1257;
  wire  _EVAL_1258;
  wire  _EVAL_1263;
  wire  _EVAL_1267;
  wire  _EVAL_1268;
  wire  _EVAL_1269;
  wire  _EVAL_1272;
  wire  _EVAL_1277;
  wire  _EVAL_1278;
  wire  _EVAL_1281;
  wire  _EVAL_1292;
  wire  _EVAL_1295;
  wire  _EVAL_1296;
  wire  _EVAL_1299;
  wire  _EVAL_1307;
  wire  _EVAL_1317;
  wire  _EVAL_1325;
  wire  _EVAL_1338;
  wire  _EVAL_1343;
  wire  _EVAL_1352;
  wire  _EVAL_1353;
  wire  _EVAL_1356;
  wire  _EVAL_1361;
  wire  _EVAL_1365;
  wire  _EVAL_1368;
  wire  _EVAL_1370;
  wire  _EVAL_1375;
  wire  _EVAL_1382;
  wire  _EVAL_1387;
  wire  _EVAL_1390;
  wire  _EVAL_1397;
  wire  _EVAL_1400;
  wire  _EVAL_1403;
  wire  _EVAL_1408;
  wire  _EVAL_1409;
  wire  _EVAL_1412;
  wire  _EVAL_1419;
  wire  _EVAL_1426;
  wire  _EVAL_1433;
  wire  _EVAL_1434;
  wire  _EVAL_1435;
  wire  _EVAL_1443;
  wire  _EVAL_1453;
  wire  _EVAL_1462;
  wire  _EVAL_1464;
  wire  _EVAL_1466;
  wire  _EVAL_1469;
  wire  _EVAL_1473;
  wire  _EVAL_1475;
  wire [2:0] _EVAL_1477;
  wire  _EVAL_1488;
  wire  _EVAL_1491;
  wire  _EVAL_1506;
  wire  _EVAL_1507;
  wire  _EVAL_1508;
  wire  _EVAL_1513;
  wire  _EVAL_1523;
  wire  _EVAL_1530;
  wire  _EVAL_1538;
  wire  _EVAL_1542;
  wire  _EVAL_1548;
  wire  _EVAL_1552;
  wire  _EVAL_1555;
  wire  _EVAL_1559;
  wire  _EVAL_1570;
  wire  _EVAL_1572;
  wire  _EVAL_1577;
  wire  _EVAL_1578;
  wire  _EVAL_1585;
  wire  _EVAL_1591;
  wire  _EVAL_1596;
  wire  _EVAL_1603;
  wire  _EVAL_1605;
  wire  _EVAL_1611;
  wire  _EVAL_1617;
  wire  _EVAL_1624;
  wire  _EVAL_1626;
  wire  _EVAL_1632;
  wire  _EVAL_1638;
  wire  _EVAL_1649;
  wire  _EVAL_1650;
  wire  _EVAL_1653;
  wire  _EVAL_1655;
  wire  _EVAL_1656;
  wire  _EVAL_1666;
  wire  _EVAL_1671;
  wire  _EVAL_1673;
  wire  _EVAL_1674;
  wire  _EVAL_1676;
  wire  _EVAL_1680;
  wire  _EVAL_1685;
  wire  _EVAL_1703;
  wire  _EVAL_1704;
  wire  _EVAL_1711;
  wire  _EVAL_1713;
  wire  _EVAL_1726;
  wire  _EVAL_1743;
  wire  _EVAL_1746;
  wire  _EVAL_1747;
  wire  _EVAL_1763;
  wire  _EVAL_1769;
  wire  _EVAL_1774;
  wire  _EVAL_1781;
  wire  _EVAL_1784;
  wire  _EVAL_1811;
  wire  _EVAL_1814;
  wire  _EVAL_1815;
  wire  _EVAL_1831;
  wire  _EVAL_1837;
  wire  _EVAL_1840;
  wire  _EVAL_1842;
  wire  _EVAL_1846;
  wire  _EVAL_1853;
  wire  _EVAL_1864;
  wire  _EVAL_1868;
  wire  _EVAL_1871;
  wire  _EVAL_1875;
  wire  _EVAL_1895;
  wire  _EVAL_1900;
  wire  _EVAL_1902;
  wire  _EVAL_1908;
  wire  _EVAL_1917;
  wire  _EVAL_1932;
  wire  _EVAL_1960;
  wire  _EVAL_1965;
  wire  _EVAL_1972;
  wire  _EVAL_1973;
  wire  _EVAL_1975;
  wire  _EVAL_1979;
  wire  _EVAL_1982;
  wire  _EVAL_1986;
  wire  _EVAL_2002;
  wire  _EVAL_2008;
  wire  _EVAL_2019;
  wire [1:0] _EVAL_2023;
  wire  _EVAL_2040;
  wire  _EVAL_2050;
  wire  _EVAL_2068;
  wire  _EVAL_2070;
  wire  _EVAL_2076;
  wire  _EVAL_2081;
  wire  _EVAL_2083;
  wire  _EVAL_2094;
  wire  _EVAL_2097;
  wire  _EVAL_2100;
  wire  _EVAL_2101;
  wire  _EVAL_2106;
  wire  _EVAL_2111;
  wire [1:0] _EVAL_2116;
  wire  _EVAL_2118;
  wire  _EVAL_2136;
  wire  _EVAL_2139;
  wire  _EVAL_2152;
  wire  _EVAL_2156;
  wire  _EVAL_2161;
  wire  _EVAL_2167;
  wire  _EVAL_2194;
  wire  _EVAL_2203;
  wire  _EVAL_2204;
  wire  _EVAL_2205;
  wire  _EVAL_2207;
  wire  _EVAL_2213;
  wire  _EVAL_2216;
  wire  _EVAL_2220;
  wire  _EVAL_2224;
  wire  _EVAL_2227;
  wire  _EVAL_2228;
  wire  _EVAL_2230;
  wire  _EVAL_2231;
  wire  _EVAL_2233;
  wire  _EVAL_2235;
  wire  _EVAL_2236;
  wire  _EVAL_2237;
  wire  _EVAL_2240;
  wire  _EVAL_2252;
  wire  _EVAL_2254;
  wire  _EVAL_2259;
  wire  _EVAL_2261;
  wire  _EVAL_2264;
  wire  _EVAL_2273;
  wire  _EVAL_2281;
  wire  _EVAL_2286;
  wire  _EVAL_2288;
  wire  _EVAL_2289;
  wire  _EVAL_2290;
  wire  _EVAL_2293;
  wire  _EVAL_2299;
  wire  _EVAL_2300;
  wire  _EVAL_2302;
  wire  _EVAL_2311;
  wire  _EVAL_2312;
  wire  _EVAL_2317;
  wire  _EVAL_2324;
  wire  _EVAL_2341;
  wire  _EVAL_2348;
  wire  _EVAL_2351;
  wire  _EVAL_2353;
  wire  _EVAL_2356;
  wire  _EVAL_2360;
  wire  _EVAL_2364;
  wire  _EVAL_2370;
  wire  _EVAL_2373;
  wire  _EVAL_2375;
  wire  _EVAL_2380;
  wire  _EVAL_2383;
  wire  _EVAL_2395;
  wire  _EVAL_2406;
  wire  _EVAL_2407;
  wire  _EVAL_2408;
  wire  _EVAL_2419;
  wire  _EVAL_2424;
  wire  _EVAL_2438;
  wire  _EVAL_2443;
  wire  _EVAL_2450;
  wire  _EVAL_2453;
  wire  _EVAL_2459;
  wire  _EVAL_2464;
  wire  _EVAL_2499;
  wire  _EVAL_2509;
  wire  _EVAL_2515;
  wire  _EVAL_2523;
  wire  _EVAL_2531;
  wire  _EVAL_2533;
  wire  _EVAL_2545;
  assign _EVAL_1267 = _EVAL_2371 & _EVAL_1061;
  assign _EVAL_1412 = _EVAL_531 == 32'h8000001b;
  assign _EVAL_2299 = _EVAL_2167 & _EVAL_1172;
  assign _EVAL_680 = _EVAL_1224 & _EVAL_2139;
  assign _EVAL_603 = _EVAL_1224 & _EVAL_2259;
  assign _EVAL_1241 = _EVAL_1224 & _EVAL_999;
  assign _EVAL_2002 = _EVAL_151 == 12'h327;
  assign _EVAL_987 = _EVAL_1224 & _EVAL_1299;
  assign _EVAL_510 = _EVAL_2167 & _EVAL_2094;
  assign _EVAL_1237 = _EVAL_2371 & _EVAL_518;
  assign _EVAL_1268 = _EVAL_1224 & _EVAL_1655;
  assign _EVAL_2300 = _EVAL_151 == 12'hc85;
  assign _EVAL_435 = _EVAL_531 == 32'h3;
  assign _EVAL_1671 = _EVAL_1224 & _EVAL_1148;
  assign _EVAL_643 = _EVAL_151 == 12'h333;
  assign _EVAL_982 = _EVAL_1224 & _EVAL_1526;
  assign _EVAL_1982 = _EVAL_1224 & _EVAL_886;
  assign _EVAL_211 = _EVAL_1224 & _EVAL_1119;
  assign _EVAL_785 = _EVAL_151 == 12'hb0d;
  assign _EVAL_2459 = _EVAL_151 == 12'hb8e;
  assign _EVAL_526 = _EVAL_151 == 12'hb96;
  assign _EVAL_2395 = _EVAL_151 == 12'hc07;
  assign _EVAL_1257 = _EVAL_1224 & _EVAL_1567;
  assign _EVAL_868 = _EVAL_1224 & _EVAL_1972;
  assign _EVAL_900 = _EVAL_151 == 12'h33b;
  assign _EVAL_2261 = _EVAL_531 == 32'h6;
  assign _EVAL_2293 = _EVAL_1224 & _EVAL_1676;
  assign _EVAL_1176 = _EVAL_151 == 12'hc8e;
  assign _EVAL_789 = _EVAL_151 == 12'hb07;
  assign _EVAL_1769 = _EVAL_151 == 12'h33e;
  assign _EVAL_698 = _EVAL_1224 & _EVAL_2220;
  assign _EVAL_669 = _EVAL_1224 & _EVAL_479;
  assign _EVAL_1338 = _EVAL_841 | _EVAL_1711;
  assign _EVAL_946 = _EVAL_1224 & _EVAL_1031;
  assign _EVAL_2351 = _EVAL_2371 & _EVAL_1412;
  assign _EVAL_2167 = _EVAL_134 == 3'h2;
  assign _EVAL_1831 = _EVAL_2167 & _EVAL_1871;
  assign _EVAL_1559 = _EVAL_151 == 12'hc9d;
  assign _EVAL_1530 = _EVAL_1224 & _EVAL_701;
  assign _EVAL_1258 = _EVAL_151 == 12'hc06;
  assign _EVAL_813 = _EVAL_2167 & _EVAL_1071;
  assign _EVAL_1837 = _EVAL_1224 & _EVAL_1409;
  assign _EVAL_2240 = _EVAL_151 == 12'hb10;
  assign _EVAL_1277 = _EVAL_151 == 12'h328;
  assign _EVAL_475 = _EVAL_2167 & _EVAL_2252;
  assign _EVAL_1973 = _EVAL_1224 & _EVAL_913;
  assign _EVAL_1409 = _EVAL_151 == 12'h7a3;
  assign _EVAL_2348 = _EVAL_2167 & _EVAL_1488;
  assign _EVAL_1148 = _EVAL_151 == 12'hb0f;
  assign _EVAL_613 = _EVAL_2371 & _EVAL_1596;
  assign _EVAL_224 = _EVAL_531 == 32'h4;
  assign _EVAL_1224 = _EVAL_1680 | _EVAL_1722;
  assign _EVAL_1908 = _EVAL_2167 & _EVAL_1443;
  assign _EVAL_2364 = _EVAL_151 == 12'hb91;
  assign _EVAL_774 = ~_EVAL_83;
  assign _EVAL_1763 = _EVAL_1224 & _EVAL_1624;
  assign _EVAL_247 = _EVAL_151 == 12'hc92;
  assign _EVAL_538 = _EVAL_1224 & _EVAL_411;
  assign _EVAL_1676 = _EVAL_151 == 12'hb0b;
  assign _EVAL_2360 = _EVAL_151 == 12'hc1c;
  assign _EVAL_1071 = _EVAL_151 == 12'hc96;
  assign _EVAL_636 = _EVAL_2167 & _EVAL_687;
  assign _EVAL_1840 = _EVAL_1224 & _EVAL_909;
  assign _EVAL_2116 = _EVAL_204 + _EVAL_102;
  assign _EVAL_2230 = _EVAL_2167 & _EVAL_247;
  assign _EVAL_376 = _EVAL_151 == 12'hb1a;
  assign _EVAL_2288 = _EVAL_1224 & _EVAL_2306;
  assign _EVAL_1026 = _EVAL_151 == 12'hb0e;
  assign _EVAL_269 = _EVAL_2167 & _EVAL_2380;
  assign _EVAL_884 = _EVAL_1224 & _EVAL_2424;
  assign _EVAL_1199 = _EVAL_1224 & _EVAL_1080;
  assign _EVAL_1466 = _EVAL_2167 & _EVAL_1453;
  assign _EVAL_1343 = _EVAL_531 == 32'h80000003;
  assign _EVAL_352 = _EVAL_2371 & _EVAL_1292;
  assign _EVAL_578 = _EVAL_1224 & _EVAL_643;
  assign _EVAL_1020 = _EVAL_1224 & _EVAL_2235;
  assign _EVAL_266 = _EVAL_2167 & _EVAL_276;
  assign _EVAL_294 = _EVAL_1603 | _EVAL_83;
  assign _EVAL_1004 = _EVAL_1224 & _EVAL_2515;
  assign _EVAL_746 = _EVAL_1224 & _EVAL_749;
  assign _EVAL_976 = _EVAL_531 == 32'h80000007;
  assign _EVAL_2281 = _EVAL_151 == 12'hb18;
  assign _EVAL_1781 = _EVAL_151 == 12'hc19;
  assign _EVAL_1008 = _EVAL_2167 & _EVAL_2136;
  assign _EVAL_742 = _EVAL_1224 & _EVAL_1626;
  assign _EVAL_758 = _EVAL_1224 & _EVAL_1473;
  assign _EVAL_2273 = ~_EVAL_294;
  assign _EVAL_1370 = _EVAL_151 == 12'hc0c;
  assign _EVAL_583 = _EVAL_151 == 12'hb87;
  assign _EVAL_908 = _EVAL_1224 & _EVAL_2530;
  assign _EVAL_2076 = _EVAL_151 == 12'hb8a;
  assign _EVAL_339 = _EVAL_1224 & _EVAL_2531;
  assign _EVAL_586 = _EVAL_2167 & _EVAL_1962;
  assign _EVAL_633 = _EVAL_2167 & _EVAL_1586;
  assign _EVAL_340 = _EVAL_151 == 12'hb08;
  assign _EVAL_1475 = _EVAL_151 == 12'h326;
  assign _EVAL_1387 = _EVAL_1224 & _EVAL_1673;
  assign _EVAL_292 = _EVAL_2167 & _EVAL_1577;
  assign _EVAL_2533 = _EVAL_1224 & _EVAL_2207;
  assign _EVAL_979 = _EVAL_531 == 32'h80000015;
  assign _EVAL_1236 = _EVAL_2167 & _EVAL_2118;
  assign _EVAL_678 = _EVAL_2167 & _EVAL_2216;
  assign _EVAL_749 = _EVAL_151 == 12'hb1d;
  assign _EVAL_764 = _EVAL_1224 & _EVAL_839;
  assign _EVAL_2083 = _EVAL_1224 & _EVAL_341;
  assign _EVAL_301 = _EVAL_1224 & _EVAL_1136;
  assign _EVAL_2353 = _EVAL_151 == 12'hc97;
  assign _EVAL_1784 = _EVAL_2371 & _EVAL_224;
  assign _EVAL_1811 = _EVAL_1224 & _EVAL_371;
  assign _EVAL_1650 = _EVAL_1224 & _EVAL_1647;
  assign _EVAL_1596 = _EVAL_531 == 32'h80000011;
  assign _EVAL_1247 = _EVAL_2371 & _EVAL_2356;
  assign _EVAL_1655 = _EVAL_151 == 12'h3b9;
  assign _EVAL_1242 = _EVAL_151 == 12'hb15;
  assign _EVAL_520 = _EVAL_1224 & _EVAL_1277;
  assign _EVAL_766 = _EVAL_151 == 12'hb8c;
  assign _EVAL_609 = _EVAL_2167 & _EVAL_1370;
  assign _EVAL_252 = _EVAL_2167 & _EVAL_1930;
  assign _EVAL_467 = _EVAL_1224 & _EVAL_1703;
  assign _EVAL_193 = _EVAL_1224 & _EVAL_1408;
  assign _EVAL_814 = _EVAL_2371 & _EVAL_1868;
  assign _EVAL_1138 = _EVAL_2167 & _EVAL_331;
  assign _EVAL_827 = _EVAL_2371 & _EVAL_2523;
  assign _EVAL_1281 = _EVAL_1338 | _EVAL_83;
  assign _EVAL_1746 = _EVAL_1224 & _EVAL_2227;
  assign _EVAL_2406 = _EVAL_151 == 12'h3ba;
  assign _EVAL_1253 = _EVAL_1224 & _EVAL_376;
  assign _EVAL_1673 = _EVAL_151 == 12'h334;
  assign _EVAL_2097 = _EVAL_1224 & _EVAL_1352;
  assign _EVAL_1435 = _EVAL_151 == 12'hb86;
  assign _EVAL_794 = _EVAL_1224 & _EVAL_406;
  assign _EVAL_2289 = _EVAL_531 == 32'h8000001e;
  assign _EVAL_2008 = _EVAL_1224 & _EVAL_1101;
  assign _EVAL_2070 = _EVAL_531 == 32'h80000013;
  assign _EVAL_887 = _EVAL_2371 & _EVAL_1513;
  assign _EVAL_2216 = _EVAL_151 == 12'hc86;
  assign _EVAL_1842 = _EVAL_151 == 12'hb88;
  assign _EVAL_479 = _EVAL_151 == 12'h332;
  assign _EVAL_1361 = _EVAL_2167 & _EVAL_645;
  assign _EVAL_1433 = _EVAL_1224 & _EVAL_1021;
  assign _EVAL_829 = _EVAL_531 == 32'h80000017;
  assign _EVAL_1234 = _EVAL_1224 & _EVAL_1726;
  assign _EVAL_826 = _EVAL_1224 & _EVAL_2291;
  assign _EVAL_838 = _EVAL_531 == 32'h2;
  assign _EVAL_1960 = _EVAL_2167 & _EVAL_1185;
  assign _EVAL_994 = _EVAL_151 == 12'hc1d;
  assign _EVAL_2373 = _EVAL_1224 & _EVAL_2064;
  assign _EVAL_1011 = _EVAL_2167 & _EVAL_2311;
  assign _EVAL_1864 = _EVAL_151 == 12'hb90;
  assign _EVAL_656 = _EVAL_1224 & _EVAL_648;
  assign _EVAL_645 = _EVAL_151 == 12'hc9f;
  assign _EVAL_864 = _EVAL_2167 & _EVAL_1419;
  assign _EVAL_544 = _EVAL_2167 & _EVAL_1098;
  assign _EVAL_2068 = _EVAL_2167 & _EVAL_470;
  assign _EVAL_1979 = _EVAL_1224 & _EVAL_992;
  assign _EVAL_953 = _EVAL_1224 & _EVAL_644;
  assign _EVAL_2213 = _EVAL_151 == 12'hb89;
  assign _EVAL_1154 = _EVAL_151 == 12'h32b;
  assign _EVAL_1713 = _EVAL_1224 & _EVAL_2393;
  assign _EVAL_1269 = _EVAL_151 == 12'hc8a;
  assign _EVAL_1207 = _EVAL_2167 & _EVAL_347;
  assign _EVAL_2203 = _EVAL_1224 & _EVAL_526;
  assign _EVAL_433 = _EVAL_1224 & _EVAL_583;
  assign _EVAL_2023 = _EVAL_2279 + _EVAL_525;
  assign _EVAL_1508 = _EVAL_2167 & _EVAL_2228;
  assign _EVAL_1473 = _EVAL_151 == 12'h337;
  assign _EVAL_2259 = _EVAL_151 == 12'h325;
  assign _EVAL_453 = _EVAL_151 == 12'hc98;
  assign _EVAL_1115 = _EVAL_1224 & _EVAL_1704;
  assign _EVAL_1307 = _EVAL_151 == 12'hb9d;
  assign _EVAL_2312 = _EVAL_151 == 12'hc16;
  assign _EVAL_347 = _EVAL_151 == 12'hc12;
  assign _EVAL_2290 = _EVAL_151 == 12'h32a;
  assign _EVAL_2419 = _EVAL_531 == 32'h5;
  assign _EVAL_2407 = _EVAL_151 == 12'hc89;
  assign _EVAL_285 = _EVAL_1224 & _EVAL_1243;
  assign _EVAL_2237 = _EVAL_151 == 12'h339;
  assign _EVAL_2081 = _EVAL_2167 & _EVAL_1731;
  assign _EVAL_1548 = _EVAL_2371 & _EVAL_1087;
  assign _EVAL_522 = _EVAL_151 == 12'hb9b;
  assign _EVAL_1375 = _EVAL_1224 & _EVAL_961;
  assign _EVAL_1685 = _EVAL_151 == 12'hc1a;
  assign _EVAL_841 = ~_EVAL_2069;
  assign _EVAL_648 = _EVAL_151 == 12'h329;
  assign _EVAL_1632 = _EVAL_2167 & _EVAL_1685;
  assign _EVAL_886 = _EVAL_151 == 12'hb12;
  assign _EVAL_2464 = _EVAL_2371 & _EVAL_435;
  assign _EVAL_259 = _EVAL_1224 & _EVAL_2505;
  assign _EVAL_2509 = _EVAL_2167 & _EVAL_1469;
  assign _EVAL_2443 = _EVAL_1224 & _EVAL_1487;
  assign _EVAL_1666 = _EVAL_2167 & _EVAL_719;
  assign _EVAL_478 = _EVAL_151 == 12'hc8f;
  assign _EVAL_2228 = _EVAL_151 == 12'hc95;
  assign _EVAL_2252 = _EVAL_151 == 12'hc11;
  assign _EVAL_1462 = _EVAL_2167 & _EVAL_1781;
  assign _EVAL_1044 = _EVAL_1224 & _EVAL_2281;
  assign _EVAL_2370 = _EVAL_2167 & _EVAL_1269;
  assign _EVAL_1488 = _EVAL_151 == 12'hc9c;
  assign _EVAL_1243 = _EVAL_151 == 12'hb14;
  assign _EVAL_1108 = _EVAL_2371 & _EVAL_1434;
  assign _EVAL_1704 = _EVAL_151 == 12'hb16;
  assign _EVAL_2111 = _EVAL_1224 & _EVAL_1435;
  assign _EVAL_2341 = _EVAL_151 == 12'hc10;
  assign _EVAL_1653 = _EVAL_1224 & _EVAL_340;
  assign _EVAL_1104 = _EVAL_151 == 12'hc90;
  assign _EVAL_406 = _EVAL_151 == 12'h330;
  assign _EVAL_961 = _EVAL_151 == 12'h33f;
  assign _EVAL_1975 = _EVAL_151 == 12'hc18;
  assign _EVAL_2264 = _EVAL_151 == 12'hc8c;
  assign _EVAL_1591 = _EVAL_151 == 12'hb13;
  assign _EVAL_1365 = _EVAL_1224 & _EVAL_2359;
  assign _EVAL_574 = _EVAL_2371 & _EVAL_1382;
  assign _EVAL_1158 = _EVAL_2167 & _EVAL_1875;
  assign _EVAL_1397 = _EVAL_1224 & _EVAL_2205;
  assign _EVAL_2311 = _EVAL_151 == 12'hc08;
  assign _EVAL_2236 = _EVAL_1224 & _EVAL_2290;
  assign _EVAL_1603 = _EVAL_1477 <= 3'h1;
  assign _EVAL_1382 = _EVAL_531 == 32'h80000019;
  assign _EVAL_588 = _EVAL_2167 & _EVAL_2019;
  assign _EVAL_808 = _EVAL_1224 & _EVAL_2076;
  assign _EVAL_1513 = _EVAL_531 == 32'h80000018;
  assign _EVAL_1871 = _EVAL_151 == 12'hc99;
  assign _EVAL_219 = _EVAL_1224 & _EVAL_496;
  assign _EVAL_2231 = _EVAL_2167 & _EVAL_2312;
  assign _EVAL_944 = ~_EVAL_1281;
  assign _EVAL_2286 = _EVAL_2371 & _EVAL_464;
  assign _EVAL_1184 = _EVAL_2371 & _EVAL_1343;
  assign _EVAL_1815 = _EVAL_1224 & _EVAL_2192;
  assign _EVAL_1656 = _EVAL_151 == 12'hb85;
  assign _EVAL_2356 = _EVAL_531 == 32'h8000000b;
  assign _EVAL_198 = _EVAL_151 == 12'hb11;
  assign _EVAL_335 = _EVAL_2167 & _EVAL_226;
  assign _EVAL_1299 = _EVAL_151 == 12'h33c;
  assign _EVAL_978 = _EVAL_1224 & _EVAL_2338;
  assign _EVAL_290 = _EVAL_1224 & _EVAL_2213;
  assign _EVAL_1638 = _EVAL_2371 & _EVAL_829;
  assign _EVAL_557 = _EVAL_1224 & _EVAL_663;
  assign _EVAL_777 = _EVAL_1224 & _EVAL_415;
  assign _EVAL_1166 = _EVAL_2167 & _EVAL_881;
  assign _EVAL_2139 = _EVAL_151 == 12'hb97;
  assign _EVAL_2302 = _EVAL_1224 & _EVAL_789;
  assign _EVAL_750 = _EVAL_2167 & _EVAL_2466;
  assign _EVAL_2324 = _EVAL_2167 & _EVAL_1747;
  assign _EVAL_1426 = _EVAL_2167 & _EVAL_2341;
  assign _EVAL_1507 = _EVAL_2167 & _EVAL_693;
  assign _EVAL_1356 = _EVAL_1224 & _EVAL_1041;
  assign _EVAL_1205 = _EVAL_151 == 12'h32d;
  assign _EVAL_644 = _EVAL_151 == 12'h3a3;
  assign _EVAL_1542 = _EVAL_1224 & _EVAL_2101;
  assign _EVAL_2254 = _EVAL_2167 & _EVAL_1555;
  assign _EVAL_1443 = _EVAL_151 == 12'hc0d;
  assign _EVAL_458 = _EVAL_2167 & _EVAL_1104;
  assign _EVAL_2453 = _EVAL_1224 & _EVAL_1902;
  assign _EVAL_2207 = _EVAL_151 == 12'hb0c;
  assign _EVAL_206 = _EVAL_151 == 12'h3bd;
  assign _EVAL_1585 = _EVAL_1224 & _EVAL_1475;
  assign _EVAL_2515 = _EVAL_151 == 12'hb8f;
  assign _EVAL_2101 = _EVAL_151 == 12'h338;
  assign _EVAL_1617 = _EVAL_531 == 32'h8000001f;
  assign _EVAL_2499 = _EVAL_1224 & _EVAL_2002;
  assign _EVAL_1101 = _EVAL_151 == 12'hb98;
  assign _EVAL_272 = _EVAL_151 == 12'hc91;
  assign _EVAL_1572 = _EVAL_2371 & _EVAL_2289;
  assign _EVAL_1453 = _EVAL_151 == 12'hc9a;
  assign _EVAL_1061 = _EVAL_531 == 32'hb;
  assign _EVAL_1649 = _EVAL_1224 & _EVAL_2041;
  assign _EVAL_1972 = _EVAL_151 == 12'hb92;
  assign _EVAL_1054 = _EVAL_1224 & _EVAL_1205;
  assign _EVAL_2317 = _EVAL_151 == 12'h3bc;
  assign _EVAL_1680 = _EVAL_2087 | _EVAL_2067;
  assign _EVAL_425 = _EVAL_2167 & _EVAL_1258;
  assign _EVAL_2531 = _EVAL_151 == 12'hb1c;
  assign _EVAL_1477 = _EVAL_2023 + _EVAL_2116;
  assign _EVAL_2118 = _EVAL_151 == 12'hc8d;
  assign _EVAL_1325 = _EVAL_151 == 12'hc1f;
  assign _EVAL_1577 = _EVAL_151 == 12'hc9b;
  assign _EVAL_1846 = _EVAL_2167 & _EVAL_2040;
  assign _EVAL_1127 = _EVAL_2371 & _EVAL_979;
  assign _EVAL_2227 = _EVAL_151 == 12'hb9c;
  assign _EVAL_2220 = _EVAL_151 == 12'hb9f;
  assign _EVAL_1419 = _EVAL_151 == 12'hc0f;
  assign _EVAL_1272 = _EVAL_1224 & _EVAL_900;
  assign _EVAL_2383 = _EVAL_1224 & _EVAL_1485;
  assign _EVAL_762 = _EVAL_2167 & _EVAL_230;
  assign _EVAL_374 = _EVAL_151 == 12'hb9a;
  assign _EVAL_1098 = _EVAL_151 == 12'hc13;
  assign _EVAL_1087 = _EVAL_531 == 32'h8000001d;
  assign _EVAL_605 = _EVAL_1224 & _EVAL_785;
  assign _EVAL_1875 = _EVAL_151 == 12'hc17;
  assign _EVAL_664 = _EVAL_2371 & _EVAL_2419;
  assign _EVAL_464 = _EVAL_531 == 32'h7;
  assign _EVAL_1506 = _EVAL_151 == 12'h32e;
  assign _EVAL_2450 = _EVAL_1224 & _EVAL_198;
  assign _EVAL_806 = _EVAL_2167 & _EVAL_478;
  assign _EVAL_1134 = _EVAL_2167 & _EVAL_2398;
  assign _EVAL_399 = _EVAL_1224 & _EVAL_2343;
  assign _EVAL_296 = _EVAL_1224 & _EVAL_1605;
  assign _EVAL_1165 = _EVAL_2371 & _EVAL_2070;
  assign _EVAL_341 = _EVAL_151 == 12'h335;
  assign _EVAL_415 = _EVAL_151 == 12'h3be;
  assign _EVAL_1932 = _EVAL_1224 & _EVAL_882;
  assign _EVAL_1317 = _EVAL_151 == 12'hb93;
  assign _EVAL_1278 = _EVAL_2167 & _EVAL_272;
  assign _EVAL_264 = _EVAL_1224 & _EVAL_1506;
  assign _EVAL_1156 = _EVAL_2371 & _EVAL_838;
  assign _EVAL_1895 = _EVAL_531 == 32'h80000012;
  assign _EVAL_998 = _EVAL_2167 & _EVAL_994;
  assign _EVAL_1296 = _EVAL_1224 & _EVAL_2063;
  assign _EVAL_2094 = _EVAL_151 == 12'hc87;
  assign _EVAL_977 = _EVAL_1224 & _EVAL_2156;
  assign _EVAL_1353 = _EVAL_1224 & _EVAL_1147;
  assign _EVAL_1711 = ~_EVAL_121;
  assign _EVAL_786 = _EVAL_2371 & _EVAL_988;
  assign _EVAL_1814 = _EVAL_1224 & _EVAL_1154;
  assign _EVAL_1089 = _EVAL_2167 & _EVAL_1106;
  assign _EVAL_1703 = _EVAL_151 == 12'hb19;
  assign _EVAL_229 = _EVAL_1224 & _EVAL_973;
  assign _EVAL_1078 = _EVAL_2371 & _EVAL_1188;
  assign _EVAL_2194 = _EVAL_1224 & _EVAL_1702;
  assign _EVAL_1403 = _EVAL_2167 & _EVAL_1559;
  assign _EVAL_984 = _EVAL_1224 & _EVAL_1842;
  assign _EVAL_1197 = _EVAL_151 == 12'h3b8;
  assign _EVAL_923 = _EVAL_1224 & _EVAL_1084;
  assign _EVAL_992 = _EVAL_151 == 12'hb9e;
  assign _EVAL_2050 = _EVAL_2167 & _EVAL_1480;
  assign _EVAL_309 = _EVAL_1224 & _EVAL_1864;
  assign _EVAL_1578 = _EVAL_2167 & _EVAL_1325;
  assign _EVAL_1902 = _EVAL_151 == 12'hb09;
  assign _EVAL_2161 = _EVAL_2167 & _EVAL_1176;
  assign _EVAL_2424 = _EVAL_151 == 12'h331;
  assign _EVAL_950 = _EVAL_1224 & _EVAL_1912;
  assign _EVAL_411 = _EVAL_151 == 12'h32c;
  assign _EVAL_2235 = _EVAL_151 == 12'hb1e;
  assign _EVAL_2205 = _EVAL_151 == 12'hb99;
  assign _EVAL_1464 = _EVAL_1224 & _EVAL_2364;
  assign _EVAL_261 = _EVAL_1224 & _EVAL_1311;
  assign _EVAL_1226 = _EVAL_1224 & _EVAL_802;
  assign _EVAL_738 = _EVAL_1224 & _EVAL_1026;
  assign _EVAL_226 = _EVAL_151 == 12'hc94;
  assign _EVAL_2523 = _EVAL_531 == 32'h80000010;
  assign _EVAL_2136 = _EVAL_151 == 12'hc1b;
  assign _EVAL_2408 = _EVAL_1224 & _EVAL_1656;
  assign _EVAL_1292 = _EVAL_531 == 32'h0;
  assign _EVAL_1225 = _EVAL_151 == 12'h33d;
  assign _EVAL_2380 = _EVAL_151 == 12'hc0a;
  assign _EVAL_1408 = _EVAL_151 == 12'h32f;
  assign _EVAL_839 = _EVAL_151 == 12'hb05;
  assign _EVAL_2224 = _EVAL_1224 & _EVAL_1769;
  assign _EVAL_940 = _EVAL_1224 & _EVAL_766;
  assign _EVAL_344 = _EVAL_2167 & _EVAL_2360;
  assign _EVAL_2204 = _EVAL_1224 & _EVAL_954;
  assign _EVAL_489 = _EVAL_1224 & _EVAL_1307;
  assign _EVAL_1747 = _EVAL_151 == 12'hc09;
  assign _EVAL_1491 = _EVAL_1224 & _EVAL_419;
  assign _EVAL_1605 = _EVAL_151 == 12'hb06;
  assign _EVAL_2156 = _EVAL_151 == 12'h33a;
  assign _EVAL_693 = _EVAL_151 == 12'hc93;
  assign _EVAL_1965 = _EVAL_1224 & _EVAL_2459;
  assign _EVAL_1295 = _EVAL_1224 & _EVAL_1225;
  assign _EVAL_331 = _EVAL_151 == 12'hc05;
  assign _EVAL_2375 = _EVAL_151 == 12'hb95;
  assign _EVAL_1523 = _EVAL_1224 & _EVAL_1839;
  assign _EVAL_1626 = _EVAL_151 == 12'hb1b;
  assign _EVAL_1726 = _EVAL_151 == 12'hb94;
  assign _EVAL_2019 = _EVAL_151 == 12'hc88;
  assign _EVAL_1093 = _EVAL_2167 & _EVAL_2300;
  assign _EVAL_2100 = _EVAL_151 == 12'hb1f;
  assign _EVAL_1570 = _EVAL_1224 & _EVAL_1917;
  assign _EVAL_948 = _EVAL_1224 & _EVAL_1039;
  assign _EVAL_1188 = _EVAL_531 == 32'h80000014;
  assign _EVAL_1400 = _EVAL_1224 & _EVAL_2237;
  assign _EVAL_1232 = _EVAL_1224 & _EVAL_2240;
  assign _EVAL_328 = _EVAL_1224 & _EVAL_1323;
  assign _EVAL_1106 = _EVAL_151 == 12'hc1e;
  assign _EVAL_1611 = _EVAL_1224 & _EVAL_2317;
  assign _EVAL_1055 = _EVAL_1224 & _EVAL_206;
  assign _EVAL_2233 = _EVAL_1224 & _EVAL_2246;
  assign _EVAL_1162 = _EVAL_1224 & _EVAL_2447;
  assign _EVAL_1868 = _EVAL_531 == 32'h1;
  assign _EVAL_518 = _EVAL_531 == 32'h8;
  assign _EVAL_2040 = _EVAL_151 == 12'hc15;
  assign _EVAL_716 = _EVAL_1224 & _EVAL_1019;
  assign _EVAL_2438 = _EVAL_2371 & _EVAL_2261;
  assign _EVAL_1390 = _EVAL_1224 & _EVAL_1317;
  assign _EVAL_2545 = _EVAL_1224 & _EVAL_2100;
  assign _EVAL_1469 = _EVAL_151 == 12'hc8b;
  assign _EVAL_1173 = _EVAL_1224 & _EVAL_1152;
  assign _EVAL_1552 = _EVAL_1224 & _EVAL_374;
  assign _EVAL_1774 = _EVAL_2167 & _EVAL_2395;
  assign _EVAL_677 = _EVAL_1224 & _EVAL_522;
  assign _EVAL_751 = _EVAL_2167 & _EVAL_2353;
  assign _EVAL_761 = _EVAL_2371 & _EVAL_1895;
  assign _EVAL_719 = _EVAL_151 == 12'hc9e;
  assign _EVAL_1021 = _EVAL_151 == 12'h336;
  assign _EVAL_276 = _EVAL_151 == 12'hc0b;
  assign _EVAL_812 = _EVAL_2167 & _EVAL_453;
  assign _EVAL_1352 = _EVAL_151 == 12'hb17;
  assign _EVAL_988 = _EVAL_531 == 32'h80000016;
  assign _EVAL_1853 = _EVAL_1224 & _EVAL_1242;
  assign _EVAL_1185 = _EVAL_151 == 12'hc0e;
  assign _EVAL_1538 = _EVAL_531 == 32'h8000001c;
  assign _EVAL_1986 = _EVAL_2167 & _EVAL_2264;
  assign _EVAL_203 = _EVAL_1224 & _EVAL_2375;
  assign _EVAL_1917 = _EVAL_151 == 12'hb8b;
  assign _EVAL_255 = _EVAL_2167 & _EVAL_1975;
  assign _EVAL_1368 = _EVAL_1224 & _EVAL_1197;
  assign _EVAL_1674 = _EVAL_1224 & _EVAL_2152;
  assign _EVAL_371 = _EVAL_151 == 12'hb8d;
  assign _EVAL_752 = _EVAL_1224 & _EVAL_1591;
  assign _EVAL_2106 = _EVAL_2371 & _EVAL_1617;
  assign _EVAL_1434 = _EVAL_531 == 32'h8000001a;
  assign _EVAL_1743 = _EVAL_1224 & _EVAL_2406;
  assign _EVAL_1900 = _EVAL_2371 & _EVAL_1538;
  assign _EVAL_1555 = _EVAL_151 == 12'hc14;
  assign _EVAL_822 = _EVAL_2167 & _EVAL_2407;
  assign _EVAL_1152 = _EVAL_151 == 12'hb0a;
  assign _EVAL_2152 = _EVAL_151 == 12'h3bb;
  assign _EVAL_1624 = _EVAL_151 == 12'h3bf;
  assign _EVAL_1263 = _EVAL_2371 & _EVAL_976;
  assign _EVAL_496 = _EVAL_151 == 12'h3a2;
  always @(posedge _EVAL_85) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_425 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f84b05d9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1982 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b2726d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_812 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(764187b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2383 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(335f766)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_669 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20e70115)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_309 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e4604e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_868 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22df21b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1207 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4aba384)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1552 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(726cc0da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_255 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d748031)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1965 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1eb2b846)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1127 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74e86945)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1267 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc52034f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2351 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2806e57)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_664 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae8e1cfb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2050 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edd6c590)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1774 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8c5c571)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2254 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d73f28ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1743 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42ab6615)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1837 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(512ed5ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_633 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26729c7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1811 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(737126bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1853 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(886b2072)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_458 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(afc44063)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1831 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a6e523)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1011 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f089853c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1368 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43e57488)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_786 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91791f0d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_467 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c120a9a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1784 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6a76e33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2068 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d98896e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1900 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51633608)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6af9aeed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1278 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d1738fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1237 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ad862db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_984 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f3d2808)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1387 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acef0569)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1932 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(642c7a43)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1004 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37093cd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_746 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a967d8e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_950 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98f13e34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1236 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d1da3cf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_822 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c4e77f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1840 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68090aeb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1268 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd43f5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1570 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17fc107c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_557 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8cdcb8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2097 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3828c185)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1585 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66d9cf17)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2499 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ebe0e95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_978 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7938427c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1578 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b46589cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_605 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(785126c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1184 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea505b2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2230 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e74656a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_344 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6534624)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1162 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62217d01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_814 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2de43d36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2453 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e281f46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2273) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da5544ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_698 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c6a8d15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_578 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fb2ecea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_433 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cec69e91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2231 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3292875)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2111 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(337522a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1530 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a34a42e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_538 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8608171)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2203 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ebea2fde)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1572 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c773c916)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1523 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80a4c0d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1653 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb66077e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2233 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44dbabfa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_887 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2a359ad4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1253 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17bba47d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1156 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7067a4eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1426 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45033694)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_813 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6e8c2a2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1403 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9208d41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2286 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98dc99b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1649 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66abcdc4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_908 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6bc21bd0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1650 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce9252b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_777 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(519cd61b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2509 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6adab0c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2081 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e93988c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1611 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72ebde33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90c4ac00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2370 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ffc7a30)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1044 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f20e67f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1375 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99097f20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1508 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9edea95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_678 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b77184d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1008 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98d88f48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_716 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99a9afcc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_750 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8011213b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1746 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b33428d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1674 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6cf461d2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1960 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff2b2a6b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_827 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4ce748d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1815 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8331b75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1247 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7eb799cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_946 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c9cbc80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_977 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c772110)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_826 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21d120d0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_296 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4577228)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2443 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d63667d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1462 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(554caf67)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_269 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c2d9f8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1713 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f2e8b53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35353d59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_761 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d9d4e7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_680 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(426741ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f9404a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1491 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b484d99e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_808 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6985cde)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1361 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4eefef2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2008 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89d20906)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_399 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67d75aed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1089 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(330c45e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_940 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5781752c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_982 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9e0c12e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2408 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdd77c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2438 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f277be5d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_352 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d3228a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1390 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f923ebce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_944) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfe5b6f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1632 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(caaae516)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_609 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52d5ab34)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1548 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d3f88c05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1115 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dbed7d2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2293 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bcb75772)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1234 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fef17256)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1666 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8fa4a617)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2299 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d91969ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_301 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25a80b6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2204 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac45bcdd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1542 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21589658)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_203 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(900006)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_636 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6d61460)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_948 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(281e91a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1397 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af463046)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1108 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(64711323)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1165 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9f4160f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1199 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edd48634)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2288 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7767f941)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1365 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd8b7535)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_656 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(102b348a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_806 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c267f081)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2464 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49db05c5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1158 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aea19b47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2545 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0854792)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_758 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bdc4da1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1173 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5f5ab85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_762 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54aa10e3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_742 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17bd09a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_544 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6db81552)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1263 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3426d500)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_764 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c78037)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_292 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c30fd74e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1814 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27bba281)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1241 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86159789)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2302 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c686f2be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2373 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(360a6e9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_211 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba3c5813)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_613 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f3b189)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_475 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82682a37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1226 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45f1c3e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1296 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec6c77c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_339 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1848f209)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1671 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3638ba6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2083 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89df614e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2236 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ea3626d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_884 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e316c29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1055 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb830853)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1400 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d0e41e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_510 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(da5e25f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1433 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81e3cd9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_586 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ddd3f597)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_752 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9cead198)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_987 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46628290)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1353 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eef2ac3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1232 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b5dbf2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2224 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43c79d32)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1356 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21d88f0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_229 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb5dff89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1295 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66718dad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2533 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1809e108)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1763 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9bc9723)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_2273) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1054 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9f13409)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_328 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(856403fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1507 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c38b4239)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_219 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f188f99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1846 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b38ef71f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_335 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9837641)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1464 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8b5bd02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_998 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4283f64)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_285 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(878eb186)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2324 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7040ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1466 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72845d46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_751 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d66435f7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2161 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b475bcb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1257 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(684adf3e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_489 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5fb8c7f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_677 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b02c8397)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1908 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4e5f55e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1093 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b98e4ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_944) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_261 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc13b121)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1272 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ecea8b6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_923 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(909530d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1020 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c8c45ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_603 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42c4e4f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_794 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d2ca5ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2106 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0ba42c4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1973 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52722d82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2348 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a79f34e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_738 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(125af846)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_864 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c67d483d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1979 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cff4640d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_290 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51fa7676)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1166 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1612798)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1986 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85861249)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1138 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4372647b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_953 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2ec65ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1638 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(661a21f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2450 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3948ccbf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_266 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95f890d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1078 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(466af74c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_574 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab7bbd55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_520 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(920dd457)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_588 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e8c4406)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2194 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(123d2eb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1134 & _EVAL_774) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28232492)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
