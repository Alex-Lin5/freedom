//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_99_assert(
  input           _EVAL_5,
  input  [2:0]    _EVAL_6,
  input           _EVAL_9,
  input  [1:0]    _EVAL_17,
  input  [2:0]    _EVAL_70,
  input  [9:0]    _EVAL_73,
  input  [3:0]    _EVAL_84,
  input           _EVAL_110,
  input           _EVAL_119,
  input  [27:0]   _EVAL_130,
  input           _EVAL_136,
  input           _EVAL_151,
  input           _EVAL_160,
  input           _EVAL_180,
  input           _EVAL_184,
  input           _EVAL_205,
  input           _EVAL_212,
  input           _EVAL_213,
  input           _EVAL_223,
  input           _EVAL_244,
  input           _EVAL_259,
  input           _EVAL_275,
  input           _EVAL_288,
  input           _EVAL_294,
  input           _EVAL_295,
  input           _EVAL_300,
  input  [126:0]  _EVAL_304,
  input           _EVAL_320,
  input           _EVAL_333,
  input           _EVAL_335,
  input           _EVAL_338,
  input           _EVAL_340,
  input           _EVAL_356,
  input           _EVAL_365,
  input           _EVAL_367,
  input           _EVAL_369,
  input           _EVAL_379,
  input           _EVAL_402,
  input           _EVAL_403,
  input           _EVAL_416,
  input           _EVAL_463,
  input  [7:0]    _EVAL_469,
  input           _EVAL_485,
  input           _EVAL_489,
  input           _EVAL_506,
  input           _EVAL_509,
  input           _EVAL_510,
  input           _EVAL_515,
  input           _EVAL_533,
  input           _EVAL_560,
  input           _EVAL_575,
  input           _EVAL_590,
  input           _EVAL_604,
  input           _EVAL_613,
  input           _EVAL_625,
  input           _EVAL_632,
  input           _EVAL_640,
  input  [1023:0] _EVAL_651,
  input           _EVAL_652,
  input           _EVAL_687,
  input           _EVAL_693,
  input           _EVAL_697,
  input           _EVAL_709,
  input           _EVAL_715,
  input           _EVAL_723,
  input           _EVAL_741,
  input           _EVAL_765,
  input           _EVAL_772,
  input           _EVAL_777,
  input           _EVAL_794,
  input           _EVAL_796,
  input           _EVAL_799,
  input           _EVAL_817,
  input           _EVAL_826,
  input           _EVAL_837,
  input           _EVAL_838,
  input           _EVAL_840,
  input           _EVAL_844,
  input           _EVAL_851,
  input           _EVAL_862,
  input           _EVAL_868,
  input           _EVAL_871,
  input           _EVAL_903,
  input           _EVAL_908,
  input           _EVAL_917,
  input           _EVAL_1012,
  input  [7:0]    _EVAL_1016,
  input           _EVAL_1022,
  input           _EVAL_1051,
  input           _EVAL_1053,
  input           _EVAL_1057,
  input           _EVAL_1066,
  input           _EVAL_1086,
  input           _EVAL_1090,
  input           _EVAL_1094,
  input           _EVAL_1103,
  input           _EVAL_1135,
  input           _EVAL_1146,
  input           _EVAL_1164,
  input           _EVAL_1170,
  input           _EVAL_1202,
  input           _EVAL_1218,
  input           _EVAL_1248,
  input           _EVAL_1250,
  input           _EVAL_1263,
  input           _EVAL_1267,
  input           _EVAL_1280,
  input           _EVAL_1301,
  input           _EVAL_1304,
  input           _EVAL_1311,
  input           _EVAL_1320,
  input           _EVAL_1328,
  input           _EVAL_1338,
  input           _EVAL_1354,
  input           _EVAL_1371,
  input           _EVAL_1396,
  input           _EVAL_1401,
  input           _EVAL_1426,
  input           _EVAL_1444,
  input           _EVAL_1476,
  input           _EVAL_1486,
  input           _EVAL_1505,
  input           _EVAL_1521,
  input           _EVAL_1532,
  input           _EVAL_1535,
  input           _EVAL_1539,
  input           _EVAL_1544,
  input           _EVAL_1560,
  input           _EVAL_1591,
  input           _EVAL_1596,
  input           _EVAL_1613,
  input           _EVAL_1644,
  input           _EVAL_1649,
  input           _EVAL_1662,
  input           _EVAL_1664,
  input           _EVAL_1712,
  input           _EVAL_1715,
  input           _EVAL_1720,
  input           _EVAL_1729,
  input           _EVAL_1731,
  input           _EVAL_1750,
  input           _EVAL_1755,
  input           _EVAL_1763,
  input           _EVAL_1769,
  input           _EVAL_1780,
  input           _EVAL_1787,
  input           _EVAL_1793,
  input           _EVAL_1797,
  input           _EVAL_1830,
  input           _EVAL_1852,
  input           _EVAL_1875,
  input           _EVAL_1877,
  input           _EVAL_1886,
  input           _EVAL_1896,
  input           _EVAL_1904,
  input           _EVAL_1905,
  input           _EVAL_1942,
  input           _EVAL_1953,
  input           _EVAL_1956,
  input           _EVAL_1972,
  input           _EVAL_1973,
  input           _EVAL_2011,
  input           _EVAL_2015,
  input           _EVAL_2027,
  input           _EVAL_2054,
  input  [2:0]    _EVAL_2084,
  input           _EVAL_2087,
  input           _EVAL_2097,
  input           _EVAL_2103,
  input           _EVAL_2113,
  input           _EVAL_2119,
  input           _EVAL_2123,
  input           _EVAL_2142,
  input           _EVAL_2152,
  input           _EVAL_2168,
  input           _EVAL_2190,
  input           _EVAL_2198,
  input           _EVAL_2206,
  input           _EVAL_2220,
  input           _EVAL_2224,
  input           _EVAL_2233,
  input           _EVAL_2234,
  input           _EVAL_2270,
  input  [126:0]  _EVAL_2296,
  input           _EVAL_2318,
  input           _EVAL_2327,
  input           _EVAL_2328,
  input           _EVAL_2329,
  input           _EVAL_2346,
  input           _EVAL_2362,
  input           _EVAL_2375,
  input           _EVAL_2403,
  input           _EVAL_2406,
  input           _EVAL_2410,
  input           _EVAL_2425,
  input           _EVAL_2454,
  input  [25:0]   _EVAL_2478,
  input           _EVAL_2484,
  input           _EVAL_2494,
  input           _EVAL_2499,
  input           _EVAL_2511,
  input           _EVAL_2577,
  input           _EVAL_2615,
  input           _EVAL_2623,
  input           _EVAL_2624,
  input           _EVAL_2633,
  input           _EVAL_2651,
  input           _EVAL_2658,
  input           _EVAL_2661,
  input           _EVAL_2689,
  input           _EVAL_2733,
  input           _EVAL_2734,
  input           _EVAL_2747,
  input           _EVAL_2756,
  input  [6:0]    _EVAL_2757,
  input           _EVAL_2773,
  input           _EVAL_2774,
  input           _EVAL_2795,
  input           _EVAL_2798,
  input           _EVAL_2814,
  input           _EVAL_2846,
  input  [31:0]   _EVAL_2850,
  input           _EVAL_2855,
  input           _EVAL_2865,
  input           _EVAL_2874,
  input           _EVAL_2879,
  input           _EVAL_2906,
  input  [7:0]    _EVAL_2914,
  input           _EVAL_2919,
  input           _EVAL_2945,
  input           _EVAL_2952,
  input           _EVAL_2963,
  input           _EVAL_2983,
  input           _EVAL_2990,
  input           _EVAL_3008,
  input           _EVAL_3036,
  input  [7:0]    _EVAL_3038,
  input           _EVAL_3056,
  input           _EVAL_3064,
  input           _EVAL_3068,
  input           _EVAL_3097,
  input           _EVAL_3099,
  input           _EVAL_3133,
  input           _EVAL_3148,
  input  [2:0]    _EVAL_3156,
  input           _EVAL_3165,
  input           _EVAL_3167,
  input           _EVAL_3179,
  input           _EVAL_3182,
  input           _EVAL_3206,
  input           _EVAL_3211,
  input           _EVAL_3223,
  input           _EVAL_3243,
  input           _EVAL_3249,
  input           _EVAL_3255,
  input           _EVAL_3286,
  input           _EVAL_3287,
  input           _EVAL_3319,
  input           _EVAL_3321,
  input           _EVAL_3339,
  input           _EVAL_3343,
  input           _EVAL_3347,
  input           _EVAL_3359,
  input           _EVAL_3368,
  input           _EVAL_3384,
  input           _EVAL_3390,
  input           _EVAL_3408,
  input           _EVAL_3410,
  input           _EVAL_3414,
  input           _EVAL_3435,
  input           _EVAL_3443,
  input           _EVAL_3456,
  input           _EVAL_3462,
  input           _EVAL_3489,
  input           _EVAL_3494,
  input           _EVAL_3519,
  input           _EVAL_3524,
  input           _EVAL_3555,
  input           _EVAL_3572,
  input           _EVAL_3588,
  input           _EVAL_3619,
  input           _EVAL_3622,
  input           _EVAL_3637,
  input           _EVAL_3651,
  input           _EVAL_3662,
  input           _EVAL_3672,
  input           _EVAL_3681,
  input           _EVAL_3696,
  input           _EVAL_3701,
  input  [6:0]    _EVAL_3702,
  input           _EVAL_3715,
  input           _EVAL_3717,
  input           _EVAL_3719,
  input           _EVAL_3720,
  input           _EVAL_3722,
  input           _EVAL_3729,
  input           _EVAL_3732,
  input           _EVAL_3735,
  input           _EVAL_3745,
  input           _EVAL_3747,
  input           _EVAL_3757,
  input           _EVAL_3787,
  input           _EVAL_3806,
  input           _EVAL_3809,
  input           _EVAL_3840,
  input           _EVAL_3852,
  input           out_back__EVAL_7,
  input  [9:0]    out_back__EVAL_11,
  input           out_back__EVAL_2,
  input  [1:0]    out_back__EVAL_6
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_145;
  wire  _EVAL_147;
  wire  _EVAL_149;
  wire  _EVAL_152;
  wire  _EVAL_154;
  wire [126:0] _EVAL_155;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_169;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_178;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire [7:0] _EVAL_194;
  wire [126:0] _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_204;
  wire  _EVAL_207;
  wire  _EVAL_211;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_226;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_237;
  wire  _EVAL_239;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_246;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_255;
  wire  _EVAL_260;
  wire  _EVAL_261;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_266;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_271;
  wire  _EVAL_277;
  wire  _EVAL_283;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_303;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_307;
  wire  _EVAL_308;
  wire  _EVAL_310;
  wire  _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire  _EVAL_319;
  wire  _EVAL_327;
  wire  _EVAL_328;
  wire  _EVAL_329;
  wire  _EVAL_332;
  wire  _EVAL_345;
  wire  _EVAL_346;
  wire  _EVAL_347;
  wire  _EVAL_348;
  wire  _EVAL_349;
  wire  _EVAL_351;
  wire  _EVAL_352;
  wire  _EVAL_357;
  wire  _EVAL_358;
  wire  _EVAL_359;
  wire  _EVAL_360;
  wire  _EVAL_361;
  wire  _EVAL_363;
  wire  _EVAL_370;
  wire  _EVAL_372;
  wire  _EVAL_373;
  wire  _EVAL_375;
  wire  _EVAL_376;
  wire  _EVAL_377;
  wire  _EVAL_380;
  wire  _EVAL_387;
  wire  _EVAL_388;
  wire  _EVAL_389;
  wire  _EVAL_391;
  wire  _EVAL_392;
  wire  _EVAL_393;
  wire  _EVAL_395;
  wire  _EVAL_397;
  wire  _EVAL_398;
  wire  _EVAL_399;
  wire  _EVAL_400;
  wire  _EVAL_401;
  wire  _EVAL_405;
  wire  _EVAL_406;
  wire  _EVAL_407;
  wire  _EVAL_409;
  wire  _EVAL_413;
  wire  _EVAL_417;
  wire  _EVAL_418;
  wire  _EVAL_419;
  wire  _EVAL_420;
  wire  _EVAL_424;
  wire  _EVAL_426;
  wire  _EVAL_430;
  wire  _EVAL_431;
  wire  _EVAL_432;
  wire  _EVAL_433;
  wire  _EVAL_436;
  wire  _EVAL_438;
  wire  _EVAL_439;
  wire  _EVAL_441;
  wire  _EVAL_442;
  wire  _EVAL_443;
  wire  _EVAL_444;
  wire  _EVAL_447;
  wire  _EVAL_448;
  wire  _EVAL_452;
  wire  _EVAL_453;
  wire [7:0] _EVAL_454;
  wire  _EVAL_455;
  wire  _EVAL_457;
  wire  _EVAL_459;
  wire [7:0] _EVAL_460;
  wire  _EVAL_464;
  wire  _EVAL_465;
  wire  _EVAL_470;
  wire  _EVAL_472;
  wire  _EVAL_474;
  wire  _EVAL_475;
  wire  _EVAL_477;
  wire  _EVAL_479;
  wire  _EVAL_481;
  wire  _EVAL_483;
  wire  _EVAL_484;
  wire  _EVAL_486;
  wire  _EVAL_491;
  wire  _EVAL_493;
  wire  _EVAL_494;
  wire  _EVAL_497;
  wire  _EVAL_501;
  wire  _EVAL_502;
  wire  _EVAL_503;
  wire  _EVAL_507;
  wire  _EVAL_508;
  wire  _EVAL_511;
  wire  _EVAL_512;
  wire  _EVAL_514;
  wire  _EVAL_519;
  wire  _EVAL_521;
  wire  _EVAL_522;
  wire  _EVAL_523;
  wire  _EVAL_525;
  wire  _EVAL_527;
  wire  _EVAL_528;
  wire  _EVAL_530;
  wire  _EVAL_535;
  wire  _EVAL_537;
  wire  _EVAL_538;
  wire  _EVAL_539;
  wire  _EVAL_541;
  wire  _EVAL_542;
  wire  _EVAL_543;
  wire  _EVAL_545;
  wire  _EVAL_546;
  wire  _EVAL_548;
  wire  _EVAL_549;
  wire  _EVAL_550;
  wire  _EVAL_551;
  wire [19:0] _EVAL_553;
  wire  _EVAL_554;
  wire  _EVAL_555;
  wire  _EVAL_556;
  wire  _EVAL_557;
  wire  _EVAL_558;
  wire  _EVAL_559;
  wire  _EVAL_561;
  wire  _EVAL_562;
  wire  _EVAL_563;
  wire  _EVAL_564;
  wire  _EVAL_565;
  wire  _EVAL_568;
  wire  _EVAL_572;
  wire  _EVAL_574;
  wire  _EVAL_577;
  wire  _EVAL_578;
  wire  _EVAL_579;
  wire  _EVAL_580;
  wire  _EVAL_581;
  wire  _EVAL_586;
  wire  _EVAL_587;
  wire  _EVAL_589;
  wire  _EVAL_591;
  wire  _EVAL_596;
  wire  _EVAL_597;
  wire  _EVAL_598;
  wire  _EVAL_599;
  wire  _EVAL_601;
  wire  _EVAL_606;
  wire  _EVAL_608;
  wire  _EVAL_611;
  wire  _EVAL_617;
  wire  _EVAL_618;
  wire  _EVAL_619;
  wire  _EVAL_620;
  wire  _EVAL_621;
  wire  _EVAL_622;
  wire  _EVAL_623;
  wire  _EVAL_624;
  wire  _EVAL_626;
  wire  _EVAL_629;
  wire  _EVAL_633;
  wire  _EVAL_634;
  wire  _EVAL_635;
  wire  _EVAL_636;
  wire  _EVAL_637;
  wire  _EVAL_649;
  wire  _EVAL_650;
  wire  _EVAL_654;
  wire  _EVAL_656;
  wire  _EVAL_658;
  wire  _EVAL_659;
  wire  _EVAL_661;
  wire  _EVAL_662;
  wire  _EVAL_663;
  wire  _EVAL_664;
  wire  _EVAL_665;
  wire  _EVAL_666;
  wire  _EVAL_671;
  wire  _EVAL_674;
  wire  _EVAL_675;
  wire  _EVAL_676;
  wire  _EVAL_680;
  wire  _EVAL_681;
  wire  _EVAL_682;
  wire  _EVAL_684;
  wire  _EVAL_686;
  wire  _EVAL_690;
  wire  _EVAL_694;
  wire  _EVAL_698;
  wire  _EVAL_701;
  wire  _EVAL_702;
  wire  _EVAL_704;
  wire  _EVAL_705;
  wire  _EVAL_706;
  wire  _EVAL_708;
  wire  _EVAL_711;
  wire  _EVAL_713;
  wire  _EVAL_714;
  wire  _EVAL_716;
  wire  _EVAL_717;
  wire  _EVAL_718;
  wire  _EVAL_720;
  wire  _EVAL_722;
  wire  _EVAL_724;
  wire  _EVAL_725;
  wire  _EVAL_728;
  wire  _EVAL_729;
  wire  _EVAL_730;
  wire  _EVAL_731;
  wire  _EVAL_734;
  wire  _EVAL_737;
  wire  _EVAL_738;
  wire  _EVAL_740;
  wire  _EVAL_742;
  wire  _EVAL_745;
  wire  _EVAL_746;
  wire  _EVAL_747;
  wire  _EVAL_748;
  wire  _EVAL_749;
  wire  _EVAL_750;
  wire  _EVAL_754;
  wire  _EVAL_756;
  wire  _EVAL_757;
  wire  _EVAL_760;
  wire  _EVAL_761;
  wire  _EVAL_763;
  wire  _EVAL_764;
  wire  _EVAL_766;
  wire  _EVAL_767;
  wire  _EVAL_768;
  wire  _EVAL_769;
  wire  _EVAL_773;
  wire  _EVAL_774;
  wire  _EVAL_781;
  wire  _EVAL_785;
  wire  _EVAL_786;
  wire  _EVAL_788;
  wire  _EVAL_790;
  wire  _EVAL_791;
  wire  _EVAL_795;
  wire  _EVAL_798;
  wire  _EVAL_800;
  wire  _EVAL_802;
  wire  _EVAL_803;
  wire  _EVAL_805;
  wire  _EVAL_806;
  wire  _EVAL_807;
  wire  _EVAL_812;
  wire  _EVAL_814;
  wire  _EVAL_816;
  wire  _EVAL_818;
  wire  _EVAL_821;
  wire  _EVAL_822;
  wire  _EVAL_823;
  wire  _EVAL_824;
  wire  _EVAL_825;
  wire  _EVAL_829;
  wire  _EVAL_830;
  wire  _EVAL_831;
  wire  _EVAL_833;
  wire  _EVAL_835;
  wire  _EVAL_836;
  wire  _EVAL_839;
  wire  _EVAL_843;
  wire  _EVAL_846;
  wire  _EVAL_852;
  wire  _EVAL_857;
  wire  _EVAL_861;
  wire  _EVAL_863;
  wire  _EVAL_864;
  wire  _EVAL_866;
  wire  _EVAL_867;
  wire  _EVAL_874;
  wire  _EVAL_875;
  wire  _EVAL_877;
  wire  _EVAL_878;
  wire  _EVAL_879;
  wire  _EVAL_881;
  wire  _EVAL_882;
  wire  _EVAL_883;
  wire  _EVAL_884;
  wire  _EVAL_885;
  wire  _EVAL_887;
  wire  _EVAL_888;
  wire  _EVAL_891;
  wire  _EVAL_893;
  wire  _EVAL_895;
  wire  _EVAL_896;
  wire  _EVAL_897;
  wire  _EVAL_898;
  wire  _EVAL_900;
  wire  _EVAL_901;
  wire  _EVAL_912;
  wire  _EVAL_914;
  wire [126:0] _EVAL_915;
  wire  _EVAL_919;
  wire  _EVAL_920;
  wire  _EVAL_922;
  wire  _EVAL_923;
  wire  _EVAL_924;
  wire  _EVAL_926;
  wire  _EVAL_927;
  wire  _EVAL_928;
  wire  _EVAL_929;
  wire  _EVAL_931;
  wire  _EVAL_932;
  wire  _EVAL_934;
  wire  _EVAL_935;
  wire  _EVAL_938;
  wire  _EVAL_940;
  wire  _EVAL_941;
  wire  _EVAL_942;
  wire  _EVAL_943;
  wire  _EVAL_945;
  wire  _EVAL_946;
  wire  _EVAL_947;
  wire  _EVAL_948;
  wire  _EVAL_950;
  wire  _EVAL_951;
  wire  _EVAL_952;
  wire  _EVAL_958;
  wire  _EVAL_960;
  wire  _EVAL_961;
  wire  _EVAL_968;
  wire  _EVAL_969;
  wire  _EVAL_971;
  wire  _EVAL_972;
  wire  _EVAL_974;
  wire  _EVAL_976;
  wire  _EVAL_977;
  wire  _EVAL_981;
  wire  _EVAL_983;
  wire  _EVAL_984;
  wire  _EVAL_985;
  wire  _EVAL_986;
  wire  _EVAL_993;
  wire  _EVAL_998;
  wire  _EVAL_999;
  wire  _EVAL_1001;
  wire  _EVAL_1003;
  wire  _EVAL_1004;
  wire  _EVAL_1006;
  wire  _EVAL_1007;
  wire  _EVAL_1013;
  wire  _EVAL_1018;
  wire  _EVAL_1019;
  wire  _EVAL_1025;
  wire  _EVAL_1027;
  wire  _EVAL_1028;
  wire  _EVAL_1029;
  wire  _EVAL_1035;
  wire  _EVAL_1037;
  wire  _EVAL_1038;
  wire  _EVAL_1042;
  wire  _EVAL_1044;
  wire  _EVAL_1045;
  wire  _EVAL_1047;
  wire  _EVAL_1048;
  wire  _EVAL_1049;
  wire  _EVAL_1050;
  wire  _EVAL_1054;
  wire  _EVAL_1055;
  wire  _EVAL_1058;
  wire  _EVAL_1059;
  wire [7:0] _EVAL_1060;
  wire  _EVAL_1063;
  wire  _EVAL_1064;
  wire  _EVAL_1067;
  wire  _EVAL_1068;
  wire  _EVAL_1069;
  wire  _EVAL_1070;
  wire  _EVAL_1075;
  wire  _EVAL_1077;
  wire  _EVAL_1078;
  wire  _EVAL_1079;
  wire  _EVAL_1080;
  wire  _EVAL_1082;
  wire  _EVAL_1083;
  wire  _EVAL_1084;
  wire  _EVAL_1091;
  wire  _EVAL_1092;
  wire  _EVAL_1095;
  wire  _EVAL_1097;
  wire  _EVAL_1098;
  wire  _EVAL_1100;
  wire  _EVAL_1104;
  wire  _EVAL_1105;
  wire  _EVAL_1106;
  wire  _EVAL_1107;
  wire  _EVAL_1108;
  wire  _EVAL_1109;
  wire  _EVAL_1110;
  wire  _EVAL_1111;
  wire  _EVAL_1113;
  wire  _EVAL_1114;
  wire  _EVAL_1115;
  wire  _EVAL_1119;
  wire  _EVAL_1121;
  wire  _EVAL_1123;
  wire  _EVAL_1125;
  wire  _EVAL_1126;
  wire  _EVAL_1128;
  wire  _EVAL_1129;
  wire  _EVAL_1131;
  wire  _EVAL_1132;
  wire  _EVAL_1136;
  wire  _EVAL_1137;
  wire  _EVAL_1139;
  wire  _EVAL_1141;
  wire  _EVAL_1142;
  wire  _EVAL_1145;
  wire  _EVAL_1149;
  wire  _EVAL_1150;
  wire  _EVAL_1152;
  wire  _EVAL_1154;
  wire  _EVAL_1155;
  wire  _EVAL_1156;
  wire  _EVAL_1157;
  wire  _EVAL_1159;
  wire  _EVAL_1160;
  wire  _EVAL_1161;
  wire  _EVAL_1162;
  wire  _EVAL_1163;
  wire  _EVAL_1165;
  wire  _EVAL_1166;
  wire  _EVAL_1168;
  wire  _EVAL_1169;
  wire  _EVAL_1173;
  wire  _EVAL_1176;
  wire  _EVAL_1177;
  wire  _EVAL_1179;
  wire  _EVAL_1186;
  wire  _EVAL_1188;
  wire  _EVAL_1189;
  wire  _EVAL_1192;
  wire  _EVAL_1194;
  wire  _EVAL_1196;
  wire  _EVAL_1197;
  wire  _EVAL_1198;
  wire  _EVAL_1201;
  wire  _EVAL_1204;
  wire  _EVAL_1205;
  wire  _EVAL_1206;
  wire  _EVAL_1207;
  wire  _EVAL_1210;
  wire  _EVAL_1212;
  wire  _EVAL_1213;
  wire  _EVAL_1214;
  wire  _EVAL_1215;
  wire  _EVAL_1216;
  wire  _EVAL_1217;
  wire  _EVAL_1219;
  wire  _EVAL_1223;
  wire  _EVAL_1225;
  wire  _EVAL_1226;
  wire  _EVAL_1227;
  wire  _EVAL_1228;
  wire  _EVAL_1229;
  wire  _EVAL_1230;
  wire  _EVAL_1231;
  wire  _EVAL_1232;
  wire  _EVAL_1233;
  wire  _EVAL_1234;
  wire  _EVAL_1235;
  wire  _EVAL_1236;
  wire  _EVAL_1240;
  wire  _EVAL_1242;
  wire  _EVAL_1244;
  wire  _EVAL_1245;
  wire [27:0] monitor__EVAL;
  wire  monitor__EVAL_0;
  wire  monitor__EVAL_1;
  wire [9:0] monitor__EVAL_2;
  wire [2:0] monitor__EVAL_3;
  wire [2:0] monitor__EVAL_4;
  wire  monitor__EVAL_5;
  wire [1:0] monitor__EVAL_6;
  wire [2:0] monitor__EVAL_7;
  wire [1:0] monitor__EVAL_8;
  wire [9:0] monitor__EVAL_9;
  wire  monitor__EVAL_10;
  wire  monitor__EVAL_11;
  wire  monitor__EVAL_12;
  wire [3:0] monitor__EVAL_13;
  wire  monitor__EVAL_14;
  wire  _EVAL_1246;
  wire  _EVAL_1247;
  wire  _EVAL_1249;
  wire  _EVAL_1253;
  wire  _EVAL_1256;
  wire  _EVAL_1258;
  wire  _EVAL_1259;
  wire  _EVAL_1260;
  wire  _EVAL_1261;
  wire  _EVAL_1265;
  wire  _EVAL_1266;
  wire  _EVAL_1271;
  wire  _EVAL_1272;
  wire  _EVAL_1273;
  wire  _EVAL_1275;
  wire  _EVAL_1276;
  wire  _EVAL_1277;
  wire  _EVAL_1279;
  wire  _EVAL_1284;
  wire  _EVAL_1285;
  wire  _EVAL_1287;
  wire  _EVAL_1289;
  wire  _EVAL_1290;
  wire  _EVAL_1291;
  wire  _EVAL_1294;
  wire  _EVAL_1295;
  wire  _EVAL_1296;
  wire  _EVAL_1297;
  wire  _EVAL_1298;
  wire  _EVAL_1300;
  wire  _EVAL_1302;
  wire  _EVAL_1305;
  wire  _EVAL_1306;
  wire  _EVAL_1309;
  wire  _EVAL_1312;
  wire  _EVAL_1313;
  wire  _EVAL_1316;
  wire  _EVAL_1317;
  wire  _EVAL_1318;
  wire  _EVAL_1319;
  wire  _EVAL_1321;
  wire  _EVAL_1322;
  wire  _EVAL_1324;
  wire  _EVAL_1326;
  wire  _EVAL_1327;
  wire  _EVAL_1330;
  wire  _EVAL_1331;
  wire  _EVAL_1332;
  wire  _EVAL_1335;
  wire  _EVAL_1337;
  wire  _EVAL_1344;
  wire  _EVAL_1345;
  wire  _EVAL_1348;
  wire  _EVAL_1351;
  wire  _EVAL_1352;
  wire  _EVAL_1353;
  wire  _EVAL_1355;
  wire  _EVAL_1356;
  wire  _EVAL_1357;
  wire  _EVAL_1360;
  wire [31:0] _EVAL_1361;
  wire  _EVAL_1362;
  wire  _EVAL_1363;
  wire  _EVAL_1370;
  wire  _EVAL_1372;
  wire  _EVAL_1373;
  wire  _EVAL_1375;
  wire  _EVAL_1376;
  wire  _EVAL_1377;
  wire  _EVAL_1378;
  wire  _EVAL_1381;
  wire  _EVAL_1383;
  wire  _EVAL_1384;
  wire  _EVAL_1386;
  wire  _EVAL_1387;
  wire  _EVAL_1388;
  wire  _EVAL_1389;
  wire  _EVAL_1390;
  wire  _EVAL_1391;
  wire  _EVAL_1393;
  wire  _EVAL_1394;
  wire  _EVAL_1397;
  wire  _EVAL_1399;
  wire  _EVAL_1402;
  wire  _EVAL_1403;
  wire  _EVAL_1404;
  wire  _EVAL_1405;
  wire  _EVAL_1406;
  wire  _EVAL_1409;
  wire  _EVAL_1410;
  wire  _EVAL_1412;
  wire  _EVAL_1414;
  wire  _EVAL_1416;
  wire  _EVAL_1420;
  wire  _EVAL_1421;
  wire  _EVAL_1423;
  wire  _EVAL_1424;
  wire  _EVAL_1425;
  wire  _EVAL_1427;
  wire  _EVAL_1429;
  wire  _EVAL_1431;
  wire  _EVAL_1432;
  wire  _EVAL_1436;
  wire  _EVAL_1437;
  wire  _EVAL_1442;
  wire  _EVAL_1445;
  wire  _EVAL_1453;
  wire  _EVAL_1454;
  wire  _EVAL_1455;
  wire [126:0] _EVAL_1456;
  wire  _EVAL_1457;
  wire  _EVAL_1458;
  wire  _EVAL_1460;
  wire  _EVAL_1461;
  wire  _EVAL_1462;
  wire  _EVAL_1463;
  wire [7:0] _EVAL_1464;
  wire  _EVAL_1465;
  wire  _EVAL_1468;
  wire  _EVAL_1469;
  wire  _EVAL_1470;
  wire  _EVAL_1474;
  wire  _EVAL_1475;
  wire  _EVAL_1477;
  wire  _EVAL_1478;
  wire  _EVAL_1479;
  wire  _EVAL_1484;
  wire  _EVAL_1487;
  wire  _EVAL_1490;
  wire  _EVAL_1491;
  wire  _EVAL_1492;
  wire  _EVAL_1493;
  wire  _EVAL_1494;
  wire  _EVAL_1495;
  wire  _EVAL_1497;
  wire  _EVAL_1501;
  wire  _EVAL_1502;
  wire  _EVAL_1503;
  wire  _EVAL_1508;
  wire  _EVAL_1511;
  wire  _EVAL_1513;
  wire  _EVAL_1514;
  wire  _EVAL_1515;
  wire  _EVAL_1519;
  wire  _EVAL_1522;
  wire  _EVAL_1523;
  wire  _EVAL_1525;
  wire  _EVAL_1526;
  wire  _EVAL_1530;
  wire  _EVAL_1531;
  wire  _EVAL_1533;
  wire  _EVAL_1538;
  wire  _EVAL_1543;
  wire  _EVAL_1545;
  wire  _EVAL_1546;
  wire  _EVAL_1551;
  wire  _EVAL_1552;
  wire  _EVAL_1553;
  wire  _EVAL_1556;
  wire  _EVAL_1557;
  wire  _EVAL_1558;
  wire  _EVAL_1559;
  wire  _EVAL_1561;
  wire  _EVAL_1562;
  wire  _EVAL_1563;
  wire  _EVAL_1566;
  wire  _EVAL_1567;
  wire  _EVAL_1570;
  wire  _EVAL_1571;
  wire  _EVAL_1572;
  wire  _EVAL_1573;
  wire  _EVAL_1574;
  wire  _EVAL_1575;
  wire  _EVAL_1577;
  wire  _EVAL_1580;
  reg  _EVAL_1581;
  wire  _EVAL_1582;
  wire  _EVAL_1583;
  wire  _EVAL_1584;
  wire  _EVAL_1585;
  wire  _EVAL_1586;
  wire  _EVAL_1588;
  wire  _EVAL_1589;
  wire  _EVAL_1590;
  wire  _EVAL_1598;
  wire  _EVAL_1599;
  wire  _EVAL_1600;
  wire  _EVAL_1602;
  wire  _EVAL_1603;
  wire  _EVAL_1606;
  wire  _EVAL_1609;
  wire  _EVAL_1611;
  wire  _EVAL_1612;
  wire  _EVAL_1614;
  wire  _EVAL_1615;
  wire  _EVAL_1616;
  wire  _EVAL_1619;
  wire  _EVAL_1620;
  wire  _EVAL_1625;
  wire  _EVAL_1626;
  wire  _EVAL_1628;
  wire  _EVAL_1629;
  wire  _EVAL_1632;
  wire  _EVAL_1633;
  wire  _EVAL_1635;
  wire  _EVAL_1636;
  wire  _EVAL_1639;
  wire  _EVAL_1640;
  wire  _EVAL_1641;
  wire  _EVAL_1642;
  wire  _EVAL_1643;
  wire  _EVAL_1646;
  wire  _EVAL_1648;
  wire  _EVAL_1650;
  wire  _EVAL_1651;
  wire  _EVAL_1652;
  wire  _EVAL_1653;
  wire  _EVAL_1654;
  wire  _EVAL_1656;
  wire  _EVAL_1660;
  wire  _EVAL_1663;
  wire  _EVAL_1665;
  wire  _EVAL_1667;
  wire  _EVAL_1668;
  wire  _EVAL_1669;
  wire  _EVAL_1671;
  wire  _EVAL_1672;
  wire  _EVAL_1676;
  wire  _EVAL_1679;
  wire  _EVAL_1682;
  wire  _EVAL_1685;
  wire  _EVAL_1686;
  wire  _EVAL_1690;
  wire  _EVAL_1691;
  wire  _EVAL_1693;
  wire  _EVAL_1699;
  wire  _EVAL_1701;
  wire  _EVAL_1704;
  wire  _EVAL_1705;
  wire  _EVAL_1708;
  wire  _EVAL_1709;
  wire  _EVAL_1713;
  wire  _EVAL_1714;
  wire  _EVAL_1716;
  wire  _EVAL_1717;
  wire  _EVAL_1719;
  wire  _EVAL_1721;
  wire  _EVAL_1724;
  wire  _EVAL_1725;
  wire  _EVAL_1726;
  wire  _EVAL_1727;
  wire  _EVAL_1728;
  wire  _EVAL_1730;
  wire  _EVAL_1732;
  wire  _EVAL_1734;
  wire  _EVAL_1735;
  wire  _EVAL_1736;
  wire  _EVAL_1737;
  wire  _EVAL_1742;
  wire  _EVAL_1744;
  wire  _EVAL_1746;
  wire  _EVAL_1747;
  wire  _EVAL_1748;
  wire  _EVAL_1753;
  wire  _EVAL_1756;
  wire  _EVAL_1759;
  wire  _EVAL_1760;
  wire  _EVAL_1766;
  wire  _EVAL_1767;
  wire  _EVAL_1770;
  wire  _EVAL_1772;
  wire  _EVAL_1775;
  wire  _EVAL_1776;
  reg [126:0] _EVAL_1777;
  wire  _EVAL_1778;
  wire  _EVAL_1782;
  wire  _EVAL_1784;
  wire  _EVAL_1786;
  wire  _EVAL_1790;
  wire  _EVAL_1791;
  wire  _EVAL_1795;
  wire  _EVAL_1798;
  wire  _EVAL_1800;
  wire  _EVAL_1803;
  wire  _EVAL_1804;
  wire  _EVAL_1806;
  wire  _EVAL_1807;
  wire  _EVAL_1808;
  wire  _EVAL_1810;
  wire  _EVAL_1811;
  wire  _EVAL_1814;
  wire  _EVAL_1816;
  wire  _EVAL_1817;
  wire  _EVAL_1818;
  wire  _EVAL_1819;
  wire  _EVAL_1820;
  wire  _EVAL_1823;
  wire  _EVAL_1825;
  wire  _EVAL_1827;
  wire  _EVAL_1829;
  wire  _EVAL_1831;
  wire  _EVAL_1834;
  wire  _EVAL_1835;
  wire  _EVAL_1836;
  wire  _EVAL_1837;
  wire  _EVAL_1838;
  wire  _EVAL_1839;
  wire  _EVAL_1840;
  wire  _EVAL_1841;
  wire  _EVAL_1842;
  wire  _EVAL_1844;
  wire  _EVAL_1845;
  wire  _EVAL_1846;
  wire  _EVAL_1848;
  wire  _EVAL_1849;
  wire  _EVAL_1850;
  wire  _EVAL_1851;
  wire  _EVAL_1856;
  wire  _EVAL_1858;
  wire  _EVAL_1859;
  wire  _EVAL_1860;
  wire  _EVAL_1861;
  wire  _EVAL_1862;
  wire  _EVAL_1863;
  wire  _EVAL_1864;
  wire  _EVAL_1865;
  wire  _EVAL_1868;
  wire  _EVAL_1870;
  wire  _EVAL_1873;
  wire  _EVAL_1874;
  wire  _EVAL_1878;
  wire  _EVAL_1881;
  wire  _EVAL_1883;
  wire  _EVAL_1885;
  wire  _EVAL_1887;
  wire  _EVAL_1888;
  wire  _EVAL_1889;
  wire  _EVAL_1891;
  wire  _EVAL_1893;
  wire  _EVAL_1894;
  wire  _EVAL_1895;
  wire  _EVAL_1897;
  wire  _EVAL_1898;
  wire  _EVAL_1906;
  wire  _EVAL_1908;
  wire  _EVAL_1909;
  wire  _EVAL_1910;
  wire  _EVAL_1911;
  wire  _EVAL_1913;
  wire  _EVAL_1914;
  wire  _EVAL_1915;
  wire  _EVAL_1916;
  wire  _EVAL_1917;
  wire  _EVAL_1919;
  wire  _EVAL_1921;
  wire  _EVAL_1922;
  wire  _EVAL_1924;
  wire  _EVAL_1926;
  wire  _EVAL_1927;
  wire  _EVAL_1929;
  wire  _EVAL_1930;
  wire  _EVAL_1931;
  wire  _EVAL_1933;
  wire  _EVAL_1934;
  wire  _EVAL_1938;
  wire  _EVAL_1939;
  wire  _EVAL_1940;
  wire  _EVAL_1941;
  wire  _EVAL_1943;
  wire  _EVAL_1945;
  wire  _EVAL_1950;
  wire  _EVAL_1951;
  wire  _EVAL_1955;
  wire  _EVAL_1958;
  wire  _EVAL_1959;
  wire  _EVAL_1961;
  wire  _EVAL_1965;
  wire  _EVAL_1967;
  wire  _EVAL_1970;
  wire  _EVAL_1971;
  wire  _EVAL_1974;
  wire  _EVAL_1975;
  wire  _EVAL_1977;
  wire  _EVAL_1979;
  wire  _EVAL_1980;
  wire  _EVAL_1981;
  wire  _EVAL_1983;
  wire  _EVAL_1984;
  wire  _EVAL_1986;
  wire  _EVAL_1989;
  wire  _EVAL_1991;
  wire  _EVAL_1992;
  wire  _EVAL_1993;
  wire  _EVAL_1995;
  wire  _EVAL_1996;
  wire  _EVAL_1999;
  wire  _EVAL_2000;
  wire  _EVAL_2001;
  wire  _EVAL_2002;
  wire  _EVAL_2003;
  wire  _EVAL_2006;
  wire  _EVAL_2007;
  wire  _EVAL_2010;
  wire  _EVAL_2013;
  wire  _EVAL_2014;
  wire  _EVAL_2016;
  wire  _EVAL_2022;
  wire  _EVAL_2024;
  wire  _EVAL_2025;
  wire  _EVAL_2026;
  wire  _EVAL_2029;
  wire  _EVAL_2031;
  wire  _EVAL_2032;
  wire  _EVAL_2033;
  wire  _EVAL_2036;
  wire  _EVAL_2037;
  wire [1023:0] _EVAL_2038;
  wire  _EVAL_2039;
  wire  _EVAL_2040;
  wire  _EVAL_2041;
  wire  _EVAL_2042;
  wire  _EVAL_2044;
  wire  _EVAL_2045;
  wire  _EVAL_2046;
  wire  _EVAL_2047;
  wire  _EVAL_2048;
  wire  _EVAL_2050;
  wire  _EVAL_2052;
  wire  _EVAL_2056;
  wire  _EVAL_2058;
  wire  _EVAL_2063;
  wire  _EVAL_2065;
  wire  _EVAL_2066;
  wire  _EVAL_2067;
  wire  _EVAL_2068;
  wire  _EVAL_2071;
  wire  _EVAL_2072;
  wire  _EVAL_2073;
  wire  _EVAL_2076;
  wire  _EVAL_2082;
  wire  _EVAL_2085;
  wire  _EVAL_2086;
  wire  _EVAL_2089;
  wire  _EVAL_2092;
  wire  _EVAL_2093;
  wire  _EVAL_2096;
  wire  _EVAL_2100;
  wire  _EVAL_2101;
  wire  _EVAL_2104;
  wire  _EVAL_2105;
  wire  _EVAL_2107;
  wire  _EVAL_2108;
  wire  _EVAL_2110;
  wire  _EVAL_2111;
  wire  _EVAL_2112;
  wire [6:0] _EVAL_2115;
  wire  _EVAL_2116;
  wire  _EVAL_2117;
  wire  _EVAL_2118;
  wire  _EVAL_2120;
  wire  _EVAL_2125;
  wire  _EVAL_2126;
  wire  _EVAL_2127;
  wire  _EVAL_2128;
  wire  _EVAL_2135;
  wire  _EVAL_2136;
  wire  _EVAL_2137;
  wire  _EVAL_2138;
  wire  _EVAL_2139;
  wire  _EVAL_2141;
  wire  _EVAL_2146;
  wire  _EVAL_2151;
  wire  _EVAL_2154;
  wire  _EVAL_2156;
  wire  _EVAL_2157;
  wire  _EVAL_2158;
  wire  _EVAL_2161;
  wire  _EVAL_2162;
  wire  _EVAL_2163;
  wire  _EVAL_2164;
  wire  _EVAL_2166;
  wire  _EVAL_2169;
  wire  _EVAL_2170;
  wire  _EVAL_2172;
  wire  _EVAL_2173;
  wire  _EVAL_2176;
  wire  _EVAL_2177;
  wire  _EVAL_2180;
  wire  _EVAL_2181;
  wire  _EVAL_2183;
  wire  _EVAL_2184;
  wire  _EVAL_2185;
  wire  _EVAL_2187;
  wire  _EVAL_2188;
  wire  _EVAL_2189;
  wire  _EVAL_2192;
  wire  _EVAL_2194;
  wire  _EVAL_2200;
  wire  _EVAL_2201;
  wire  _EVAL_2203;
  wire  _EVAL_2208;
  wire  _EVAL_2209;
  wire  _EVAL_2210;
  wire  _EVAL_2212;
  wire  _EVAL_2213;
  wire  _EVAL_2214;
  wire  _EVAL_2215;
  wire  _EVAL_2219;
  wire  _EVAL_2223;
  wire  _EVAL_2225;
  wire  _EVAL_2228;
  wire  _EVAL_2229;
  wire  _EVAL_2232;
  wire  _EVAL_2235;
  wire  _EVAL_2237;
  wire  _EVAL_2238;
  wire  _EVAL_2239;
  wire  _EVAL_2240;
  wire  _EVAL_2241;
  wire  _EVAL_2242;
  wire  _EVAL_2243;
  wire  _EVAL_2244;
  wire  _EVAL_2245;
  wire  _EVAL_2246;
  wire  _EVAL_2247;
  wire  _EVAL_2250;
  wire  _EVAL_2255;
  wire  _EVAL_2256;
  wire  _EVAL_2259;
  wire  _EVAL_2260;
  wire  _EVAL_2261;
  wire  _EVAL_2265;
  wire  _EVAL_2266;
  wire  _EVAL_2267;
  wire  _EVAL_2269;
  wire  _EVAL_2271;
  wire  _EVAL_2272;
  wire  _EVAL_2273;
  wire  _EVAL_2277;
  wire  _EVAL_2278;
  wire  _EVAL_2280;
  wire  _EVAL_2283;
  wire  _EVAL_2286;
  wire  _EVAL_2287;
  wire  _EVAL_2288;
  wire  _EVAL_2290;
  wire  _EVAL_2291;
  wire  _EVAL_2292;
  wire  _EVAL_2295;
  wire  _EVAL_2299;
  wire  _EVAL_2301;
  wire  _EVAL_2302;
  wire  _EVAL_2304;
  wire  _EVAL_2305;
  wire  _EVAL_2307;
  wire  _EVAL_2310;
  wire  _EVAL_2317;
  wire  _EVAL_2319;
  wire  _EVAL_2323;
  wire  _EVAL_2324;
  wire  _EVAL_2325;
  wire  _EVAL_2326;
  wire  _EVAL_2330;
  wire  _EVAL_2331;
  wire  _EVAL_2332;
  wire  _EVAL_2333;
  wire  _EVAL_2334;
  wire  _EVAL_2335;
  wire  _EVAL_2336;
  wire  _EVAL_2338;
  wire  _EVAL_2339;
  wire  _EVAL_2340;
  wire  _EVAL_2343;
  wire  _EVAL_2351;
  wire  _EVAL_2353;
  wire  _EVAL_2355;
  wire  _EVAL_2356;
  wire  _EVAL_2357;
  wire  _EVAL_2358;
  wire  _EVAL_2359;
  wire  _EVAL_2360;
  wire  _EVAL_2363;
  wire  _EVAL_2364;
  wire  _EVAL_2365;
  wire  _EVAL_2367;
  wire  _EVAL_2368;
  wire  _EVAL_2371;
  wire  _EVAL_2372;
  wire  _EVAL_2373;
  wire  _EVAL_2374;
  wire  _EVAL_2376;
  wire  _EVAL_2382;
  wire  _EVAL_2383;
  wire  _EVAL_2387;
  wire  _EVAL_2388;
  wire  _EVAL_2390;
  wire  _EVAL_2393;
  wire  _EVAL_2394;
  wire  _EVAL_2395;
  wire  _EVAL_2398;
  wire  _EVAL_2400;
  wire  _EVAL_2401;
  wire  _EVAL_2402;
  wire  _EVAL_2404;
  wire  _EVAL_2405;
  wire  _EVAL_2407;
  wire  _EVAL_2409;
  wire  _EVAL_2411;
  wire  _EVAL_2412;
  wire  _EVAL_2413;
  wire  _EVAL_2414;
  wire  _EVAL_2419;
  wire  _EVAL_2420;
  wire  _EVAL_2421;
  wire  _EVAL_2422;
  wire  _EVAL_2423;
  wire  _EVAL_2426;
  wire  _EVAL_2429;
  wire  _EVAL_2430;
  wire  _EVAL_2432;
  wire  _EVAL_2433;
  wire  _EVAL_2434;
  wire  _EVAL_2435;
  wire  _EVAL_2436;
  wire  _EVAL_2437;
  wire  _EVAL_2442;
  wire  _EVAL_2443;
  wire  _EVAL_2445;
  wire  _EVAL_2446;
  wire  _EVAL_2447;
  wire  _EVAL_2448;
  wire  _EVAL_2449;
  wire  _EVAL_2452;
  wire  _EVAL_2456;
  wire  _EVAL_2457;
  wire  _EVAL_2458;
  wire  _EVAL_2459;
  wire  _EVAL_2461;
  wire  _EVAL_2463;
  wire  _EVAL_2464;
  wire  _EVAL_2467;
  wire  _EVAL_2468;
  wire  _EVAL_2470;
  wire  _EVAL_2471;
  wire  _EVAL_2475;
  wire  _EVAL_2480;
  wire  _EVAL_2481;
  wire  _EVAL_2485;
  wire  _EVAL_2487;
  wire  _EVAL_2489;
  wire  _EVAL_2491;
  wire  _EVAL_2493;
  wire  _EVAL_2496;
  wire  _EVAL_2497;
  wire  _EVAL_2500;
  wire  _EVAL_2501;
  wire  _EVAL_2504;
  wire  _EVAL_2505;
  wire  _EVAL_2506;
  wire  _EVAL_2507;
  wire  _EVAL_2508;
  wire  _EVAL_2510;
  wire  _EVAL_2512;
  wire  _EVAL_2513;
  wire  _EVAL_2514;
  wire  _EVAL_2516;
  wire  _EVAL_2519;
  wire  _EVAL_2522;
  wire  _EVAL_2524;
  wire  _EVAL_2526;
  wire  _EVAL_2528;
  wire  _EVAL_2529;
  wire  _EVAL_2532;
  wire  _EVAL_2535;
  wire  _EVAL_2536;
  wire  _EVAL_2538;
  wire  _EVAL_2539;
  wire  _EVAL_2540;
  wire  _EVAL_2541;
  wire  _EVAL_2543;
  wire  _EVAL_2544;
  wire  _EVAL_2545;
  wire  _EVAL_2546;
  wire  _EVAL_2547;
  wire  _EVAL_2548;
  wire  _EVAL_2550;
  wire  _EVAL_2551;
  wire  _EVAL_2552;
  wire  _EVAL_2553;
  wire  _EVAL_2560;
  wire  _EVAL_2562;
  wire  _EVAL_2563;
  wire  _EVAL_2564;
  wire  _EVAL_2566;
  wire  _EVAL_2567;
  wire  _EVAL_2569;
  wire  _EVAL_2570;
  wire  _EVAL_2573;
  wire  _EVAL_2574;
  wire  _EVAL_2578;
  wire  _EVAL_2579;
  wire  _EVAL_2581;
  wire  _EVAL_2582;
  wire  _EVAL_2583;
  wire  _EVAL_2584;
  wire  _EVAL_2585;
  wire  _EVAL_2587;
  wire  _EVAL_2588;
  wire  _EVAL_2590;
  wire  _EVAL_2591;
  wire  _EVAL_2592;
  wire  _EVAL_2594;
  wire  _EVAL_2595;
  wire  _EVAL_2596;
  wire  _EVAL_2597;
  wire  _EVAL_2598;
  wire  _EVAL_2599;
  wire  _EVAL_2600;
  wire  _EVAL_2602;
  wire  _EVAL_2603;
  wire  _EVAL_2605;
  wire  _EVAL_2606;
  wire  _EVAL_2608;
  wire  _EVAL_2609;
  wire [126:0] _EVAL_2610;
  wire  _EVAL_2611;
  wire  _EVAL_2613;
  wire  _EVAL_2620;
  wire  _EVAL_2625;
  wire  _EVAL_2630;
  wire  _EVAL_2631;
  wire  _EVAL_2634;
  wire  _EVAL_2635;
  wire  _EVAL_2636;
  wire  _EVAL_2638;
  wire  _EVAL_2640;
  wire  _EVAL_2641;
  wire  _EVAL_2642;
  wire  _EVAL_2643;
  wire  _EVAL_2644;
  wire  _EVAL_2645;
  wire  _EVAL_2646;
  wire  _EVAL_2647;
  wire  _EVAL_2648;
  wire  _EVAL_2652;
  wire  _EVAL_2656;
  wire  _EVAL_2657;
  wire  _EVAL_2662;
  wire  _EVAL_2664;
  wire  _EVAL_2665;
  wire  _EVAL_2666;
  wire  _EVAL_2669;
  wire  _EVAL_2670;
  wire  _EVAL_2673;
  wire  _EVAL_2674;
  wire  _EVAL_2675;
  wire  _EVAL_2677;
  wire  _EVAL_2678;
  wire  _EVAL_2679;
  wire  _EVAL_2680;
  wire  _EVAL_2681;
  wire  _EVAL_2683;
  wire  _EVAL_2684;
  wire  _EVAL_2687;
  wire  _EVAL_2688;
  wire  _EVAL_2690;
  wire  _EVAL_2691;
  wire  _EVAL_2695;
  wire [1:0] _EVAL_2699;
  wire  _EVAL_2703;
  wire  _EVAL_2704;
  wire  _EVAL_2706;
  wire  _EVAL_2707;
  wire  _EVAL_2708;
  wire  _EVAL_2709;
  wire  _EVAL_2713;
  wire  _EVAL_2714;
  wire  _EVAL_2718;
  wire  _EVAL_2721;
  wire  _EVAL_2723;
  wire  _EVAL_2725;
  wire  _EVAL_2726;
  wire  _EVAL_2729;
  wire  _EVAL_2731;
  wire  _EVAL_2735;
  wire  _EVAL_2736;
  wire  _EVAL_2740;
  wire  _EVAL_2741;
  wire  _EVAL_2743;
  wire  _EVAL_2744;
  wire  _EVAL_2746;
  wire [3:0] _EVAL_2748;
  wire  _EVAL_2749;
  wire  _EVAL_2750;
  wire  _EVAL_2751;
  wire  _EVAL_2752;
  wire  _EVAL_2754;
  wire  _EVAL_2755;
  wire  _EVAL_2760;
  wire  _EVAL_2761;
  wire  _EVAL_2762;
  wire  _EVAL_2764;
  wire  _EVAL_2766;
  wire  _EVAL_2768;
  wire  _EVAL_2769;
  wire  _EVAL_2771;
  wire [19:0] _EVAL_2775;
  wire  _EVAL_2776;
  wire  _EVAL_2778;
  wire  _EVAL_2780;
  wire  _EVAL_2783;
  wire  _EVAL_2785;
  wire  _EVAL_2786;
  wire  _EVAL_2790;
  wire  _EVAL_2792;
  wire  _EVAL_2794;
  wire  _EVAL_2796;
  wire  _EVAL_2797;
  wire  _EVAL_2802;
  wire  _EVAL_2804;
  wire  _EVAL_2806;
  wire  _EVAL_2807;
  wire  _EVAL_2808;
  wire  _EVAL_2809;
  wire  _EVAL_2813;
  wire  _EVAL_2815;
  wire  _EVAL_2816;
  wire  _EVAL_2818;
  wire  _EVAL_2819;
  wire  _EVAL_2820;
  wire  _EVAL_2821;
  wire  _EVAL_2823;
  wire  _EVAL_2824;
  wire  _EVAL_2825;
  wire  _EVAL_2826;
  wire  _EVAL_2827;
  wire  _EVAL_2829;
  wire  _EVAL_2830;
  wire  _EVAL_2831;
  wire  _EVAL_2834;
  wire  _EVAL_2835;
  wire  _EVAL_2836;
  wire  _EVAL_2837;
  wire  _EVAL_2839;
  wire  _EVAL_2840;
  wire  _EVAL_2843;
  wire  _EVAL_2847;
  wire  _EVAL_2848;
  wire  _EVAL_2851;
  wire  _EVAL_2854;
  wire  _EVAL_2857;
  wire  _EVAL_2858;
  wire  _EVAL_2859;
  wire  _EVAL_2864;
  wire  _EVAL_2866;
  wire  _EVAL_2867;
  wire  _EVAL_2869;
  wire  _EVAL_2870;
  wire  _EVAL_2875;
  wire  _EVAL_2876;
  wire  _EVAL_2882;
  wire  _EVAL_2883;
  wire  _EVAL_2884;
  wire  _EVAL_2886;
  wire  _EVAL_2887;
  reg  _EVAL_2890;
  wire  _EVAL_2891;
  wire  _EVAL_2893;
  wire  _EVAL_2894;
  wire  _EVAL_2895;
  wire  _EVAL_2897;
  wire  _EVAL_2898;
  wire  _EVAL_2899;
  wire  _EVAL_2901;
  wire  _EVAL_2905;
  wire  _EVAL_2908;
  wire  _EVAL_2909;
  wire  _EVAL_2912;
  wire  _EVAL_2916;
  wire  _EVAL_2920;
  wire  _EVAL_2923;
  wire  _EVAL_2924;
  wire  _EVAL_2925;
  wire  _EVAL_2930;
  wire  _EVAL_2931;
  wire  _EVAL_2933;
  wire  _EVAL_2937;
  wire  _EVAL_2939;
  wire  _EVAL_2940;
  wire  _EVAL_2941;
  wire  _EVAL_2943;
  wire  _EVAL_2947;
  wire  _EVAL_2948;
  wire  _EVAL_2949;
  wire  _EVAL_2950;
  wire  _EVAL_2953;
  wire  _EVAL_2954;
  wire  _EVAL_2955;
  wire  _EVAL_2958;
  wire  _EVAL_2959;
  wire  _EVAL_2960;
  wire  _EVAL_2962;
  wire  _EVAL_2964;
  wire  _EVAL_2967;
  wire  _EVAL_2971;
  wire  _EVAL_2972;
  wire  _EVAL_2973;
  wire  _EVAL_2976;
  wire  _EVAL_2984;
  wire  _EVAL_2991;
  wire  _EVAL_2993;
  wire  _EVAL_2994;
  wire  _EVAL_2995;
  wire  _EVAL_3003;
  wire  _EVAL_3004;
  wire  _EVAL_3006;
  wire  _EVAL_3009;
  wire  _EVAL_3010;
  wire  _EVAL_3012;
  wire  _EVAL_3016;
  wire  _EVAL_3018;
  wire  _EVAL_3019;
  wire  _EVAL_3020;
  wire  _EVAL_3021;
  wire  _EVAL_3022;
  wire  _EVAL_3023;
  wire  _EVAL_3024;
  wire  _EVAL_3025;
  wire  _EVAL_3026;
  wire  _EVAL_3028;
  wire  _EVAL_3031;
  wire  _EVAL_3032;
  wire  _EVAL_3041;
  wire  _EVAL_3042;
  wire  _EVAL_3044;
  wire  _EVAL_3045;
  wire  _EVAL_3046;
  wire  _EVAL_3048;
  wire  _EVAL_3049;
  wire  _EVAL_3050;
  wire  _EVAL_3051;
  wire  _EVAL_3052;
  wire  _EVAL_3053;
  wire  _EVAL_3054;
  wire  _EVAL_3057;
  wire  _EVAL_3058;
  wire  _EVAL_3060;
  wire  _EVAL_3062;
  wire  _EVAL_3065;
  wire  _EVAL_3066;
  wire  _EVAL_3070;
  wire  _EVAL_3073;
  wire  _EVAL_3078;
  wire  _EVAL_3079;
  wire  _EVAL_3083;
  wire  _EVAL_3085;
  wire  _EVAL_3087;
  wire  _EVAL_3088;
  wire  _EVAL_3090;
  wire  _EVAL_3091;
  wire  _EVAL_3092;
  wire [127:0] _EVAL_3093;
  wire  _EVAL_3098;
  wire  _EVAL_3103;
  wire  _EVAL_3109;
  wire  _EVAL_3110;
  wire  _EVAL_3113;
  wire  _EVAL_3116;
  wire  _EVAL_3117;
  wire  _EVAL_3118;
  wire  _EVAL_3119;
  wire  _EVAL_3120;
  wire  _EVAL_3121;
  wire  _EVAL_3125;
  wire  _EVAL_3126;
  wire  _EVAL_3128;
  wire  _EVAL_3131;
  wire  _EVAL_3132;
  wire  _EVAL_3135;
  wire  _EVAL_3136;
  wire  _EVAL_3137;
  wire  _EVAL_3139;
  wire  _EVAL_3141;
  wire  _EVAL_3143;
  wire  _EVAL_3144;
  wire  _EVAL_3146;
  wire  _EVAL_3149;
  wire  _EVAL_3154;
  wire  _EVAL_3158;
  wire  _EVAL_3159;
  wire  _EVAL_3160;
  wire  _EVAL_3163;
  wire  _EVAL_3164;
  wire  _EVAL_3168;
  wire [6:0] _EVAL_3169;
  wire  _EVAL_3170;
  wire  _EVAL_3173;
  wire  _EVAL_3175;
  wire  _EVAL_3176;
  wire  _EVAL_3178;
  wire  _EVAL_3180;
  wire  _EVAL_3181;
  wire  _EVAL_3184;
  wire [28:0] _EVAL_3187;
  wire  _EVAL_3188;
  wire  _EVAL_3190;
  wire  _EVAL_3192;
  wire  _EVAL_3194;
  wire  _EVAL_3195;
  wire  _EVAL_3196;
  wire  _EVAL_3197;
  wire  _EVAL_3203;
  wire  _EVAL_3207;
  wire  _EVAL_3208;
  wire  _EVAL_3212;
  wire  _EVAL_3215;
  wire  _EVAL_3224;
  wire  _EVAL_3226;
  wire  _EVAL_3227;
  wire  _EVAL_3228;
  wire  _EVAL_3229;
  wire  _EVAL_3230;
  wire  _EVAL_3231;
  wire  _EVAL_3232;
  wire  _EVAL_3233;
  wire  _EVAL_3234;
  wire  _EVAL_3235;
  wire  _EVAL_3238;
  wire  _EVAL_3239;
  wire  _EVAL_3247;
  wire  _EVAL_3248;
  wire  _EVAL_3250;
  wire  _EVAL_3252;
  wire  _EVAL_3253;
  wire  _EVAL_3254;
  wire  _EVAL_3257;
  wire  _EVAL_3258;
  wire  _EVAL_3269;
  wire  _EVAL_3272;
  wire  _EVAL_3273;
  wire  _EVAL_3274;
  wire  _EVAL_3277;
  wire  _EVAL_3279;
  wire  _EVAL_3280;
  wire  _EVAL_3281;
  wire  _EVAL_3282;
  wire  _EVAL_3283;
  wire  _EVAL_3289;
  wire  _EVAL_3292;
  wire  _EVAL_3293;
  wire  _EVAL_3294;
  wire  _EVAL_3295;
  wire  _EVAL_3296;
  wire  _EVAL_3297;
  wire  _EVAL_3298;
  wire  _EVAL_3300;
  wire  _EVAL_3301;
  wire  _EVAL_3306;
  wire  _EVAL_3308;
  wire  _EVAL_3309;
  wire  _EVAL_3310;
  wire [28:0] _EVAL_3313;
  wire  _EVAL_3314;
  wire  _EVAL_3320;
  wire  _EVAL_3323;
  wire  _EVAL_3325;
  wire  _EVAL_3332;
  wire  _EVAL_3333;
  wire  _EVAL_3334;
  wire  _EVAL_3338;
  wire  _EVAL_3344;
  wire  _EVAL_3348;
  wire  _EVAL_3350;
  wire  _EVAL_3351;
  wire  _EVAL_3352;
  wire  _EVAL_3356;
  wire  _EVAL_3360;
  wire  _EVAL_3362;
  wire  _EVAL_3364;
  wire  _EVAL_3365;
  wire  _EVAL_3369;
  wire  _EVAL_3371;
  wire  _EVAL_3372;
  wire  _EVAL_3377;
  wire  _EVAL_3379;
  wire  _EVAL_3380;
  wire  _EVAL_3382;
  wire  _EVAL_3383;
  wire  _EVAL_3385;
  wire  _EVAL_3389;
  wire  _EVAL_3396;
  wire  _EVAL_3398;
  wire  _EVAL_3400;
  wire [2:0] _EVAL_3403;
  wire  _EVAL_3405;
  wire  _EVAL_3406;
  wire  _EVAL_3407;
  wire  _EVAL_3411;
  wire  _EVAL_3413;
  wire  _EVAL_3415;
  wire  _EVAL_3419;
  wire  _EVAL_3421;
  wire  _EVAL_3423;
  wire  _EVAL_3424;
  wire  _EVAL_3428;
  wire [9:0] _EVAL_3429;
  wire  _EVAL_3432;
  wire  _EVAL_3439;
  wire  _EVAL_3441;
  wire  _EVAL_3445;
  wire  _EVAL_3447;
  wire  _EVAL_3448;
  wire  _EVAL_3451;
  wire  _EVAL_3452;
  wire  _EVAL_3453;
  wire  _EVAL_3458;
  wire  _EVAL_3459;
  wire  _EVAL_3464;
  wire  _EVAL_3466;
  wire  _EVAL_3470;
  wire  _EVAL_3472;
  wire  _EVAL_3473;
  wire  _EVAL_3477;
  wire  _EVAL_3478;
  wire  _EVAL_3482;
  wire  _EVAL_3484;
  wire  _EVAL_3487;
  wire  _EVAL_3491;
  wire  _EVAL_3492;
  wire  _EVAL_3493;
  wire  _EVAL_3495;
  wire  _EVAL_3496;
  wire  _EVAL_3497;
  wire  _EVAL_3498;
  wire [7:0] _EVAL_3499;
  wire  _EVAL_3500;
  wire  _EVAL_3501;
  wire  _EVAL_3502;
  wire  _EVAL_3503;
  wire  _EVAL_3506;
  wire  _EVAL_3507;
  wire  _EVAL_3509;
  wire  _EVAL_3511;
  wire  _EVAL_3512;
  wire  _EVAL_3514;
  wire  _EVAL_3515;
  wire  _EVAL_3517;
  wire  _EVAL_3518;
  wire  _EVAL_3522;
  wire  _EVAL_3525;
  wire  _EVAL_3532;
  wire  _EVAL_3535;
  wire  _EVAL_3536;
  wire  _EVAL_3539;
  wire  _EVAL_3540;
  wire  _EVAL_3541;
  wire  _EVAL_3542;
  wire  _EVAL_3543;
  wire  _EVAL_3544;
  wire  _EVAL_3546;
  wire  _EVAL_3547;
  wire  _EVAL_3549;
  wire  _EVAL_3550;
  wire  _EVAL_3551;
  wire  _EVAL_3552;
  wire  _EVAL_3553;
  wire  _EVAL_3554;
  wire  _EVAL_3556;
  wire  _EVAL_3558;
  wire  _EVAL_3561;
  wire  _EVAL_3562;
  wire  _EVAL_3563;
  wire  _EVAL_3565;
  wire  _EVAL_3570;
  wire  _EVAL_3573;
  wire  _EVAL_3574;
  wire  _EVAL_3578;
  wire  _EVAL_3580;
  wire  _EVAL_3581;
  wire  _EVAL_3582;
  wire  _EVAL_3583;
  wire  _EVAL_3584;
  wire  _EVAL_3585;
  wire  _EVAL_3586;
  wire  _EVAL_3592;
  wire  _EVAL_3594;
  wire  _EVAL_3598;
  wire  _EVAL_3601;
  wire  _EVAL_3602;
  wire  _EVAL_3604;
  wire  _EVAL_3605;
  wire  _EVAL_3606;
  wire  _EVAL_3607;
  wire  _EVAL_3608;
  wire  _EVAL_3609;
  wire  _EVAL_3611;
  wire  _EVAL_3614;
  wire  _EVAL_3617;
  wire  _EVAL_3621;
  wire  _EVAL_3623;
  wire  _EVAL_3625;
  wire  _EVAL_3628;
  wire  _EVAL_3629;
  wire  _EVAL_3630;
  wire  _EVAL_3631;
  wire  _EVAL_3634;
  wire  _EVAL_3640;
  wire  _EVAL_3641;
  wire  _EVAL_3645;
  wire  _EVAL_3647;
  wire  _EVAL_3648;
  wire  _EVAL_3649;
  wire  _EVAL_3650;
  wire  _EVAL_3655;
  wire  _EVAL_3658;
  wire  _EVAL_3659;
  wire  _EVAL_3660;
  wire  _EVAL_3661;
  wire  _EVAL_3664;
  wire  _EVAL_3665;
  wire  _EVAL_3666;
  wire  _EVAL_3668;
  wire  _EVAL_3669;
  wire  _EVAL_3670;
  wire  _EVAL_3671;
  wire  _EVAL_3673;
  wire  _EVAL_3674;
  wire  _EVAL_3675;
  wire  _EVAL_3676;
  wire  _EVAL_3677;
  wire  _EVAL_3678;
  wire  _EVAL_3679;
  wire  _EVAL_3682;
  wire  _EVAL_3687;
  wire  _EVAL_3688;
  wire  _EVAL_3689;
  wire  _EVAL_3690;
  wire  _EVAL_3691;
  wire  _EVAL_3693;
  wire  _EVAL_3694;
  wire  _EVAL_3697;
  wire  _EVAL_3698;
  wire  _EVAL_3699;
  wire  _EVAL_3703;
  wire  _EVAL_3705;
  wire  _EVAL_3707;
  wire  _EVAL_3709;
  wire  _EVAL_3710;
  wire  _EVAL_3712;
  wire  _EVAL_3713;
  wire  _EVAL_3721;
  wire  _EVAL_3724;
  wire  _EVAL_3727;
  wire  _EVAL_3728;
  wire  _EVAL_3730;
  wire  _EVAL_3731;
  wire  _EVAL_3733;
  wire  _EVAL_3736;
  wire  _EVAL_3738;
  wire  _EVAL_3739;
  wire  _EVAL_3740;
  wire  _EVAL_3741;
  wire  _EVAL_3748;
  wire  _EVAL_3749;
  wire  _EVAL_3750;
  wire  _EVAL_3752;
  wire  _EVAL_3753;
  wire  _EVAL_3754;
  wire  _EVAL_3755;
  wire  _EVAL_3758;
  wire  _EVAL_3761;
  wire  _EVAL_3763;
  wire  _EVAL_3764;
  wire  _EVAL_3765;
  wire  _EVAL_3766;
  wire  _EVAL_3767;
  wire  _EVAL_3768;
  wire  _EVAL_3769;
  wire  _EVAL_3771;
  wire  _EVAL_3773;
  wire  _EVAL_3774;
  wire [1:0] _EVAL_3776;
  wire  _EVAL_3778;
  wire  _EVAL_3779;
  wire [7:0] _EVAL_3780;
  wire  _EVAL_3781;
  wire  _EVAL_3783;
  wire  _EVAL_3784;
  wire  _EVAL_3785;
  wire  _EVAL_3788;
  wire  _EVAL_3789;
  wire  _EVAL_3790;
  wire  _EVAL_3792;
  wire  _EVAL_3795;
  wire  _EVAL_3796;
  wire  _EVAL_3799;
  wire [7:0] _EVAL_3805;
  wire  _EVAL_3808;
  wire  _EVAL_3810;
  wire  _EVAL_3812;
  wire  _EVAL_3813;
  wire  _EVAL_3814;
  wire  _EVAL_3816;
  wire  _EVAL_3817;
  wire  _EVAL_3818;
  wire  _EVAL_3820;
  wire  _EVAL_3821;
  wire  _EVAL_3822;
  wire  _EVAL_3823;
  wire  _EVAL_3826;
  wire  _EVAL_3827;
  wire  _EVAL_3829;
  wire  _EVAL_3830;
  wire  _EVAL_3833;
  wire  _EVAL_3836;
  wire  _EVAL_3837;
  wire  _EVAL_3838;
  wire  _EVAL_3839;
  wire  _EVAL_3841;
  wire  _EVAL_3843;
  wire  _EVAL_3846;
  wire  _EVAL_3853;
  wire  _EVAL_3854;
  _EVAL_95_assert monitor (
    ._EVAL(monitor__EVAL),
    ._EVAL_0(monitor__EVAL_0),
    ._EVAL_1(monitor__EVAL_1),
    ._EVAL_2(monitor__EVAL_2),
    ._EVAL_3(monitor__EVAL_3),
    ._EVAL_4(monitor__EVAL_4),
    ._EVAL_5(monitor__EVAL_5),
    ._EVAL_6(monitor__EVAL_6),
    ._EVAL_7(monitor__EVAL_7),
    ._EVAL_8(monitor__EVAL_8),
    ._EVAL_9(monitor__EVAL_9),
    ._EVAL_10(monitor__EVAL_10),
    ._EVAL_11(monitor__EVAL_11),
    ._EVAL_12(monitor__EVAL_12),
    ._EVAL_13(monitor__EVAL_13),
    ._EVAL_14(monitor__EVAL_14)
  );
  assign _EVAL_1814 = _EVAL_2532 & _EVAL_2764;
  assign _EVAL_477 = _EVAL_623 & _EVAL_2047;
  assign _EVAL_3752 = _EVAL_2356 & _EVAL_3830;
  assign _EVAL_551 = _EVAL_3774 & _EVAL_2540;
  assign _EVAL_1229 = _EVAL_1649 & _EVAL_3133;
  assign _EVAL_3606 = |_EVAL_1272;
  assign _EVAL_1859 = _EVAL_1424 & _EVAL_2047;
  assign _EVAL_1107 = _EVAL_173 & _EVAL_405;
  assign _EVAL_1562 = _EVAL_1927 & _EVAL_2273;
  assign _EVAL_2519 = _EVAL_2991 & _EVAL_2047;
  assign _EVAL_729 = _EVAL_1927 & _EVAL_3792;
  assign _EVAL_1888 = _EVAL_1649 & _EVAL_2395;
  assign _EVAL_867 = _EVAL_2584 & _EVAL_1004;
  assign _EVAL_3296 = _EVAL_920 & _EVAL_802;
  assign _EVAL_2513 = _EVAL_702 & _EVAL_701;
  assign _EVAL_3020 = _EVAL_1361[9];
  assign _EVAL_2166 = _EVAL_1361[17];
  assign _EVAL_2755 = _EVAL_3604 & _EVAL_2047;
  assign _EVAL_2448 = _EVAL_2532 & _EVAL_3060;
  assign _EVAL_1979 = _EVAL_895 & _EVAL_2047;
  assign _EVAL_1289 = _EVAL_2948 & _EVAL_2047;
  assign _EVAL_345 = _EVAL_2850[16];
  assign _EVAL_237 = _EVAL_1649 & _EVAL_2152;
  assign _EVAL_2642 = _EVAL_2993 & _EVAL_2096;
  assign _EVAL_3385 = _EVAL_1927 & _EVAL_1378;
  assign _EVAL_1893 = _EVAL_2532 & _EVAL_1685;
  assign _EVAL_622 = _EVAL_3749 & _EVAL_3827;
  assign _EVAL_1234 = _EVAL_3585 & _EVAL_914;
  assign _EVAL_803 = _EVAL_1776 & _EVAL_2941;
  assign _EVAL_1206 = _EVAL_376 & _EVAL_701;
  assign _EVAL_2305 = _EVAL_3546 & _EVAL_701;
  assign _EVAL_395 = _EVAL_3573 & _EVAL_1004;
  assign _EVAL_431 = _EVAL_2993 & _EVAL_1730;
  assign _EVAL_2536 = _EVAL_173 & _EVAL_3498;
  assign _EVAL_887 = _EVAL_3125 & _EVAL_1245;
  assign _EVAL_1125 = |_EVAL_1839;
  assign _EVAL_2022 = _EVAL_2993 & _EVAL_2540;
  assign _EVAL_399 = _EVAL_2038[259];
  assign _EVAL_3103 = _EVAL_1927 & _EVAL_2834;
  assign _EVAL_974 = _EVAL_2038[23];
  assign _EVAL_2214 = _EVAL_2038[58];
  assign _EVAL_3141 = _EVAL_2746 & _EVAL_701;
  assign _EVAL_3400 = _EVAL_2532 & _EVAL_3405;
  assign _EVAL_1603 = _EVAL_3383 & _EVAL_2047;
  assign _EVAL_2830 = _EVAL_1649 & _EVAL_3489;
  assign _EVAL_2442 = _EVAL_1927 & _EVAL_1619;
  assign _EVAL_1611 = _EVAL_1421 & _EVAL_826;
  assign _EVAL_1004 = |_EVAL_3403;
  assign _EVAL_481 = |_EVAL_1070;
  assign _EVAL_900 = _EVAL_2687 & _EVAL_826;
  assign _EVAL_3025 = _EVAL_2203 & _EVAL_2941;
  assign _EVAL_409 = _EVAL_152 & _EVAL_826;
  assign _EVAL_204 = _EVAL_2038[76];
  assign _EVAL_3348 = _EVAL_3585 & _EVAL_3407;
  assign _EVAL_2419 = _EVAL_1649 & _EVAL_3757;
  assign _EVAL_2422 = _EVAL_2038[10];
  assign _EVAL_3671 = _EVAL_2532 & _EVAL_1665;
  assign _EVAL_1841 = _EVAL_3562 & _EVAL_2436;
  assign _EVAL_3607 = _EVAL_1927 & _EVAL_2826;
  assign _EVAL_3143 = _EVAL_1649 & _EVAL_2224;
  assign _EVAL_2487 = |_EVAL_586;
  assign _EVAL_3645 = _EVAL_920 & _EVAL_154;
  assign _EVAL_187 = _EVAL_2038[49];
  assign _EVAL_969 = _EVAL_2038[89];
  assign _EVAL_290 = |_EVAL_1035;
  assign _EVAL_1461 = _EVAL_665 & _EVAL_826;
  assign _EVAL_2112 = _EVAL_1381 & _EVAL_2047;
  assign _EVAL_3535 = _EVAL_1927 & _EVAL_3823;
  assign _EVAL_3184 = _EVAL_2038[106];
  assign _EVAL_2120 = _EVAL_2277 & _EVAL_2047;
  assign _EVAL_701 = &_EVAL_3403;
  assign _EVAL_1497 = _EVAL_2038[128];
  assign _EVAL_1457 = _EVAL_651[129];
  assign _EVAL_3197 = _EVAL_3749 & _EVAL_1811;
  assign _EVAL_2127 = _EVAL_1425 & _EVAL_826;
  assign _EVAL_555 = _EVAL_3503 & _EVAL_826;
  assign _EVAL_1360 = _EVAL_2677 & _EVAL_2047;
  assign _EVAL_2266 = _EVAL_3774 & _EVAL_1442;
  assign _EVAL_2766 = _EVAL_2597 & _EVAL_1004;
  assign _EVAL_3736 = _EVAL_1927 & _EVAL_1950;
  assign _EVAL_3788 = _EVAL_2707 & _EVAL_826;
  assign _EVAL_3674 = _EVAL_1384 & _EVAL_826;
  assign _EVAL_1406 = _EVAL_1649 & _EVAL_2983;
  assign _EVAL_2948 = _EVAL_2532 & _EVAL_2255;
  assign _EVAL_2925 = _EVAL_2014 & _EVAL_701;
  assign _EVAL_2181 = _EVAL_2670 & _EVAL_2047;
  assign _EVAL_211 = _EVAL_2532 & _EVAL_1378;
  assign _EVAL_3423 = |_EVAL_3020;
  assign _EVAL_790 = _EVAL_2038[104];
  assign _EVAL_3158 = _EVAL_2038[99];
  assign _EVAL_1492 = _EVAL_3352 & _EVAL_2047;
  assign _EVAL_1306 = _EVAL_1795 & _EVAL_826;
  assign _EVAL_3238 = _EVAL_1927 & _EVAL_768;
  assign _EVAL_2943 = _EVAL_308 & _EVAL_2047;
  assign _EVAL_3658 = _EVAL_1767 & _EVAL_2941;
  assign _EVAL_1067 = _EVAL_1856 & _EVAL_826;
  assign _EVAL_1558 = _EVAL_2532 & _EVAL_2118;
  assign _EVAL_2407 = _EVAL_2038[62];
  assign _EVAL_1084 = _EVAL_3535 & _EVAL_2047;
  assign _EVAL_1145 = _EVAL_2532 & _EVAL_3698;
  assign _EVAL_587 = _EVAL_1927 & _EVAL_3765;
  assign _EVAL_2215 = _EVAL_2514 & _EVAL_826;
  assign _EVAL_1214 = _EVAL_1927 & _EVAL_3758;
  assign _EVAL_1705 = _EVAL_173 & _EVAL_290;
  assign _EVAL_1458 = _EVAL_2238 & _EVAL_1004;
  assign _EVAL_2695 = _EVAL_1636 & _EVAL_2047;
  assign _EVAL_1469 = _EVAL_3562 & _EVAL_914;
  assign _EVAL_1938 = _EVAL_3126 & _EVAL_1730;
  assign _EVAL_3629 = _EVAL_1064 & _EVAL_1004;
  assign _EVAL_597 = _EVAL_1649 & _EVAL_817;
  assign _EVAL_401 = _EVAL_1927 & _EVAL_1667;
  assign _EVAL_2240 = _EVAL_1927 & _EVAL_3057;
  assign _EVAL_3466 = _EVAL_920 & _EVAL_3605;
  assign _EVAL_3608 = _EVAL_3451 & _EVAL_2941;
  assign _EVAL_983 = _EVAL_1981 & _EVAL_826;
  assign _EVAL_2405 = _EVAL_2532 & _EVAL_188;
  assign _EVAL_2118 = _EVAL_2038[82];
  assign _EVAL_1321 = _EVAL_397 & _EVAL_3764;
  assign _EVAL_2373 = _EVAL_1927 & _EVAL_3308;
  assign _EVAL_2657 = _EVAL_1897 & _EVAL_154;
  assign _EVAL_1313 = _EVAL_543 & _EVAL_826;
  assign _EVAL_3843 = _EVAL_1927 & _EVAL_2422;
  assign _EVAL_1205 = _EVAL_2038[92];
  assign _EVAL_2485 = _EVAL_3109 & _EVAL_826;
  assign _EVAL_2459 = _EVAL_3514 & _EVAL_2047;
  assign _EVAL_1049 = _EVAL_360 & _EVAL_2941;
  assign _EVAL_3707 = _EVAL_2376 & _EVAL_701;
  assign _EVAL_2201 = _EVAL_3154 & _EVAL_701;
  assign _EVAL_2870 = _EVAL_1927 & _EVAL_635;
  assign _EVAL_1155 = _EVAL_3774 & _EVAL_417;
  assign _EVAL_2071 = _EVAL_268 & _EVAL_2047;
  assign _EVAL_2261 = |_EVAL_1955;
  assign _EVAL_3113 = _EVAL_409 & _EVAL_2941;
  assign _EVAL_260 = _EVAL_2532 & _EVAL_2543;
  assign _EVAL_2792 = _EVAL_2038[12];
  assign _EVAL_444 = _EVAL_3585 & _EVAL_2194;
  assign _EVAL_2126 = _EVAL_1927 & _EVAL_263;
  assign _EVAL_2656 = _EVAL_1649 & _EVAL_2906;
  assign _EVAL_3012 = _EVAL_2532 & _EVAL_2056;
  assign _EVAL_2748 = {1'h1,_EVAL_3156};
  assign _EVAL_3837 = _EVAL_1927 & _EVAL_1721;
  assign _EVAL_2706 = _EVAL_1927 & _EVAL_204;
  assign _EVAL_2125 = _EVAL_1649 & _EVAL_379;
  assign _EVAL_2741 = _EVAL_3585 & _EVAL_3232;
  assign _EVAL_3542 = _EVAL_3774 & _EVAL_370;
  assign _EVAL_1846 = _EVAL_1927 & _EVAL_1236;
  assign _EVAL_694 = _EVAL_1653 & _EVAL_2047;
  assign _EVAL_3126 = _EVAL_1410 & _EVAL_2047;
  assign _EVAL_3109 = _EVAL_1649 & _EVAL_1280;
  assign _EVAL_3168 = _EVAL_397 & _EVAL_3407;
  assign _EVAL_2847 = _EVAL_1810 & _EVAL_2047;
  assign _EVAL_821 = _EVAL_3495 & _EVAL_701;
  assign _EVAL_1463 = _EVAL_2532 & _EVAL_768;
  assign _EVAL_3314 = _EVAL_2993 & _EVAL_405;
  assign _EVAL_3215 = _EVAL_1649 & _EVAL_402;
  assign _EVAL_1305 = _EVAL_397 & _EVAL_2456;
  assign _EVAL_745 = _EVAL_2532 & _EVAL_1431;
  assign _EVAL_2546 = _EVAL_3562 & _EVAL_3224;
  assign _EVAL_1590 = _EVAL_1927 & _EVAL_2792;
  assign _EVAL_1726 = _EVAL_3125 & _EVAL_481;
  assign _EVAL_2749 = _EVAL_1927 & _EVAL_1029;
  assign _EVAL_812 = _EVAL_2587 & _EVAL_2047;
  assign _EVAL_1219 = _EVAL_2680 & _EVAL_826;
  assign _EVAL_3176 = _EVAL_3774 & _EVAL_2024;
  assign _EVAL_750 = _EVAL_2164 & _EVAL_2941;
  assign _EVAL_738 = _EVAL_2532 & _EVAL_3765;
  assign _EVAL_2420 = _EVAL_3585 & _EVAL_3606;
  assign _EVAL_3300 = |_EVAL_2797;
  assign _EVAL_773 = _EVAL_2325 & _EVAL_2047;
  assign _EVAL_2325 = _EVAL_1927 & _EVAL_2821;
  assign _EVAL_606 = _EVAL_3774 & _EVAL_1551;
  assign _EVAL_1337 = _EVAL_1927 & _EVAL_722;
  assign _EVAL_1210 = |_EVAL_380;
  assign _EVAL_3676 = _EVAL_1580 & _EVAL_2941;
  assign monitor__EVAL_5 = out_back__EVAL_7;
  assign _EVAL_1416 = _EVAL_1927 & _EVAL_2691;
  assign _EVAL_1300 = _EVAL_1296 & _EVAL_2047;
  assign _EVAL_2594 = _EVAL_1372 & _EVAL_1004;
  assign _EVAL_1961 = _EVAL_1908 & _EVAL_1004;
  assign _EVAL_2093 = _EVAL_3721 & _EVAL_701;
  assign _EVAL_3413 = _EVAL_2850[24];
  assign _EVAL_2335 = |_EVAL_1641;
  assign _EVAL_3740 = _EVAL_3333 & _EVAL_701;
  assign _EVAL_2548 = _EVAL_2038[131];
  assign _EVAL_1027 = _EVAL_1649 & _EVAL_3729;
  assign _EVAL_621 = _EVAL_2535 & _EVAL_2047;
  assign _EVAL_528 = _EVAL_1375 & _EVAL_2941;
  assign _EVAL_527 = _EVAL_1927 & _EVAL_3280;
  assign _EVAL_2046 = _EVAL_2897 & _EVAL_701;
  assign _EVAL_508 = _EVAL_3125 & _EVAL_1177;
  assign _EVAL_3558 = _EVAL_1361[10];
  assign _EVAL_413 = _EVAL_2850[18];
  assign _EVAL_1503 = _EVAL_1649 & _EVAL_416;
  assign _EVAL_3625 = _EVAL_1649 & _EVAL_2855;
  assign _EVAL_1665 = _EVAL_2038[257];
  assign _EVAL_1060 = _EVAL_1361[23:16];
  assign _EVAL_2491 = _EVAL_1927 & _EVAL_2407;
  assign _EVAL_1842 = _EVAL_3472 & _EVAL_826;
  assign _EVAL_3079 = _EVAL_3774 & _EVAL_405;
  assign _EVAL_3333 = _EVAL_2595 & _EVAL_2047;
  assign _EVAL_624 = _EVAL_1927 & _EVAL_3496;
  assign _EVAL_2709 = _EVAL_1927 & _EVAL_1028;
  assign _EVAL_2493 = _EVAL_1803 & _EVAL_826;
  assign _EVAL_2333 = _EVAL_3774 & _EVAL_1583;
  assign _EVAL_2640 = _EVAL_2038[117];
  assign _EVAL_948 = _EVAL_352 & _EVAL_826;
  assign _EVAL_3309 = _EVAL_502 & _EVAL_701;
  assign _EVAL_3010 = _EVAL_1159 & _EVAL_802;
  assign _EVAL_2818 = _EVAL_1025 & _EVAL_1004;
  assign _EVAL_2510 = _EVAL_2993 & _EVAL_2335;
  assign _EVAL_348 = _EVAL_852 & _EVAL_701;
  assign _EVAL_2169 = _EVAL_2038[97];
  assign _EVAL_3118 = _EVAL_2850[14];
  assign _EVAL_1553 = _EVAL_2656 & _EVAL_826;
  assign _EVAL_788 = _EVAL_1927 & _EVAL_3046;
  assign _EVAL_2678 = |_EVAL_307;
  assign _EVAL_2625 = _EVAL_1244 & _EVAL_826;
  assign _EVAL_2480 = _EVAL_3585 & _EVAL_2436;
  assign _EVAL_2242 = _EVAL_948 & _EVAL_2941;
  assign _EVAL_2219 = _EVAL_173 & _EVAL_2024;
  assign _EVAL_2158 = _EVAL_1361[0];
  assign _EVAL_2569 = _EVAL_2532 & _EVAL_3758;
  assign _EVAL_1803 = _EVAL_1649 & _EVAL_1763;
  assign _EVAL_682 = _EVAL_1889 & _EVAL_2047;
  assign _EVAL_2600 = _EVAL_3231 & _EVAL_2941;
  assign _EVAL_1958 = _EVAL_2459 & _EVAL_1004;
  assign _EVAL_1047 = _EVAL_1848 & _EVAL_2941;
  assign _EVAL_863 = _EVAL_220 & _EVAL_1004;
  assign _EVAL_1412 = _EVAL_2532 & _EVAL_2452;
  assign _EVAL_1295 = _EVAL_1999 & _EVAL_2047;
  assign _EVAL_2665 = _EVAL_3585 & _EVAL_2162;
  assign _EVAL_3540 = _EVAL_2038[5];
  assign _EVAL_1330 = _EVAL_2038[24];
  assign _EVAL_1215 = _EVAL_173 & _EVAL_2096;
  assign _EVAL_3796 = _EVAL_1649 & _EVAL_3747;
  assign _EVAL_601 = _EVAL_3235 & _EVAL_2047;
  assign _EVAL_2225 = _EVAL_3295 & _EVAL_701;
  assign _EVAL_3383 = _EVAL_2532 & _EVAL_974;
  assign _EVAL_3093 = _EVAL_2610 - 127'h1;
  assign _EVAL_261 = _EVAL_1927 & _EVAL_2550;
  assign _EVAL_2761 = _EVAL_2827 & _EVAL_826;
  assign _EVAL_2063 = _EVAL_3502 & _EVAL_826;
  assign _EVAL_619 = _EVAL_3125 & _EVAL_2261;
  assign _EVAL_748 = _EVAL_2883 & _EVAL_826;
  assign _EVAL_2398 = _EVAL_3432 & _EVAL_826;
  assign _EVAL_2645 = _EVAL_3556 & _EVAL_2047;
  assign _EVAL_1910 = _EVAL_2532 & _EVAL_2834;
  assign _EVAL_617 = _EVAL_3628 & _EVAL_2047;
  assign _EVAL_3565 = _EVAL_2426 & _EVAL_826;
  assign _EVAL_521 = _EVAL_173 & _EVAL_417;
  assign _EVAL_3814 = _EVAL_2598 & _EVAL_1004;
  assign _EVAL_3570 = _EVAL_2101 & _EVAL_2047;
  assign _EVAL_2602 = _EVAL_266 & _EVAL_2941;
  assign _EVAL_2731 = _EVAL_2038[121];
  assign _EVAL_2647 = _EVAL_2500 & _EVAL_1004;
  assign _EVAL_1111 = |_EVAL_1602;
  assign _EVAL_1690 = _EVAL_2532 & _EVAL_969;
  assign _EVAL_1232 = |_EVAL_3702;
  assign _EVAL_1373 = _EVAL_2188 & _EVAL_826;
  assign _EVAL_3673 = _EVAL_1560 & _EVAL_2890;
  assign _EVAL_2382 = _EVAL_3822 & _EVAL_1004;
  assign _EVAL_3484 = _EVAL_2050 & _EVAL_701;
  assign _EVAL_884 = _EVAL_3647 & _EVAL_701;
  assign _EVAL_3078 = _EVAL_1092 & _EVAL_1004;
  assign _EVAL_3790 = |_EVAL_3441;
  assign _EVAL_2681 = _EVAL_1927 & _EVAL_523;
  assign _EVAL_1508 = _EVAL_2532 & _EVAL_2640;
  assign _EVAL_1080 = _EVAL_2993 & _EVAL_3423;
  assign _EVAL_3250 = _EVAL_2850[28];
  assign monitor__EVAL_6 = _EVAL_17;
  assign _EVAL_3761 = |_EVAL_3753;
  assign _EVAL_545 = _EVAL_251 & _EVAL_701;
  assign _EVAL_2170 = _EVAL_1165 & _EVAL_701;
  assign _EVAL_537 = _EVAL_2993 & _EVAL_1986;
  assign _EVAL_1242 = _EVAL_1649 & _EVAL_1486;
  assign _EVAL_1156 = _EVAL_3507 & _EVAL_2047;
  assign _EVAL_1727 = _EVAL_3679 & _EVAL_1004;
  assign _EVAL_1110 = _EVAL_3125 & _EVAL_2162;
  assign _EVAL_3247 = _EVAL_1649 & _EVAL_3167;
  assign _EVAL_3415 = _EVAL_1405 & _EVAL_2971;
  assign _EVAL_1429 = &_EVAL_1464;
  assign _EVAL_1614 = _EVAL_3562 & _EVAL_443;
  assign _EVAL_3293 = _EVAL_2038[114];
  assign _EVAL_2950 = _EVAL_1082 & _EVAL_826;
  assign _EVAL_924 = _EVAL_397 & _EVAL_2261;
  assign _EVAL_2794 = _EVAL_2496 & _EVAL_826;
  assign _EVAL_2905 = _EVAL_1927 & _EVAL_574;
  assign _EVAL_3774 = _EVAL_1416 & _EVAL_2047;
  assign _EVAL_2543 = _EVAL_2038[85];
  assign _EVAL_885 = _EVAL_173 & _EVAL_3810;
  assign _EVAL_1721 = _EVAL_2038[79];
  assign _EVAL_375 = _EVAL_3050 & _EVAL_826;
  assign _EVAL_2522 = _EVAL_3774 & _EVAL_2335;
  assign _EVAL_470 = _EVAL_2532 & _EVAL_1619;
  assign _EVAL_1188 = _EVAL_3562 & _EVAL_3272;
  assign _EVAL_3682 = _EVAL_2448 & _EVAL_2047;
  assign _EVAL_690 = _EVAL_882 & _EVAL_3120;
  assign _EVAL_1913 = _EVAL_3562 & _EVAL_2162;
  assign _EVAL_391 = _EVAL_2532 & _EVAL_1029;
  assign _EVAL_2013 = _EVAL_2532 & _EVAL_2826;
  assign _EVAL_1941 = _EVAL_1927 & _EVAL_2223;
  assign _EVAL_795 = _EVAL_3585 & _EVAL_3761;
  assign _EVAL_2785 = _EVAL_3294 & _EVAL_1004;
  assign _EVAL_2646 = _EVAL_3126 & _EVAL_3810;
  assign _EVAL_2751 = _EVAL_2802 & _EVAL_2941;
  assign _EVAL_1197 = _EVAL_483 & _EVAL_2047;
  assign _EVAL_901 = _EVAL_940 & _EVAL_701;
  assign _EVAL_271 = _EVAL_2038[112];
  assign _EVAL_1851 = _EVAL_310 & _EVAL_826;
  assign _EVAL_3453 = _EVAL_3562 & _EVAL_3764;
  assign _EVAL_1376 = _EVAL_3774 & _EVAL_1986;
  assign _EVAL_3630 = _EVAL_2038[53];
  assign _EVAL_162 = _EVAL_3254 & _EVAL_2941;
  assign _EVAL_1279 = _EVAL_3562 & _EVAL_3761;
  assign _EVAL_3816 = _EVAL_2405 & _EVAL_2047;
  assign _EVAL_2933 = _EVAL_1927 & _EVAL_720;
  assign _EVAL_3332 = ~_EVAL_110;
  assign _EVAL_243 = _EVAL_2038[61];
  assign _EVAL_1977 = _EVAL_2532 & _EVAL_2301;
  assign _EVAL_3022 = _EVAL_717 & _EVAL_1429;
  assign _EVAL_2839 = _EVAL_1927 & _EVAL_187;
  assign _EVAL_3292 = _EVAL_1649 & _EVAL_506;
  assign _EVAL_947 = ~_EVAL_2116;
  assign _EVAL_754 = _EVAL_3774 & _EVAL_3854;
  assign _EVAL_3226 = _EVAL_1361[14];
  assign _EVAL_1950 = _EVAL_2038[14];
  assign _EVAL_2512 = _EVAL_1770 & _EVAL_2047;
  assign _EVAL_2754 = _EVAL_2038[256];
  assign _EVAL_3054 = _EVAL_1996 & _EVAL_2047;
  assign _EVAL_3586 = _EVAL_717 & _EVAL_3233;
  assign monitor__EVAL_2 = out_back__EVAL_11;
  assign _EVAL_1204 = _EVAL_397 & _EVAL_3790;
  assign _EVAL_702 = _EVAL_823 & _EVAL_2047;
  assign _EVAL_2292 = _EVAL_1091 & _EVAL_2047;
  assign _EVAL_1348 = ~_EVAL_1393;
  assign _EVAL_2259 = _EVAL_1679 & _EVAL_1004;
  assign _EVAL_3092 = _EVAL_2532 & _EVAL_3821;
  assign _EVAL_1992 = _EVAL_173 & _EVAL_2678;
  assign _EVAL_3675 = _EVAL_738 & _EVAL_2047;
  assign _EVAL_2250 = _EVAL_3666 & _EVAL_826;
  assign _EVAL_359 = _EVAL_1766 & _EVAL_2047;
  assign _EVAL_2104 = _EVAL_2532 & _EVAL_3132;
  assign monitor__EVAL_10 = _EVAL_136;
  assign _EVAL_3808 = _EVAL_2038[258];
  assign _EVAL_722 = _EVAL_2038[90];
  assign _EVAL_756 = _EVAL_1800 & _EVAL_2047;
  assign _EVAL_564 = _EVAL_1927 & _EVAL_1497;
  assign _EVAL_2497 = _EVAL_1313 & _EVAL_2941;
  assign _EVAL_2449 = _EVAL_1927 & _EVAL_3132;
  assign _EVAL_1772 = _EVAL_3126 & _EVAL_2678;
  assign _EVAL_2563 = _EVAL_1927 & _EVAL_1316;
  assign _EVAL_493 = _EVAL_1095 & _EVAL_2941;
  assign _EVAL_3514 = _EVAL_1927 & _EVAL_3818;
  assign _EVAL_1273 = _EVAL_3125 & _EVAL_3252;
  assign _EVAL_3634 = _EVAL_3585 & _EVAL_3764;
  assign _EVAL_1991 = _EVAL_303 & _EVAL_701;
  assign _EVAL_3459 = _EVAL_207 & _EVAL_2047;
  assign _EVAL_1456 = ~_EVAL_1777;
  assign _EVAL_1612 = _EVAL_1503 & _EVAL_826;
  assign _EVAL_169 = _EVAL_486 & _EVAL_2047;
  assign _EVAL_3279 = _EVAL_2038[27];
  assign _EVAL_452 = _EVAL_3562 & _EVAL_3252;
  assign _EVAL_2898 = _EVAL_2038[69];
  assign _EVAL_1173 = _EVAL_2532 & _EVAL_2411;
  assign _EVAL_519 = _EVAL_351 & _EVAL_2941;
  assign _EVAL_1575 = _EVAL_277 & _EVAL_2026;
  assign _EVAL_3062 = _EVAL_1553 & _EVAL_2941;
  assign _EVAL_417 = |_EVAL_3085;
  assign _EVAL_1654 = _EVAL_2048 & _EVAL_1004;
  assign _EVAL_3360 = _EVAL_2532 & _EVAL_2187;
  assign _EVAL_3561 = _EVAL_874 & _EVAL_2047;
  assign _EVAL_2535 = _EVAL_1927 & _EVAL_3258;
  assign _EVAL_1068 = _EVAL_1842 & _EVAL_2941;
  assign _EVAL_3473 = _EVAL_2775[2];
  assign _EVAL_235 = _EVAL_2532 & _EVAL_1887;
  assign _EVAL_2884 = _EVAL_3126 & _EVAL_2635;
  assign _EVAL_2326 = _EVAL_1649 & _EVAL_1973;
  assign _EVAL_1225 = _EVAL_3125 & _EVAL_2908;
  assign _EVAL_3429 = {_EVAL_1141,_EVAL_3128,_EVAL_216,_EVAL_3687,_EVAL_2508,_EVAL_2714,_EVAL_542,_EVAL_3473,_EVAL_2464,
    _EVAL_1285};
  assign _EVAL_1216 = _EVAL_3585 & _EVAL_942;
  assign _EVAL_807 = _EVAL_1361[19];
  assign _EVAL_1157 = _EVAL_1927 & _EVAL_985;
  assign _EVAL_2815 = _EVAL_173 & _EVAL_3703;
  assign _EVAL_3496 = _EVAL_2038[42];
  assign _EVAL_3778 = _EVAL_1561 & _EVAL_2047;
  assign _EVAL_248 = _EVAL_2532 & _EVAL_464;
  assign _EVAL_2920 = _EVAL_740 & _EVAL_701;
  assign _EVAL_1636 = _EVAL_2532 & _EVAL_2573;
  assign _EVAL_3741 = _EVAL_1927 & _EVAL_3630;
  assign _EVAL_277 = _EVAL_2125 & _EVAL_826;
  assign _EVAL_2475 = _EVAL_3669 & _EVAL_701;
  assign _EVAL_1192 = _EVAL_2532 & _EVAL_1650;
  assign _EVAL_3282 = _EVAL_3298 & _EVAL_1004;
  assign _EVAL_912 = _EVAL_3178 & _EVAL_1004;
  assign _EVAL_1646 = _EVAL_1361[22];
  assign _EVAL_3380 = _EVAL_2901 & _EVAL_701;
  assign _EVAL_3539 = _EVAL_2993 & _EVAL_1223;
  assign _EVAL_3730 = _EVAL_217 & _EVAL_2941;
  assign _EVAL_3447 = _EVAL_717 & _EVAL_3830;
  assign _EVAL_3738 = _EVAL_2993 & _EVAL_2780;
  assign _EVAL_3234 = _EVAL_2953 & _EVAL_826;
  assign _EVAL_3445 = _EVAL_1137 & _EVAL_701;
  assign _EVAL_543 = _EVAL_1649 & _EVAL_838;
  assign _EVAL_2072 = _EVAL_617 & _EVAL_701;
  assign _EVAL_2394 = _EVAL_2532 & _EVAL_2359;
  assign _EVAL_3846 = _EVAL_6 == 3'h4;
  assign _EVAL_1106 = _EVAL_1649 & _EVAL_3319;
  assign _EVAL_2876 = _EVAL_2867 & _EVAL_1004;
  assign _EVAL_654 = _EVAL_2684 & _EVAL_1811;
  assign _EVAL_2560 = _EVAL_3125 & _EVAL_3606;
  assign _EVAL_2033 = |_EVAL_413;
  assign _EVAL_2778 = _EVAL_3607 & _EVAL_2047;
  assign _EVAL_3660 = _EVAL_1629 & _EVAL_826;
  assign _EVAL_802 = |_EVAL_1060;
  assign _EVAL_2775 = _EVAL_2478[19:0];
  assign _EVAL_3018 = _EVAL_2128 & _EVAL_2047;
  assign _EVAL_298 = _EVAL_2532 & _EVAL_2169;
  assign _EVAL_591 = _EVAL_2532 & _EVAL_2445;
  assign _EVAL_2265 = _EVAL_1271 & _EVAL_1004;
  assign _EVAL_1970 = _EVAL_2850[13];
  assign _EVAL_857 = _EVAL_2434 & _EVAL_701;
  assign _EVAL_2163 = _EVAL_2532 & _EVAL_3496;
  assign _EVAL_3441 = _EVAL_2850[2];
  assign _EVAL_2135 = _EVAL_3098 & _EVAL_2047;
  assign _EVAL_1272 = _EVAL_2850[25];
  assign _EVAL_3753 = _EVAL_2850[7];
  assign _EVAL_1538 = _EVAL_397 & _EVAL_3649;
  assign _EVAL_2670 = _EVAL_2532 & _EVAL_650;
  assign _EVAL_2256 = _EVAL_2491 & _EVAL_2047;
  assign _EVAL_1298 = _EVAL_2373 & _EVAL_2047;
  assign _EVAL_763 = _EVAL_3377 & _EVAL_826;
  assign _EVAL_1037 = _EVAL_2139 & _EVAL_2941;
  assign _EVAL_3396 = _EVAL_1114 & _EVAL_2047;
  assign _EVAL_1588 = _EVAL_525 & _EVAL_2047;
  assign _EVAL_441 = _EVAL_1405 & _EVAL_3233;
  assign _EVAL_2243 = _EVAL_1927 & _EVAL_2169;
  assign _EVAL_589 = _EVAL_791 & _EVAL_2047;
  assign _EVAL_2840 = _EVAL_2184 & _EVAL_826;
  assign _EVAL_1231 = _EVAL_3562 & _EVAL_1930;
  assign _EVAL_2954 = _EVAL_2603 & _EVAL_1004;
  assign _EVAL_1878 = _EVAL_2937 & _EVAL_2047;
  assign _EVAL_3830 = &_EVAL_1060;
  assign monitor__EVAL_11 = out_back__EVAL_2;
  assign _EVAL_149 = |_EVAL_1361;
  assign _EVAL_2357 = _EVAL_1556 & _EVAL_2941;
  assign _EVAL_658 = _EVAL_1018 & _EVAL_701;
  assign _EVAL_879 = _EVAL_1927 & _EVAL_2754;
  assign _EVAL_360 = _EVAL_3003 & _EVAL_826;
  assign _EVAL_3767 = _EVAL_2038[31];
  assign _EVAL_1543 = _EVAL_1649 & _EVAL_3524;
  assign _EVAL_1332 = _EVAL_2532 & _EVAL_2962;
  assign _EVAL_1917 = _EVAL_2123 & _EVAL_3841;
  assign _EVAL_2726 = _EVAL_2038[95];
  assign _EVAL_1344 = _EVAL_3234 & _EVAL_2941;
  assign _EVAL_717 = _EVAL_438 & _EVAL_2047;
  assign _EVAL_1967 = _EVAL_2532 & _EVAL_1566;
  assign _EVAL_1586 = _EVAL_3126 & _EVAL_2096;
  assign _EVAL_877 = _EVAL_512 & _EVAL_2047;
  assign _EVAL_2797 = _EVAL_2850[22];
  assign _EVAL_2006 = _EVAL_3829 & _EVAL_1004;
  assign _EVAL_2532 = _EVAL_159 & _EVAL_1113;
  assign _EVAL_3208 = _EVAL_147 & _EVAL_2941;
  assign _EVAL_3500 = _EVAL_359 & _EVAL_701;
  assign _EVAL_1455 = _EVAL_2532 & _EVAL_698;
  assign _EVAL_1557 = _EVAL_1625 & _EVAL_826;
  assign _EVAL_1619 = _EVAL_2038[122];
  assign _EVAL_2288 = _EVAL_3238 & _EVAL_2047;
  assign _EVAL_2939 = _EVAL_3562 & _EVAL_3606;
  assign _EVAL_1424 = _EVAL_2532 & _EVAL_1370;
  assign _EVAL_1487 = _EVAL_1784 & _EVAL_2047;
  assign _EVAL_2082 = _EVAL_484 & _EVAL_2941;
  assign _EVAL_2958 = _EVAL_1895 & _EVAL_1004;
  assign _EVAL_1951 = _EVAL_3512 & _EVAL_1004;
  assign _EVAL_2591 = _EVAL_2563 & _EVAL_2047;
  assign _EVAL_1921 = _EVAL_1814 & _EVAL_2047;
  assign _EVAL_1129 = _EVAL_2038[46];
  assign _EVAL_1397 = _EVAL_3781 & _EVAL_1526;
  assign _EVAL_2136 = _EVAL_2836 & _EVAL_2047;
  assign _EVAL_1491 = _EVAL_173 & _EVAL_1986;
  assign _EVAL_3369 = _EVAL_2038[512];
  assign _EVAL_2834 = _EVAL_2038[30];
  assign _EVAL_818 = _EVAL_3625 & _EVAL_826;
  assign _EVAL_3773 = _EVAL_875 & _EVAL_826;
  assign _EVAL_3323 = _EVAL_2850[8];
  assign _EVAL_1840 = _EVAL_1943 & _EVAL_2047;
  assign _EVAL_3839 = _EVAL_1306 & _EVAL_2941;
  assign _EVAL_351 = _EVAL_1126 & _EVAL_826;
  assign _EVAL_3554 = _EVAL_1649 & _EVAL_160;
  assign _EVAL_1533 = _EVAL_1798 & _EVAL_2047;
  assign _EVAL_1845 = _EVAL_3126 & _EVAL_2024;
  assign _EVAL_1931 = _EVAL_1348 | _EVAL_110;
  assign _EVAL_3780 = _EVAL_3584 ? 8'hff : 8'h0;
  assign _EVAL_2529 = _EVAL_1317 & _EVAL_826;
  assign _EVAL_1835 = _EVAL_1361[29];
  assign _EVAL_2930 = _EVAL_397 & _EVAL_1177;
  assign _EVAL_2157 = _EVAL_1786 & _EVAL_2047;
  assign _EVAL_2514 = _EVAL_1649 & _EVAL_3255;
  assign _EVAL_2032 = _EVAL_2778 & _EVAL_1004;
  assign _EVAL_2038 = 1024'h1 << _EVAL_3429;
  assign _EVAL_1887 = _EVAL_2038[54];
  assign _EVAL_1895 = _EVAL_1058 & _EVAL_2047;
  assign _EVAL_373 = _EVAL_1649 & _EVAL_560;
  assign _EVAL_3598 = _EVAL_2847 & _EVAL_1004;
  assign _EVAL_188 = _EVAL_2038[109];
  assign _EVAL_3512 = _EVAL_2240 & _EVAL_2047;
  assign _EVAL_1383 = _EVAL_1159 & _EVAL_3605;
  assign _EVAL_623 = _EVAL_1927 & _EVAL_1330;
  assign _EVAL_2235 = |_EVAL_1970;
  assign _EVAL_262 = _EVAL_2641 & _EVAL_1004;
  assign _EVAL_2790 = _EVAL_2528 & _EVAL_701;
  assign _EVAL_2837 = _EVAL_2400 & _EVAL_1004;
  assign _EVAL_1625 = _EVAL_1649 & _EVAL_2865;
  assign _EVAL_525 = _EVAL_2532 & _EVAL_935;
  assign _EVAL_1351 = _EVAL_1927 & _EVAL_2640;
  assign _EVAL_2066 = _EVAL_397 & _EVAL_3232;
  assign _EVAL_419 = _EVAL_1201 & _EVAL_826;
  assign _EVAL_308 = _EVAL_1927 & _EVAL_549;
  assign _EVAL_1389 = _EVAL_2816 & _EVAL_2941;
  assign _EVAL_1778 = _EVAL_1059 & _EVAL_2941;
  assign _EVAL_684 = _EVAL_785 & _EVAL_1232;
  assign _EVAL_1196 = _EVAL_3126 & _EVAL_3854;
  assign _EVAL_1643 = _EVAL_2850[23];
  assign _EVAL_430 = _EVAL_1589 & _EVAL_826;
  assign _EVAL_2421 = _EVAL_1649 & _EVAL_3343;
  assign _EVAL_1236 = _EVAL_2038[35];
  assign _EVAL_1894 = _EVAL_2769 & _EVAL_2047;
  assign _EVAL_1063 = _EVAL_3837 & _EVAL_2047;
  assign _EVAL_3781 = _EVAL_2757 > 7'h8;
  assign _EVAL_1582 = _EVAL_1927 & _EVAL_3421;
  assign _EVAL_2452 = _EVAL_2038[71];
  assign _EVAL_548 = _EVAL_1897 & _EVAL_3605;
  assign _EVAL_2286 = _EVAL_455 & _EVAL_2047;
  assign _EVAL_3677 = _EVAL_1993 & _EVAL_1004;
  assign _EVAL_3580 = _EVAL_2532 & _EVAL_1950;
  assign _EVAL_1583 = |_EVAL_2893;
  assign _EVAL_3230 = _EVAL_397 & _EVAL_1245;
  assign _EVAL_1479 = _EVAL_1501 & _EVAL_826;
  assign _EVAL_1891 = _EVAL_2532 & _EVAL_3184;
  assign _EVAL_2010 = _EVAL_3585 & _EVAL_3272;
  assign _EVAL_896 = _EVAL_2071 & _EVAL_701;
  assign _EVAL_1108 = _EVAL_433 & _EVAL_1004;
  assign _EVAL_220 = _EVAL_3406 & _EVAL_2047;
  assign _EVAL_1493 = _EVAL_598 & _EVAL_2047;
  assign _EVAL_432 = _EVAL_3788 & _EVAL_2941;
  assign _EVAL_3601 = _EVAL_3562 & _EVAL_2908;
  assign _EVAL_266 = _EVAL_2463 & _EVAL_826;
  assign _EVAL_2429 = _EVAL_1967 & _EVAL_2047;
  assign _EVAL_3137 = _EVAL_3562 & _EVAL_2194;
  assign _EVAL_2984 = _EVAL_2940 & _EVAL_826;
  assign _EVAL_2461 = _EVAL_3041 & _EVAL_2047;
  assign _EVAL_579 = _EVAL_747 & _EVAL_701;
  assign _EVAL_805 = _EVAL_84[1];
  assign _EVAL_2188 = _EVAL_1649 & _EVAL_2814;
  assign _EVAL_1168 = _EVAL_2993 & _EVAL_2487;
  assign _EVAL_178 = _EVAL_2993 & _EVAL_1125;
  assign _EVAL_2371 = _EVAL_397 & _EVAL_2194;
  assign _EVAL_1515 = _EVAL_1940 & _EVAL_2047;
  assign _EVAL_550 = _EVAL_2461 & _EVAL_1004;
  assign _EVAL_2137 = _EVAL_1649 & _EVAL_3243;
  assign _EVAL_2897 = _EVAL_952 & _EVAL_2047;
  assign _EVAL_554 = _EVAL_2287 & _EVAL_2047;
  assign _EVAL_1628 = _EVAL_3562 & _EVAL_846;
  assign _EVAL_866 = _EVAL_1927 & _EVAL_464;
  assign _EVAL_455 = _EVAL_1927 & _EVAL_2445;
  assign _EVAL_2187 = _EVAL_2038[119];
  assign _EVAL_1432 = _EVAL_2532 & _EVAL_2792;
  assign _EVAL_1996 = _EVAL_2532 & _EVAL_329;
  assign _EVAL_447 = _EVAL_397 & _EVAL_2436;
  assign _EVAL_2570 = _EVAL_328 & _EVAL_826;
  assign _EVAL_1266 = _EVAL_3126 & _EVAL_1125;
  assign _EVAL_1574 = _EVAL_1258 & _EVAL_2941;
  assign _EVAL_242 = _EVAL_2532 & _EVAL_1205;
  assign _EVAL_2581 = _EVAL_2835 & _EVAL_2047;
  assign _EVAL_1223 = |_EVAL_2393;
  assign _EVAL_287 = _EVAL_3470 & _EVAL_2047;
  assign _EVAL_3424 = _EVAL_3562 & _EVAL_2456;
  assign _EVAL_2708 = _EVAL_2808 & _EVAL_826;
  assign _EVAL_1786 = _EVAL_2532 & _EVAL_574;
  assign _EVAL_503 = _EVAL_1682 & _EVAL_701;
  assign _EVAL_708 = _EVAL_1063 & _EVAL_1004;
  assign _EVAL_2506 = _EVAL_1557 & _EVAL_2941;
  assign _EVAL_2351 = _EVAL_546 & _EVAL_2941;
  assign _EVAL_400 = _EVAL_1927 & _EVAL_3710;
  assign _EVAL_3248 = _EVAL_2127 & _EVAL_2941;
  assign _EVAL_846 = |_EVAL_1734;
  assign _EVAL_3169 = {{3'd0}, _EVAL_2748};
  assign _EVAL_1207 = _EVAL_2755 & _EVAL_701;
  assign _EVAL_2807 = _EVAL_993 & _EVAL_1004;
  assign _EVAL_3690 = _EVAL_3092 & _EVAL_2047;
  assign _EVAL_2401 = _EVAL_1322 & _EVAL_2941;
  assign _EVAL_3403 = _EVAL_1361[2:0];
  assign _EVAL_2674 = _EVAL_2891 & _EVAL_826;
  assign _EVAL_1770 = _EVAL_2532 & _EVAL_722;
  assign _EVAL_3016 = _EVAL_1229 & _EVAL_826;
  assign _EVAL_2962 = _EVAL_2038[4];
  assign _EVAL_3277 = _EVAL_2364 & _EVAL_2941;
  assign _EVAL_1915 = _EVAL_1927 & _EVAL_1129;
  assign _EVAL_2255 = _EVAL_2038[48];
  assign _EVAL_1766 = _EVAL_2532 & _EVAL_1316;
  assign _EVAL_2228 = _EVAL_1454 & _EVAL_826;
  assign _EVAL_1651 = _EVAL_1492 & _EVAL_1004;
  assign _EVAL_2445 = _EVAL_2038[80];
  assign _EVAL_2967 = _EVAL_1671 & _EVAL_2941;
  assign _EVAL_1244 = _EVAL_1649 & _EVAL_3099;
  assign _EVAL_2128 = _EVAL_1927 & _EVAL_2056;
  assign _EVAL_1044 = _EVAL_3018 & _EVAL_1004;
  assign _EVAL_2809 = _EVAL_1870 & _EVAL_826;
  assign _EVAL_2050 = _EVAL_211 & _EVAL_2047;
  assign _EVAL_2597 = _EVAL_1335 & _EVAL_2047;
  assign _EVAL_2752 = _EVAL_3585 & _EVAL_481;
  assign _EVAL_1620 = _EVAL_3690 & _EVAL_701;
  assign _EVAL_1522 = _EVAL_1487 & _EVAL_701;
  assign _EVAL_1791 = _EVAL_1212 & _EVAL_1004;
  assign _EVAL_3421 = _EVAL_2038[67];
  assign _EVAL_1189 = _EVAL_1337 & _EVAL_2047;
  assign _EVAL_387 = _EVAL_1067 & _EVAL_2941;
  assign _EVAL_1064 = _EVAL_3741 & _EVAL_2047;
  assign _EVAL_1981 = _EVAL_1649 & _EVAL_2624;
  assign _EVAL_1230 = _EVAL_3749 & _EVAL_3087;
  assign _EVAL_586 = _EVAL_1361[7];
  assign _EVAL_972 = _EVAL_3016 & _EVAL_2941;
  assign _EVAL_305 = _EVAL_3585 & _EVAL_2456;
  assign _EVAL_785 = _EVAL_349 & _EVAL_826;
  assign _EVAL_1059 = _EVAL_1345 & _EVAL_826;
  assign _EVAL_507 = |_EVAL_3313;
  assign _EVAL_3679 = _EVAL_3648 & _EVAL_2047;
  assign _EVAL_1121 = _EVAL_601 & _EVAL_1004;
  assign _EVAL_3452 = _EVAL_3125 & _EVAL_3649;
  assign monitor__EVAL_7 = _EVAL_70;
  assign _EVAL_2909 = _EVAL_2123 & _EVAL_3724;
  assign _EVAL_2995 = _EVAL_1649 & _EVAL_840;
  assign _EVAL_2664 = _EVAL_3125 & _EVAL_1111;
  assign _EVAL_946 = _EVAL_1927 & _EVAL_3184;
  assign _EVAL_961 = _EVAL_1995 & _EVAL_1004;
  assign _EVAL_3053 = _EVAL_397 & _EVAL_3272;
  assign _EVAL_3313 = _EVAL_2850[31:3];
  assign _EVAL_3792 = _EVAL_2038[11];
  assign _EVAL_3091 = _EVAL_3126 & _EVAL_2541;
  assign _EVAL_2783 = _EVAL_2532 & _EVAL_511;
  assign _EVAL_2916 = _EVAL_3774 & _EVAL_290;
  assign _EVAL_2044 = _EVAL_1804 & _EVAL_1004;
  assign _EVAL_1810 = _EVAL_1927 & _EVAL_3279;
  assign _EVAL_2723 = _EVAL_1977 & _EVAL_2047;
  assign _EVAL_1906 = _EVAL_565 & _EVAL_2941;
  assign _EVAL_1109 = _EVAL_943 & _EVAL_701;
  assign _EVAL_3364 = _EVAL_2157 & _EVAL_701;
  assign _EVAL_2443 = _EVAL_397 & _EVAL_1111;
  assign _EVAL_1652 = _EVAL_2894 & _EVAL_1004;
  assign _EVAL_2432 = _EVAL_2993 & _EVAL_3549;
  assign _EVAL_1468 = _EVAL_1186 & _EVAL_701;
  assign _EVAL_327 = _EVAL_3126 & _EVAL_1583;
  assign _EVAL_3810 = |_EVAL_3783;
  assign _EVAL_835 = _EVAL_2161 & _EVAL_2941;
  assign _EVAL_2489 = _EVAL_2135 & _EVAL_701;
  assign _EVAL_935 = _EVAL_2038[72];
  assign _EVAL_2813 = _EVAL_246 & _EVAL_2047;
  assign _EVAL_2245 = _EVAL_1543 & _EVAL_826;
  assign _EVAL_3506 = _EVAL_1649 & _EVAL_1090;
  assign _EVAL_676 = _EVAL_663 & _EVAL_701;
  assign _EVAL_3116 = _EVAL_1736 & _EVAL_2047;
  assign _EVAL_874 = _EVAL_1927 & _EVAL_457;
  assign _EVAL_2317 = _EVAL_2038[18];
  assign _EVAL_1370 = _EVAL_2038[59];
  assign _EVAL_3090 = _EVAL_2404 & _EVAL_1004;
  assign _EVAL_2964 = _EVAL_1917 & _EVAL_1581;
  assign _EVAL_2283 = _EVAL_397 & _EVAL_914;
  assign _EVAL_1808 = _EVAL_2356 & _EVAL_3233;
  assign _EVAL_1563 = _EVAL_3125 & _EVAL_942;
  assign _EVAL_927 = _EVAL_2831 & _EVAL_826;
  assign _EVAL_3224 = |_EVAL_919;
  assign _EVAL_3509 = _EVAL_2704 & _EVAL_1004;
  assign _EVAL_2505 = _EVAL_1927 & _EVAL_1566;
  assign _EVAL_1318 = _EVAL_2038[7];
  assign _EVAL_1980 = _EVAL_2388 & _EVAL_1004;
  assign _EVAL_1933 = _EVAL_1716 & _EVAL_701;
  assign _EVAL_3160 = _EVAL_3126 & _EVAL_1551;
  assign _EVAL_1131 = _EVAL_1649 & _EVAL_212;
  assign _EVAL_749 = _EVAL_3562 & _EVAL_1275;
  assign _EVAL_1823 = _EVAL_3126 & _EVAL_1470;
  assign _EVAL_1217 = _EVAL_2993 & _EVAL_290;
  assign _EVAL_2620 = _EVAL_589 & _EVAL_701;
  assign _EVAL_926 = _EVAL_1649 & _EVAL_1877;
  assign _EVAL_1247 = _EVAL_1649 & _EVAL_2027;
  assign monitor__EVAL_4 = _EVAL_6;
  assign _EVAL_1464 = _EVAL_1361[31:24];
  assign _EVAL_1265 = _EVAL_986 & _EVAL_2047;
  assign _EVAL_3823 = _EVAL_2038[63];
  assign _EVAL_3239 = _EVAL_781 & _EVAL_2047;
  assign _EVAL_1600 = _EVAL_1927 & _EVAL_2185;
  assign _EVAL_3709 = _EVAL_2038[26];
  assign _EVAL_194 = _EVAL_3044 ? 8'hff : 8'h0;
  assign _EVAL_3563 = _EVAL_877 & _EVAL_701;
  assign _EVAL_734 = _EVAL_3774 & _EVAL_1125;
  assign _EVAL_2463 = _EVAL_1649 & _EVAL_2220;
  assign _EVAL_895 = _EVAL_1927 & _EVAL_935;
  assign _EVAL_2744 = _EVAL_3126 & _EVAL_290;
  assign _EVAL_1477 = _EVAL_2228 & _EVAL_2941;
  assign _EVAL_3131 = _EVAL_661 & _EVAL_1004;
  assign _EVAL_1285 = _EVAL_2775[0];
  assign _EVAL_2302 = _EVAL_2532 & _EVAL_1028;
  assign _EVAL_2209 = _EVAL_1649 & _EVAL_2484;
  assign _EVAL_2820 = _EVAL_173 & _EVAL_3854;
  assign _EVAL_1523 = _EVAL_1361[16];
  assign _EVAL_1105 = _EVAL_3126 & _EVAL_1478;
  assign _EVAL_2173 = _EVAL_2326 & _EVAL_826;
  assign _EVAL_1384 = _EVAL_1649 & _EVAL_3384;
  assign _EVAL_2339 = _EVAL_1649 & _EVAL_1830;
  assign _EVAL_1162 = _EVAL_2532 & _EVAL_3258;
  assign _EVAL_3546 = _EVAL_1163 & _EVAL_2047;
  assign _EVAL_2707 = _EVAL_1649 & _EVAL_2346;
  assign _EVAL_426 = _EVAL_1277 & _EVAL_701;
  assign _EVAL_2446 = _EVAL_1361[4];
  assign _EVAL_1598 = _EVAL_2038[37];
  assign _EVAL_1844 = _EVAL_3143 & _EVAL_826;
  assign _EVAL_2827 = _EVAL_1649 & _EVAL_1354;
  assign _EVAL_951 = _EVAL_2532 & _EVAL_2566;
  assign _EVAL_800 = _EVAL_2943 & _EVAL_1004;
  assign _EVAL_511 = _EVAL_2038[44];
  assign _EVAL_1327 = _EVAL_3774 & _EVAL_2780;
  assign _EVAL_3573 = _EVAL_718 & _EVAL_2047;
  assign _EVAL_3779 = _EVAL_1084 & _EVAL_1004;
  assign _EVAL_556 = _EVAL_1582 & _EVAL_2047;
  assign _EVAL_3623 = _EVAL_3126 & _EVAL_1223;
  assign _EVAL_3066 = _EVAL_3448 & _EVAL_2047;
  assign _EVAL_2471 = _EVAL_1649 & _EVAL_2798;
  assign _EVAL_2721 = _EVAL_2850[5];
  assign _EVAL_3338 = _EVAL_2363 & _EVAL_2941;
  assign _EVAL_420 = _EVAL_173 & _EVAL_1868;
  assign _EVAL_2002 = _EVAL_651[130];
  assign _EVAL_538 = _EVAL_557 & _EVAL_826;
  assign _EVAL_1756 = _EVAL_2212 & _EVAL_1004;
  assign _EVAL_2358 = _EVAL_2993 & _EVAL_3498;
  assign _EVAL_2007 = _EVAL_2413 & _EVAL_2047;
  assign _EVAL_2959 = _EVAL_250 & _EVAL_701;
  assign _EVAL_3117 = _EVAL_3774 & _EVAL_2447;
  assign _EVAL_1381 = _EVAL_2532 & _EVAL_475;
  assign _EVAL_2583 = _EVAL_3697 & _EVAL_1004;
  assign _EVAL_2895 = _EVAL_2850[29];
  assign _EVAL_3817 = _EVAL_2544 & _EVAL_826;
  assign _EVAL_3274 = _EVAL_1927 & _EVAL_2543;
  assign _EVAL_2229 = _EVAL_1420 & _EVAL_701;
  assign _EVAL_774 = _EVAL_2138 & _EVAL_826;
  assign _EVAL_3724 = _EVAL_3776[0];
  assign _EVAL_549 = _EVAL_2038[98];
  assign _EVAL_3818 = _EVAL_2038[29];
  assign _EVAL_1829 = _EVAL_173 & _EVAL_2541;
  assign _EVAL_3371 = _EVAL_2250 & _EVAL_2941;
  assign _EVAL_1152 = _EVAL_843 & _EVAL_701;
  assign _EVAL_311 = _EVAL_277 & _EVAL_1811;
  assign _EVAL_3482 = _EVAL_3774 & _EVAL_1478;
  assign _EVAL_3464 = _EVAL_2137 & _EVAL_826;
  assign _EVAL_1635 = _EVAL_2038[55];
  assign _EVAL_2991 = _EVAL_1927 & _EVAL_2643;
  assign _EVAL_3748 = _EVAL_1927 & _EVAL_398;
  assign _EVAL_2115 = _EVAL_1361[7:1];
  assign _EVAL_535 = _EVAL_1927 & _EVAL_1598;
  assign _EVAL_1816 = _EVAL_2156 & _EVAL_436;
  assign _EVAL_1571 = |_EVAL_824;
  assign _EVAL_1633 = _EVAL_2703 & _EVAL_826;
  assign _EVAL_2447 = |_EVAL_3558;
  assign _EVAL_3710 = _EVAL_2038[22];
  assign _EVAL_159 = _EVAL_5 & _EVAL_3491;
  assign _EVAL_3584 = _EVAL_84[3];
  assign monitor__EVAL = _EVAL_130;
  assign _EVAL_3301 = _EVAL_3769 & _EVAL_2047;
  assign _EVAL_1513 = _EVAL_2120 & _EVAL_1429;
  assign _EVAL_3356 = _EVAL_3126 & _EVAL_1708;
  assign _EVAL_999 = _EVAL_1649 & _EVAL_2375;
  assign _EVAL_2573 = _EVAL_2038[68];
  assign _EVAL_1839 = _EVAL_1361[18];
  assign _EVAL_1404 = _EVAL_581 & _EVAL_2047;
  assign _EVAL_2526 = _EVAL_2215 & _EVAL_2941;
  assign _EVAL_3493 = _EVAL_2532 & _EVAL_3308;
  assign _EVAL_2899 = _EVAL_621 & _EVAL_1004;
  assign _EVAL_443 = |_EVAL_3833;
  assign _EVAL_1294 = _EVAL_1927 & _EVAL_1318;
  assign _EVAL_1484 = _EVAL_287 & _EVAL_1004;
  assign _EVAL_2887 = _EVAL_2605 & _EVAL_701;
  assign _EVAL_3771 = _EVAL_3125 & _EVAL_3232;
  assign _EVAL_2541 = |_EVAL_1835;
  assign _EVAL_1776 = _EVAL_686 & _EVAL_826;
  assign _EVAL_263 = _EVAL_2038[6];
  assign _EVAL_1873 = _EVAL_2850[12];
  assign _EVAL_2528 = _EVAL_391 & _EVAL_2047;
  assign _EVAL_1856 = _EVAL_1649 & _EVAL_3206;
  assign _EVAL_3758 = _EVAL_2038[16];
  assign _EVAL_2430 = _EVAL_3125 & _EVAL_1275;
  assign _EVAL_2029 = _EVAL_2532 & _EVAL_226;
  assign _EVAL_1335 = _EVAL_1927 & _EVAL_974;
  assign _EVAL_3585 = _EVAL_1119 & _EVAL_826;
  assign _EVAL_3298 = _EVAL_479 & _EVAL_2047;
  assign _EVAL_530 = _EVAL_186 & _EVAL_2941;
  assign _EVAL_1926 = _EVAL_1927 & _EVAL_1370;
  assign _EVAL_1048 = _EVAL_931 & _EVAL_826;
  assign _EVAL_3228 = _EVAL_1156 & _EVAL_701;
  assign _EVAL_1848 = _EVAL_2421 & _EVAL_826;
  assign _EVAL_3273 = _EVAL_829 & _EVAL_826;
  assign _EVAL_1526 = _EVAL_2757 <= _EVAL_3169;
  assign _EVAL_3836 = _EVAL_1649 & _EVAL_3165;
  assign _EVAL_297 = _EVAL_999 & _EVAL_826;
  assign _EVAL_3382 = _EVAL_3562 & _EVAL_3407;
  assign _EVAL_1119 = _EVAL_1649 & _EVAL_2002;
  assign _EVAL_3149 = _EVAL_2809 & _EVAL_2941;
  assign _EVAL_472 = _EVAL_2031 & _EVAL_2047;
  assign _EVAL_3689 = _EVAL_1361[2];
  assign _EVAL_1393 = _EVAL_1560 & _EVAL_1142;
  assign _EVAL_716 = _EVAL_1546 & _EVAL_1004;
  assign _EVAL_3006 = _EVAL_1649 & _EVAL_1444;
  assign _EVAL_2638 = _EVAL_2875 & _EVAL_2941;
  assign _EVAL_2780 = |_EVAL_514;
  assign _EVAL_637 = _EVAL_1246 & _EVAL_701;
  assign _EVAL_2835 = _EVAL_2532 & _EVAL_2538;
  assign _EVAL_2338 = _EVAL_419 & _EVAL_2941;
  assign _EVAL_1676 = _EVAL_1588 & _EVAL_701;
  assign _EVAL_2631 = _EVAL_3774 & _EVAL_3549;
  assign _EVAL_1881 = _EVAL_1649 & _EVAL_1942;
  assign _EVAL_3821 = _EVAL_2038[83];
  assign _EVAL_674 = _EVAL_1927 & _EVAL_3767;
  assign _EVAL_3428 = _EVAL_2038[86];
  assign _EVAL_2609 = _EVAL_3774 & _EVAL_2635;
  assign _EVAL_1889 = _EVAL_2532 & _EVAL_713;
  assign _EVAL_2324 = _EVAL_2532 & _EVAL_671;
  assign _EVAL_1909 = _EVAL_1927 & _EVAL_3369;
  assign _EVAL_3733 = _EVAL_3749 & _EVAL_2026;
  assign _EVAL_173 = _EVAL_1453 & _EVAL_2047;
  assign _EVAL_2831 = _EVAL_1649 & _EVAL_2406;
  assign _EVAL_3755 = _EVAL_2532 & _EVAL_2272;
  assign _EVAL_665 = _EVAL_1649 & _EVAL_844;
  assign _EVAL_2456 = |_EVAL_1836;
  assign _EVAL_724 = _EVAL_2532 & _EVAL_2726;
  assign _EVAL_1615 = _EVAL_2993 & _EVAL_3854;
  assign _EVAL_1240 = _EVAL_1276 & _EVAL_701;
  assign _EVAL_898 = _EVAL_1713 & _EVAL_701;
  assign _EVAL_2464 = _EVAL_2775[1];
  assign _EVAL_2340 = _EVAL_2532 & _EVAL_1667;
  assign _EVAL_479 = _EVAL_1927 & _EVAL_3540;
  assign _EVAL_3406 = _EVAL_1927 & _EVAL_2452;
  assign _EVAL_2110 = _EVAL_3126 & _EVAL_3703;
  assign _EVAL_2578 = _EVAL_3126 & _EVAL_3549;
  assign _EVAL_2603 = _EVAL_3712 & _EVAL_2047;
  assign _EVAL_464 = _EVAL_2038[111];
  assign _EVAL_3351 = _EVAL_3585 & _EVAL_3790;
  assign _EVAL_3838 = _EVAL_173 & _EVAL_2780;
  assign _EVAL_3605 = |_EVAL_1464;
  assign _EVAL_363 = ~_EVAL_2909;
  assign _EVAL_3498 = |_EVAL_2446;
  assign _EVAL_1317 = _EVAL_1649 & _EVAL_2795;
  assign _EVAL_1095 = _EVAL_230 & _EVAL_826;
  assign _EVAL_1275 = |_EVAL_1873;
  assign _EVAL_1427 = _EVAL_1909 & _EVAL_2047;
  assign _EVAL_1775 = _EVAL_2038[130];
  assign _EVAL_2383 = _EVAL_2532 & _EVAL_3818;
  assign _EVAL_881 = _EVAL_1649 & _EVAL_1544;
  assign _EVAL_2630 = _EVAL_3562 & _EVAL_2235;
  assign _EVAL_1545 = _EVAL_1894 & _EVAL_1004;
  assign _EVAL_358 = _EVAL_1704 & _EVAL_701;
  assign _EVAL_3362 = _EVAL_459 & _EVAL_826;
  assign _EVAL_3120 = |_EVAL_3499;
  assign _EVAL_2003 = _EVAL_2532 & _EVAL_243;
  assign _EVAL_2740 = _EVAL_2067 & _EVAL_1004;
  assign _EVAL_2677 = _EVAL_1927 & _EVAL_2947;
  assign _EVAL_1179 = _EVAL_1927 & _EVAL_1635;
  assign _EVAL_199 = _EVAL_1361[25];
  assign _EVAL_928 = _EVAL_173 & _EVAL_2635;
  assign _EVAL_1930 = |_EVAL_1643;
  assign _EVAL_3583 = _EVAL_2532 & _EVAL_2273;
  assign _EVAL_2089 = _EVAL_173 & _EVAL_1730;
  assign _EVAL_1584 = _EVAL_2761 & _EVAL_2941;
  assign _EVAL_1641 = _EVAL_1361[31];
  assign _EVAL_861 = _EVAL_3774 & _EVAL_3498;
  assign _EVAL_1245 = |_EVAL_345;
  assign _EVAL_2042 = _EVAL_2213 & _EVAL_1004;
  assign _EVAL_181 = _EVAL_1649 & _EVAL_3651;
  assign _EVAL_596 = _EVAL_3125 & _EVAL_3272;
  assign _EVAL_829 = _EVAL_1649 & _EVAL_3368;
  assign _EVAL_3320 = _EVAL_1145 & _EVAL_2047;
  assign _EVAL_2776 = _EVAL_1649 & _EVAL_1457;
  assign _EVAL_1919 = _EVAL_2532 & _EVAL_3279;
  assign _EVAL_2364 = _EVAL_1247 & _EVAL_826;
  assign _EVAL_1672 = _EVAL_3774 & _EVAL_1730;
  assign _EVAL_3164 = _EVAL_2532 & _EVAL_1129;
  assign _EVAL_3621 = _EVAL_1858 & _EVAL_2941;
  assign _EVAL_3272 = |_EVAL_3458;
  assign _EVAL_1423 = _EVAL_3125 & _EVAL_3300;
  assign _EVAL_3614 = _EVAL_2713 & _EVAL_701;
  assign _EVAL_769 = _EVAL_3125 & _EVAL_3790;
  assign _EVAL_2151 = _EVAL_3562 & _EVAL_1176;
  assign _EVAL_3258 = _EVAL_2038[107];
  assign _EVAL_3350 = _EVAL_2038[70];
  assign _EVAL_2073 = _EVAL_3774 & _EVAL_1223;
  assign _EVAL_706 = _EVAL_3274 & _EVAL_2047;
  assign _EVAL_578 = _EVAL_2419 & _EVAL_826;
  assign _EVAL_2161 = _EVAL_3554 & _EVAL_826;
  assign _EVAL_2280 = _EVAL_1295 & _EVAL_701;
  assign _EVAL_306 = _EVAL_1649 & _EVAL_1875;
  assign _EVAL_286 = _EVAL_522 & _EVAL_149;
  assign _EVAL_629 = _EVAL_1640 & _EVAL_701;
  assign _EVAL_718 = _EVAL_1927 & _EVAL_2898;
  assign _EVAL_760 = _EVAL_2387 & _EVAL_826;
  assign _EVAL_1648 = _EVAL_2532 & _EVAL_1850;
  assign _EVAL_3458 = _EVAL_2850[26];
  assign _EVAL_764 = _EVAL_3585 & _EVAL_443;
  assign _EVAL_2848 = _EVAL_1927 & _EVAL_2538;
  assign _EVAL_2507 = _EVAL_2532 & _EVAL_3280;
  assign _EVAL_945 = _EVAL_1361[3];
  assign _EVAL_3750 = _EVAL_1927 & _EVAL_3207;
  assign _EVAL_1975 = _EVAL_1069 & _EVAL_1004;
  assign _EVAL_1050 = _EVAL_763 & _EVAL_2941;
  assign _EVAL_1850 = _EVAL_2038[96];
  assign _EVAL_2277 = _EVAL_2532 & _EVAL_399;
  assign _EVAL_1386 = _EVAL_1878 & _EVAL_701;
  assign _EVAL_1874 = _EVAL_883 & _EVAL_2941;
  assign _EVAL_2567 = _EVAL_3144 & _EVAL_1004;
  assign _EVAL_3609 = _EVAL_173 & _EVAL_1470;
  assign _EVAL_1309 = _EVAL_173 & _EVAL_1223;
  assign _EVAL_1804 = _EVAL_2505 & _EVAL_2047;
  assign _EVAL_985 = _EVAL_2038[94];
  assign _EVAL_1078 = _EVAL_3247 & _EVAL_826;
  assign monitor__EVAL_8 = out_back__EVAL_6;
  assign _EVAL_2608 = _EVAL_1361[26];
  assign _EVAL_1403 = _EVAL_1838 & _EVAL_2047;
  assign _EVAL_3009 = _EVAL_2768 & _EVAL_826;
  assign _EVAL_798 = _EVAL_3585 & _EVAL_3252;
  assign _EVAL_433 = _EVAL_3659 & _EVAL_2047;
  assign _EVAL_3377 = _EVAL_1649 & _EVAL_3223;
  assign _EVAL_3789 = _EVAL_1414 & _EVAL_2941;
  assign _EVAL_852 = _EVAL_2104 & _EVAL_2047;
  assign _EVAL_3041 = _EVAL_1927 & _EVAL_475;
  assign _EVAL_1212 = _EVAL_2442 & _EVAL_2047;
  assign _EVAL_1361 = {_EVAL_3780,_EVAL_454,_EVAL_460,_EVAL_194};
  assign _EVAL_3511 = _EVAL_1649 & _EVAL_697;
  assign _EVAL_2829 = _EVAL_2295 & _EVAL_1004;
  assign _EVAL_361 = _EVAL_1927 & _EVAL_2566;
  assign _EVAL_1514 = _EVAL_2532 & _EVAL_1701;
  assign _EVAL_2750 = _EVAL_2993 & _EVAL_1559;
  assign _EVAL_1377 = _EVAL_3125 & _EVAL_443;
  assign _EVAL_1160 = _EVAL_3125 & _EVAL_2456;
  assign _EVAL_1235 = _EVAL_3125 & _EVAL_846;
  assign _EVAL_2679 = _EVAL_1649 & _EVAL_2747;
  assign _EVAL_1559 = |_EVAL_199;
  assign _EVAL_3031 = _EVAL_927 & _EVAL_2941;
  assign _EVAL_2026 = |_EVAL_2914;
  assign _EVAL_418 = _EVAL_155 != 127'h0;
  assign _EVAL_3128 = _EVAL_2775[11];
  assign _EVAL_720 = _EVAL_2038[88];
  assign _EVAL_182 = _EVAL_397 & _EVAL_2235;
  assign _EVAL_2598 = _EVAL_2933 & _EVAL_2047;
  assign _EVAL_216 = _EVAL_2775[10];
  assign _EVAL_2336 = _EVAL_2292 & _EVAL_1004;
  assign _EVAL_3502 = _EVAL_1649 & _EVAL_3696;
  assign _EVAL_971 = _EVAL_3774 & _EVAL_3810;
  assign _EVAL_1462 = _EVAL_3562 & _EVAL_3300;
  assign _EVAL_2611 = _EVAL_983 & _EVAL_2941;
  assign _EVAL_2041 = _EVAL_1649 & _EVAL_3287;
  assign _EVAL_2675 = _EVAL_1649 & _EVAL_1338;
  assign _EVAL_1166 = _EVAL_2729 & _EVAL_826;
  assign _EVAL_3763 = _EVAL_173 & _EVAL_1559;
  assign _EVAL_3046 = _EVAL_2038[43];
  assign _EVAL_3207 = _EVAL_2038[25];
  assign _EVAL_1249 = _EVAL_1965 & _EVAL_701;
  assign _EVAL_3611 = _EVAL_2532 & _EVAL_3540;
  assign _EVAL_3132 = _EVAL_2038[110];
  assign _EVAL_3820 = _EVAL_568 & _EVAL_1004;
  assign _EVAL_2949 = _EVAL_2532 & _EVAL_3293;
  assign _EVAL_2331 = _EVAL_1927 & _EVAL_2187;
  assign _EVAL_2048 = _EVAL_624 & _EVAL_2047;
  assign _EVAL_3669 = _EVAL_1898 & _EVAL_2047;
  assign _EVAL_2786 = _EVAL_556 & _EVAL_1004;
  assign _EVAL_3119 = _EVAL_2850[4];
  assign _EVAL_1573 = _EVAL_2690 & _EVAL_701;
  assign _EVAL_221 = _EVAL_1001 & _EVAL_701;
  assign _EVAL_3543 = _EVAL_3585 & _EVAL_1210;
  assign _EVAL_1261 = _EVAL_2950 & _EVAL_2941;
  assign _EVAL_3487 = _EVAL_2485 & _EVAL_2941;
  assign _EVAL_2610 = _EVAL_915 & _EVAL_1456;
  assign _EVAL_1475 = _EVAL_2038[21];
  assign _EVAL_3813 = _EVAL_2343 & _EVAL_701;
  assign _EVAL_154 = |_EVAL_3805;
  assign _EVAL_3647 = _EVAL_1460 & _EVAL_2047;
  assign _EVAL_2437 = _EVAL_1649 & _EVAL_294;
  assign _EVAL_2291 = _EVAL_2120 & _EVAL_3830;
  assign _EVAL_539 = _EVAL_1927 & _EVAL_2731;
  assign _EVAL_1132 = _EVAL_3125 & _EVAL_3407;
  assign _EVAL_3024 = _EVAL_1412 & _EVAL_2047;
  assign _EVAL_1838 = _EVAL_1927 & _EVAL_1431;
  assign _EVAL_1114 = _EVAL_1927 & _EVAL_1475;
  assign _EVAL_968 = _EVAL_392 & _EVAL_701;
  assign _EVAL_2584 = _EVAL_878 & _EVAL_2047;
  assign _EVAL_768 = _EVAL_2038[87];
  assign _EVAL_2100 = _EVAL_3585 & _EVAL_1245;
  assign _EVAL_2635 = |_EVAL_1356;
  assign _EVAL_1860 = _EVAL_825 & _EVAL_1004;
  assign _EVAL_2390 = _EVAL_173 & _EVAL_1442;
  assign _EVAL_398 = _EVAL_2038[123];
  assign _EVAL_2768 = _EVAL_1649 & _EVAL_1057;
  assign _EVAL_1864 = _EVAL_3739 & _EVAL_701;
  assign _EVAL_577 = _EVAL_1927 & _EVAL_226;
  assign _EVAL_1042 = _EVAL_3778 & _EVAL_701;
  assign _EVAL_1531 = _EVAL_2493 & _EVAL_2941;
  assign _EVAL_405 = |_EVAL_1929;
  assign _EVAL_1642 = _EVAL_2245 & _EVAL_2941;
  assign _EVAL_3853 = _EVAL_2562 & _EVAL_2047;
  assign _EVAL_3088 = _EVAL_3175 & _EVAL_2941;
  assign _EVAL_1668 = _EVAL_3257 & _EVAL_2047;
  assign _EVAL_3594 = _EVAL_3562 & _EVAL_3790;
  assign _EVAL_661 = _EVAL_2126 & _EVAL_2047;
  assign _EVAL_666 = _EVAL_2695 & _EVAL_701;
  assign _EVAL_2821 = _EVAL_2038[102];
  assign _EVAL_1055 = _EVAL_173 & _EVAL_1125;
  assign _EVAL_2673 = _EVAL_3562 & _EVAL_481;
  assign _EVAL_3693 = _EVAL_3774 & _EVAL_1559;
  assign _EVAL_2413 = _EVAL_2532 & _EVAL_457;
  assign _EVAL_283 = _EVAL_929 & _EVAL_701;
  assign _EVAL_1038 = _EVAL_3682 & _EVAL_701;
  assign _EVAL_3728 = _EVAL_1603 & _EVAL_701;
  assign _EVAL_483 = _EVAL_1927 & _EVAL_713;
  assign _EVAL_2564 = _EVAL_1649 & _EVAL_1793;
  assign _EVAL_501 = _EVAL_1927 & _EVAL_950;
  assign _EVAL_3283 = _EVAL_173 & _EVAL_1478;
  assign _EVAL_3602 = _EVAL_430 & _EVAL_2941;
  assign _EVAL_2356 = _EVAL_1983 & _EVAL_2047;
  assign _EVAL_2819 = _EVAL_1298 & _EVAL_1004;
  assign _EVAL_1490 = _EVAL_2433 & _EVAL_701;
  assign _EVAL_3306 = _EVAL_597 & _EVAL_826;
  assign _EVAL_2433 = _EVAL_1690 & _EVAL_2047;
  assign _EVAL_307 = _EVAL_1361[15];
  assign _EVAL_1748 = _EVAL_2993 & _EVAL_417;
  assign _EVAL_1660 = _EVAL_1157 & _EVAL_2047;
  assign _EVAL_766 = _EVAL_2241 & _EVAL_2047;
  assign _EVAL_1025 = _EVAL_3501 & _EVAL_2047;
  assign _EVAL_3551 = _EVAL_1649 & _EVAL_1304;
  assign _EVAL_439 = _EVAL_3126 & _EVAL_2447;
  assign _EVAL_3552 = _EVAL_2045 & _EVAL_1004;
  assign _EVAL_2068 = _EVAL_2794 & _EVAL_507;
  assign _EVAL_3252 = |_EVAL_2721;
  assign _EVAL_2736 = _EVAL_1197 & _EVAL_1004;
  assign _EVAL_2056 = _EVAL_2038[81];
  assign _EVAL_269 = _EVAL_1927 & _EVAL_1665;
  assign _EVAL_349 = _EVAL_1649 & _EVAL_1371;
  assign _EVAL_713 = _EVAL_2038[64];
  assign _EVAL_1137 = _EVAL_728 & _EVAL_2047;
  assign _EVAL_523 = _EVAL_2038[118];
  assign _EVAL_2613 = _EVAL_2532 & _EVAL_720;
  assign _EVAL_2058 = _EVAL_3754 & _EVAL_826;
  assign _EVAL_1029 = _EVAL_2038[66];
  assign _EVAL_3045 = _EVAL_538 & _EVAL_2941;
  assign _EVAL_329 = _EVAL_2038[32];
  assign _EVAL_977 = _EVAL_3544 & _EVAL_701;
  assign _EVAL_2634 = _EVAL_2239 & _EVAL_2047;
  assign _EVAL_1924 = _EVAL_3344 & _EVAL_2047;
  assign _EVAL_1570 = _EVAL_2512 & _EVAL_701;
  assign _EVAL_2353 = _EVAL_1927 & _EVAL_1205;
  assign _EVAL_2260 = _EVAL_1226 & _EVAL_2047;
  assign _EVAL_993 = _EVAL_1214 & _EVAL_2047;
  assign _EVAL_2208 = _EVAL_3459 & _EVAL_701;
  assign _EVAL_2244 = _EVAL_1693 & _EVAL_2047;
  assign _EVAL_3154 = _EVAL_951 & _EVAL_2047;
  assign _EVAL_3026 = _EVAL_1289 & _EVAL_701;
  assign _EVAL_3023 = _EVAL_3562 & _EVAL_1571;
  assign _EVAL_1159 = _EVAL_3253 & _EVAL_2047;
  assign _EVAL_1355 = _EVAL_1927 & _EVAL_2214;
  assign _EVAL_2404 = _EVAL_2243 & _EVAL_2047;
  assign _EVAL_3159 = _EVAL_3126 & _EVAL_405;
  assign _EVAL_2177 = _EVAL_3585 & _EVAL_2261;
  assign _EVAL_1849 = _EVAL_3582 & _EVAL_2047;
  assign _EVAL_2290 = _EVAL_2532 & _EVAL_2176;
  assign _EVAL_1868 = |_EVAL_1807;
  assign _EVAL_3648 = _EVAL_1927 & _EVAL_2718;
  assign _EVAL_3173 = _EVAL_3562 & _EVAL_3649;
  assign _EVAL_1058 = _EVAL_1927 & _EVAL_234;
  assign _EVAL_442 = _EVAL_3774 & _EVAL_2678;
  assign _EVAL_3032 = _EVAL_183 & _EVAL_2941;
  assign _EVAL_915 = _EVAL_2296 & _EVAL_304;
  assign _EVAL_2203 = _EVAL_2437 & _EVAL_826;
  assign _EVAL_2436 = |_EVAL_1945;
  assign _EVAL_1916 = _EVAL_1934 & _EVAL_1004;
  assign _EVAL_598 = _EVAL_2532 & _EVAL_3709;
  assign _EVAL_581 = _EVAL_2532 & _EVAL_1330;
  assign _EVAL_1885 = _EVAL_173 & _EVAL_2335;
  assign _EVAL_2524 = _EVAL_3477 & _EVAL_2047;
  assign _EVAL_2295 = _EVAL_1562 & _EVAL_2047;
  assign _EVAL_553 = _EVAL_2775 & 20'h7f380;
  assign _EVAL_2804 = _EVAL_2839 & _EVAL_2047;
  assign _EVAL_1599 = _EVAL_1294 & _EVAL_2047;
  assign _EVAL_3439 = _EVAL_1917 | _EVAL_1560;
  assign _EVAL_3065 = _EVAL_766 & _EVAL_1004;
  assign _EVAL_1986 = |_EVAL_3226;
  assign _EVAL_3541 = _EVAL_2684 & _EVAL_2026;
  assign _EVAL_3668 = _EVAL_3755 & _EVAL_2047;
  assign _EVAL_1054 = _EVAL_3306 & _EVAL_2941;
  assign _EVAL_1989 = _EVAL_1927 & _EVAL_1887;
  assign _EVAL_1324 = _EVAL_748 & _EVAL_2941;
  assign _EVAL_958 = _EVAL_249 & _EVAL_701;
  assign _EVAL_1943 = _EVAL_1927 & _EVAL_671;
  assign monitor__EVAL_1 = _EVAL_110;
  assign _EVAL_2869 = _EVAL_1649 & _EVAL_1656;
  assign _EVAL_2363 = _EVAL_2564 & _EVAL_826;
  assign _EVAL_332 = _EVAL_1173 & _EVAL_2047;
  assign _EVAL_3501 = _EVAL_1927 & _EVAL_790;
  assign _EVAL_1736 = _EVAL_2532 & _EVAL_3497;
  assign _EVAL_635 = _EVAL_2038[33];
  assign _EVAL_152 = _EVAL_1649 & _EVAL_1852;
  assign _EVAL_3731 = _EVAL_608 & _EVAL_2047;
  assign _EVAL_1028 = _EVAL_2038[51];
  assign _EVAL_2426 = _EVAL_1649 & _EVAL_1532;
  assign _EVAL_1356 = _EVAL_1361[27];
  assign _EVAL_2395 = _EVAL_651[128];
  assign _EVAL_3592 = _EVAL_1897 & _EVAL_802;
  assign _EVAL_484 = _EVAL_881 & _EVAL_826;
  assign _EVAL_1357 = _EVAL_2260 & _EVAL_1004;
  assign _EVAL_1271 = _EVAL_527 & _EVAL_2047;
  assign _EVAL_1708 = |_EVAL_2608;
  assign _EVAL_1136 = _EVAL_316 & _EVAL_701;
  assign _EVAL_1150 = _EVAL_1626 & _EVAL_1004;
  assign _EVAL_233 = _EVAL_2804 & _EVAL_1004;
  assign _EVAL_3196 = _EVAL_1897 & _EVAL_3120;
  assign _EVAL_1818 = _EVAL_711 & _EVAL_701;
  assign _EVAL_608 = _EVAL_1927 & _EVAL_960;
  assign monitor__EVAL_14 = _EVAL_5;
  assign _EVAL_2247 = _EVAL_785 & _EVAL_1811;
  assign _EVAL_671 = _EVAL_2038[57];
  assign _EVAL_1685 = _EVAL_2038[1];
  assign _EVAL_1316 = _EVAL_2038[127];
  assign _EVAL_3822 = _EVAL_1989 & _EVAL_2047;
  assign _EVAL_2973 = _EVAL_785 & _EVAL_481;
  assign _EVAL_2367 = _EVAL_3774 & _EVAL_2541;
  assign _EVAL_891 = _EVAL_3125 & _EVAL_1176;
  assign _EVAL_546 = _EVAL_306 & _EVAL_826;
  assign _EVAL_2857 = _EVAL_1649 & _EVAL_1086;
  assign _EVAL_291 = _EVAL_773 & _EVAL_1004;
  assign _EVAL_1551 = |_EVAL_1646;
  assign _EVAL_2972 = _EVAL_1649 & _EVAL_3701;
  assign _EVAL_1079 = _EVAL_2813 & _EVAL_701;
  assign _EVAL_3212 = _EVAL_3126 & _EVAL_2487;
  assign _EVAL_251 = _EVAL_1508 & _EVAL_2047;
  assign _EVAL_1233 = _EVAL_1361[23];
  assign _EVAL_3727 = _EVAL_2319 & _EVAL_2047;
  assign _EVAL_3257 = _EVAL_1927 & _EVAL_3293;
  assign _EVAL_3659 = _EVAL_1927 & _EVAL_3405;
  assign _EVAL_3180 = _EVAL_397 & _EVAL_1571;
  assign _EVAL_663 = _EVAL_2507 & _EVAL_2047;
  assign _EVAL_599 = _EVAL_2470 & _EVAL_701;
  assign _EVAL_2931 = _EVAL_1599 & _EVAL_1004;
  assign _EVAL_3517 = _EVAL_1515 & _EVAL_701;
  assign _EVAL_1445 = _EVAL_2063 & _EVAL_2941;
  assign _EVAL_2368 = _EVAL_2108 & _EVAL_2941;
  assign _EVAL_1746 = _EVAL_2645 & _EVAL_701;
  assign _EVAL_1258 = _EVAL_2458 & _EVAL_826;
  assign _EVAL_920 = _EVAL_879 & _EVAL_2047;
  assign _EVAL_3125 = _EVAL_2776 & _EVAL_826;
  assign _EVAL_1176 = |_EVAL_3119;
  assign _EVAL_2924 = _EVAL_1927 & _EVAL_2118;
  assign _EVAL_1460 = _EVAL_2532 & _EVAL_2821;
  assign _EVAL_1194 = _EVAL_3103 & _EVAL_2047;
  assign _EVAL_239 = _EVAL_3125 & _EVAL_1571;
  assign _EVAL_1276 = _EVAL_998 & _EVAL_2047;
  assign _EVAL_1123 = _EVAL_1649 & _EVAL_3717;
  assign _EVAL_3254 = _EVAL_1291 & _EVAL_826;
  assign _EVAL_2052 = _EVAL_1360 & _EVAL_1004;
  assign _EVAL_1609 = _EVAL_397 & _EVAL_2033;
  assign _EVAL_888 = _EVAL_2993 & _EVAL_1442;
  assign _EVAL_312 = _EVAL_812 & _EVAL_1004;
  assign _EVAL_147 = _EVAL_2675 & _EVAL_826;
  assign _EVAL_246 = _EVAL_2532 & _EVAL_3710;
  assign _EVAL_2691 = _EVAL_2038[129];
  assign _EVAL_2826 = _EVAL_2038[15];
  assign _EVAL_1831 = _EVAL_3562 & _EVAL_1177;
  assign _EVAL_264 = _EVAL_397 & _EVAL_3224;
  assign _EVAL_843 = _EVAL_298 & _EVAL_2047;
  assign _EVAL_3536 = _EVAL_3493 & _EVAL_2047;
  assign _EVAL_436 = &_EVAL_1361;
  assign _EVAL_454 = _EVAL_2111 ? 8'hff : 8'h0;
  assign _EVAL_3048 = _EVAL_3125 & _EVAL_2235;
  assign _EVAL_3739 = _EVAL_3400 & _EVAL_2047;
  assign _EVAL_457 = _EVAL_2038[3];
  assign _EVAL_3028 = _EVAL_3126 & _EVAL_417;
  assign _EVAL_1256 = _EVAL_920 & _EVAL_3854;
  assign _EVAL_1744 = _EVAL_2355 & _EVAL_1004;
  assign _EVAL_2189 = _EVAL_2993 & _EVAL_1708;
  assign _EVAL_976 = _EVAL_1649 & _EVAL_340;
  assign _EVAL_704 = _EVAL_397 & _EVAL_2908;
  assign _EVAL_2468 = |_EVAL_2115;
  assign _EVAL_514 = _EVAL_1361[21];
  assign _EVAL_1246 = _EVAL_2340 & _EVAL_2047;
  assign _EVAL_1883 = _EVAL_1649 & _EVAL_794;
  assign _EVAL_1409 = _EVAL_3126 & _EVAL_370;
  assign _EVAL_2504 = _EVAL_277 & _EVAL_3827;
  assign _EVAL_563 = _EVAL_173 & _EVAL_2447;
  assign _EVAL_1501 = _EVAL_1649 & _EVAL_640;
  assign _EVAL_816 = _EVAL_1668 & _EVAL_1004;
  assign _EVAL_1322 = _EVAL_1302 & _EVAL_826;
  assign _EVAL_1713 = _EVAL_1558 & _EVAL_2047;
  assign _EVAL_3227 = _EVAL_1533 & _EVAL_701;
  assign _EVAL_1800 = _EVAL_2532 & _EVAL_523;
  assign _EVAL_2141 = _EVAL_2993 & _EVAL_1551;
  assign _EVAL_2590 = _EVAL_920 & _EVAL_2468;
  assign _EVAL_2762 = _EVAL_3024 & _EVAL_701;
  assign _EVAL_1353 = _EVAL_477 & _EVAL_1004;
  assign _EVAL_2387 = _EVAL_1649 & _EVAL_3637;
  assign _EVAL_2323 = _EVAL_1649 & _EVAL_184;
  assign _EVAL_1097 = _EVAL_1844 & _EVAL_2941;
  assign _EVAL_3661 = _EVAL_2681 & _EVAL_2047;
  assign _EVAL_2825 = _EVAL_1859 & _EVAL_701;
  assign _EVAL_380 = _EVAL_2850[17];
  assign _EVAL_3110 = _EVAL_248 & _EVAL_2047;
  assign _EVAL_2307 = _EVAL_3585 & _EVAL_3649;
  assign _EVAL_2941 = |_EVAL_2084;
  assign _EVAL_2652 = _EVAL_1083 & _EVAL_2047;
  assign _EVAL_2891 = _EVAL_1649 & _EVAL_2234;
  assign _EVAL_2683 = _EVAL_2065 & _EVAL_1004;
  assign _EVAL_1352 = _EVAL_2570 & _EVAL_2941;
  assign _EVAL_1983 = _EVAL_2532 & _EVAL_2754;
  assign _EVAL_3451 = _EVAL_2995 & _EVAL_826;
  assign _EVAL_2595 = _EVAL_2532 & _EVAL_3421;
  assign _EVAL_2496 = _EVAL_1649 & _EVAL_213;
  assign _EVAL_2138 = _EVAL_1649 & _EVAL_1170;
  assign _EVAL_3235 = _EVAL_1927 & _EVAL_650;
  assign _EVAL_1421 = _EVAL_1649 & _EVAL_1396;
  assign _EVAL_1959 = _EVAL_2532 & _EVAL_960;
  assign _EVAL_2388 = _EVAL_656 & _EVAL_2047;
  assign _EVAL_1820 = _EVAL_664 & _EVAL_1004;
  assign _EVAL_3187 = _EVAL_1361[31:3];
  assign _EVAL_2704 = _EVAL_539 & _EVAL_2047;
  assign _EVAL_3049 = _EVAL_1660 & _EVAL_1004;
  assign _EVAL_1511 = _EVAL_2532 & _EVAL_985;
  assign _EVAL_1098 = _EVAL_3768 & _EVAL_2941;
  assign _EVAL_392 = _EVAL_2796 & _EVAL_2047;
  assign _EVAL_2501 = _EVAL_397 & _EVAL_942;
  assign _EVAL_3232 = |_EVAL_3118;
  assign _EVAL_2735 = _EVAL_2850[1];
  assign _EVAL_3784 = _EVAL_774 & _EVAL_2941;
  assign _EVAL_883 = _EVAL_2471 & _EVAL_826;
  assign _EVAL_1013 = _EVAL_3585 & _EVAL_846;
  assign _EVAL_407 = _EVAL_2288 & _EVAL_1004;
  assign _EVAL_1699 = _EVAL_675 & _EVAL_2941;
  assign _EVAL_1436 = &_EVAL_2115;
  assign _EVAL_2808 = _EVAL_1649 & _EVAL_709;
  assign _EVAL_1169 = _EVAL_1927 & _EVAL_2255;
  assign _EVAL_680 = _EVAL_3585 & _EVAL_1177;
  assign _EVAL_833 = _EVAL_277 & _EVAL_3087;
  assign _EVAL_698 = _EVAL_2038[101];
  assign _EVAL_2550 = _EVAL_2038[513];
  assign _EVAL_1984 = _EVAL_2013 & _EVAL_2047;
  assign _EVAL_1686 = _EVAL_1404 & _EVAL_701;
  assign _EVAL_3799 = _EVAL_169 & _EVAL_1004;
  assign _EVAL_1922 = _EVAL_397 & _EVAL_1210;
  assign _EVAL_1454 = _EVAL_1649 & _EVAL_3211;
  assign _EVAL_3713 = _EVAL_3125 & _EVAL_3761;
  assign _EVAL_1693 = _EVAL_2532 & _EVAL_2898;
  assign _EVAL_919 = _EVAL_2850[30];
  assign _EVAL_3553 = _EVAL_3562 & _EVAL_942;
  assign _EVAL_2376 = _EVAL_3360 & _EVAL_2047;
  assign _EVAL_1414 = _EVAL_1242 & _EVAL_826;
  assign _EVAL_3289 = _EVAL_2038[105];
  assign _EVAL_1577 = _EVAL_2579 & _EVAL_2047;
  assign _EVAL_1837 = _EVAL_2524 & _EVAL_1004;
  assign _EVAL_163 = _EVAL_1649 & _EVAL_3435;
  assign _EVAL_3703 = |_EVAL_2955;
  assign _EVAL_2858 = _EVAL_3674 & _EVAL_2941;
  assign _EVAL_3655 = _EVAL_1927 & _EVAL_1650;
  assign _EVAL_2588 = _EVAL_3585 & _EVAL_1111;
  assign _EVAL_1018 = _EVAL_2324 & _EVAL_2047;
  assign _EVAL_1556 = _EVAL_2209 & _EVAL_826;
  assign _EVAL_2269 = _EVAL_1300 & _EVAL_1004;
  assign _EVAL_3325 = _EVAL_1465 & _EVAL_1004;
  assign _EVAL_1494 = _EVAL_2823 & _EVAL_1004;
  assign _EVAL_3769 = _EVAL_1927 & _EVAL_243;
  assign _EVAL_572 = _EVAL_3766 & _EVAL_2941;
  assign _EVAL_3352 = _EVAL_1927 & _EVAL_511;
  assign _EVAL_1807 = _EVAL_1361[20];
  assign _EVAL_376 = _EVAL_1192 & _EVAL_2047;
  assign _EVAL_2713 = _EVAL_724 & _EVAL_2047;
  assign _EVAL_1719 = _EVAL_1219 & _EVAL_2941;
  assign _EVAL_929 = _EVAL_2606 & _EVAL_2047;
  assign _EVAL_2319 = _EVAL_2532 & _EVAL_3289;
  assign _EVAL_633 = _EVAL_2136 & _EVAL_1004;
  assign _EVAL_1141 = _EVAL_2775[19];
  assign _EVAL_1228 = _EVAL_3125 & _EVAL_2033;
  assign _EVAL_3805 = _EVAL_1361[15:8];
  assign _EVAL_3308 = _EVAL_2038[13];
  assign _EVAL_2402 = _EVAL_785 & _EVAL_3827;
  assign _EVAL_1399 = _EVAL_3536 & _EVAL_701;
  assign _EVAL_191 = _EVAL_3125 & _EVAL_1210;
  assign _EVAL_3294 = _EVAL_729 & _EVAL_2047;
  assign _EVAL_2552 = _EVAL_3215 & _EVAL_826;
  assign _EVAL_1704 = _EVAL_897 & _EVAL_2047;
  assign _EVAL_1227 = _EVAL_3389 & _EVAL_1004;
  assign _EVAL_2180 = _EVAL_2200 & _EVAL_1004;
  assign _EVAL_1001 = _EVAL_1891 & _EVAL_2047;
  assign _EVAL_3665 = _EVAL_173 & _EVAL_3549;
  assign _EVAL_303 = _EVAL_1862 & _EVAL_2047;
  assign _EVAL_1388 = _EVAL_836 & _EVAL_2941;
  assign _EVAL_3492 = _EVAL_1649 & _EVAL_3619;
  assign _EVAL_2882 = _EVAL_2708 & _EVAL_2941;
  assign _EVAL_998 = _EVAL_2532 & _EVAL_1635;
  assign _EVAL_252 = _EVAL_2794 & _EVAL_2941;
  assign _EVAL_1465 = _EVAL_400 & _EVAL_2047;
  assign _EVAL_2582 = _EVAL_2581 & _EVAL_701;
  assign _EVAL_565 = _EVAL_2679 & _EVAL_826;
  assign _EVAL_1861 = _EVAL_2993 & _EVAL_1583;
  assign _EVAL_839 = _EVAL_1881 & _EVAL_826;
  assign _EVAL_3146 = _EVAL_388 & _EVAL_701;
  assign _EVAL_357 = _EVAL_1649 & _EVAL_1780;
  assign _EVAL_2185 = _EVAL_2038[100];
  assign _EVAL_1405 = _EVAL_3671 & _EVAL_2047;
  assign _EVAL_1561 = _EVAL_2532 & _EVAL_3046;
  assign _EVAL_1691 = _EVAL_3774 & _EVAL_2487;
  assign _EVAL_1626 = _EVAL_3655 & _EVAL_2047;
  assign _EVAL_2562 = _EVAL_2532 & _EVAL_3792;
  assign _EVAL_1003 = _EVAL_1361[8];
  assign _EVAL_3057 = _EVAL_2038[56];
  assign _EVAL_2688 = _EVAL_2993 & _EVAL_3703;
  assign _EVAL_3641 = _EVAL_173 & _EVAL_1708;
  assign _EVAL_1302 = _EVAL_1649 & _EVAL_515;
  assign _EVAL_742 = _EVAL_3506 & _EVAL_826;
  assign _EVAL_3280 = _EVAL_2038[75];
  assign _EVAL_1478 = |_EVAL_945;
  assign _EVAL_502 = _EVAL_1432 & _EVAL_2047;
  assign _EVAL_1819 = _EVAL_2532 & _EVAL_234;
  assign _EVAL_2769 = _EVAL_1927 & _EVAL_3365;
  assign _EVAL_714 = _EVAL_2652 & _EVAL_701;
  assign _EVAL_3617 = _EVAL_3116 & _EVAL_701;
  assign _EVAL_2213 = _EVAL_3297 & _EVAL_2047;
  assign _EVAL_3432 = _EVAL_1649 & _EVAL_2874;
  assign _EVAL_2411 = _EVAL_2038[39];
  assign _EVAL_1284 = _EVAL_2029 & _EVAL_2047;
  assign _EVAL_2001 = _EVAL_173 & _EVAL_1551;
  assign _EVAL_1442 = |_EVAL_807;
  assign _EVAL_372 = _EVAL_1259 & _EVAL_2941;
  assign _EVAL_3229 = _EVAL_2039 & _EVAL_701;
  assign _EVAL_1767 = _EVAL_1883 & _EVAL_826;
  assign _EVAL_1663 = _EVAL_1525 & _EVAL_1004;
  assign _EVAL_1402 = _EVAL_2552 & _EVAL_2941;
  assign _EVAL_218 = _EVAL_3126 & _EVAL_1442;
  assign _EVAL_580 = _EVAL_2993 & _EVAL_3810;
  assign _EVAL_1784 = _EVAL_2532 & _EVAL_1236;
  assign _EVAL_3192 = _EVAL_3320 & _EVAL_701;
  assign _EVAL_2976 = _EVAL_2092 & _EVAL_701;
  assign _EVAL_2241 = _EVAL_1927 & _EVAL_2272;
  assign _EVAL_3281 = _EVAL_1194 & _EVAL_1004;
  assign _EVAL_2703 = _EVAL_1649 & _EVAL_2623;
  assign _EVAL_3379 = _EVAL_3562 & _EVAL_2033;
  assign _EVAL_1502 = _EVAL_3126 & _EVAL_1868;
  assign _EVAL_1862 = _EVAL_2532 & _EVAL_1598;
  assign _EVAL_2232 = _EVAL_3585 & _EVAL_2235;
  assign _EVAL_3687 = _EVAL_2775[6];
  assign _EVAL_541 = _EVAL_2146 & _EVAL_701;
  assign _EVAL_3649 = |_EVAL_3550;
  assign _EVAL_2760 = _EVAL_1511 & _EVAL_2047;
  assign _EVAL_1372 = _EVAL_1846 & _EVAL_2047;
  assign _EVAL_1999 = _EVAL_2532 & _EVAL_659;
  assign _EVAL_1394 = _EVAL_3675 & _EVAL_701;
  assign _EVAL_268 = _EVAL_2532 & _EVAL_3428;
  assign _EVAL_2372 = _EVAL_3585 & _EVAL_1571;
  assign _EVAL_1667 = _EVAL_2038[73];
  assign _EVAL_512 = _EVAL_2532 & _EVAL_398;
  assign _EVAL_1113 = ~_EVAL_3846;
  assign _EVAL_3297 = _EVAL_1927 & _EVAL_3158;
  assign _EVAL_3419 = _EVAL_2516 & _EVAL_1004;
  assign _EVAL_2457 = _EVAL_1585 & _EVAL_701;
  assign _EVAL_1709 = _EVAL_1078 & _EVAL_2941;
  assign _EVAL_1201 = _EVAL_1649 & _EVAL_3036;
  assign _EVAL_814 = _EVAL_3565 & _EVAL_2941;
  assign _EVAL_2096 = |_EVAL_424;
  assign _EVAL_3190 = _EVAL_1612 & _EVAL_2941;
  assign _EVAL_1552 = _EVAL_2648 & _EVAL_2941;
  assign _EVAL_2481 = _EVAL_3736 & _EVAL_2047;
  assign _EVAL_1075 = _EVAL_1189 & _EVAL_1004;
  assign _EVAL_3085 = _EVAL_1361[28];
  assign _EVAL_1115 = _EVAL_2532 & _EVAL_3767;
  assign _EVAL_1213 = _EVAL_1405 & _EVAL_1429;
  assign _EVAL_377 = _EVAL_1984 & _EVAL_701;
  assign _EVAL_2146 = _EVAL_1893 & _EVAL_2047;
  assign _EVAL_1083 = _EVAL_2532 & _EVAL_2718;
  assign _EVAL_1939 = _EVAL_1979 & _EVAL_1004;
  assign _EVAL_3556 = _EVAL_2532 & _EVAL_2643;
  assign _EVAL_940 = _EVAL_2613 & _EVAL_2047;
  assign _EVAL_2864 = _EVAL_694 & _EVAL_701;
  assign _EVAL_3826 = _EVAL_1649 & _EVAL_338;
  assign _EVAL_1825 = _EVAL_375 & _EVAL_2941;
  assign _EVAL_1806 = _EVAL_2532 & _EVAL_2550;
  assign _EVAL_3052 = _EVAL_397 & _EVAL_2162;
  assign _EVAL_1724 = _EVAL_472 & _EVAL_1004;
  assign _EVAL_740 = _EVAL_2394 & _EVAL_2047;
  assign _EVAL_183 = _EVAL_3006 & _EVAL_826;
  assign _EVAL_3578 = _EVAL_2532 & _EVAL_549;
  assign _EVAL_3697 = _EVAL_2706 & _EVAL_2047;
  assign _EVAL_1453 = _EVAL_1927 & _EVAL_2548;
  assign _EVAL_3139 = _EVAL_3562 & _EVAL_2261;
  assign _EVAL_725 = _EVAL_3126 & _EVAL_1986;
  assign _EVAL_1363 = _EVAL_1405 & _EVAL_3830;
  assign _EVAL_561 = _EVAL_1461 & _EVAL_2941;
  assign _EVAL_1863 = _EVAL_3126 & _EVAL_2335;
  assign _EVAL_824 = _EVAL_2850[11];
  assign _EVAL_217 = _EVAL_976 & _EVAL_826;
  assign _EVAL_1782 = _EVAL_2356 & _EVAL_1436;
  assign _EVAL_3021 = _EVAL_2532 & _EVAL_3057;
  assign _EVAL_2355 = _EVAL_2331 & _EVAL_2047;
  assign _EVAL_3253 = _EVAL_1927 & _EVAL_3808;
  assign _EVAL_1589 = _EVAL_1649 & _EVAL_1053;
  assign _EVAL_2374 = _EVAL_2923 & _EVAL_2941;
  assign _EVAL_2105 = _EVAL_3385 & _EVAL_2047;
  assign _EVAL_2669 = _EVAL_1927 & _EVAL_1701;
  assign _EVAL_2599 = _EVAL_1123 & _EVAL_826;
  assign _EVAL_3628 = _EVAL_2532 & _EVAL_2214;
  assign _EVAL_2238 = _EVAL_1351 & _EVAL_2047;
  assign _EVAL_2435 = _EVAL_1921 & _EVAL_701;
  assign _EVAL_3515 = _EVAL_397 & _EVAL_443;
  assign _EVAL_3574 = _EVAL_2723 & _EVAL_701;
  assign _EVAL_1387 = _EVAL_578 & _EVAL_2941;
  assign _EVAL_2334 = _EVAL_3362 & _EVAL_2941;
  assign _EVAL_730 = _EVAL_1427 & _EVAL_731;
  assign _EVAL_1747 = _EVAL_882 & _EVAL_3605;
  assign _EVAL_2641 = _EVAL_1600 & _EVAL_2047;
  assign _EVAL_2067 = _EVAL_1260 & _EVAL_2047;
  assign _EVAL_2836 = _EVAL_1927 & _EVAL_2726;
  assign _EVAL_1297 = _EVAL_2993 & _EVAL_1470;
  assign _EVAL_3495 = _EVAL_1632 & _EVAL_2047;
  assign _EVAL_316 = _EVAL_1162 & _EVAL_2047;
  assign _EVAL_1006 = _EVAL_2850[19];
  assign _EVAL_352 = _EVAL_1649 & _EVAL_3806;
  assign _EVAL_2605 = _EVAL_2383 & _EVAL_2047;
  assign _EVAL_1817 = _EVAL_3562 & _EVAL_1210;
  assign _EVAL_3712 = _EVAL_1927 & _EVAL_3497;
  assign _EVAL_2666 = _EVAL_3585 & _EVAL_2033;
  assign _EVAL_3749 = _EVAL_3551 & _EVAL_826;
  assign _EVAL_2360 = _EVAL_157 & _EVAL_1004;
  assign _EVAL_310 = _EVAL_1649 & _EVAL_1135;
  assign _EVAL_2579 = _EVAL_1927 & _EVAL_201;
  assign _EVAL_1753 = _EVAL_1290 & _EVAL_1004;
  assign _EVAL_822 = _EVAL_2286 & _EVAL_1004;
  assign _EVAL_3705 = _EVAL_3748 & _EVAL_2047;
  assign _EVAL_1650 = _EVAL_2038[113];
  assign _EVAL_3691 = _EVAL_3650 & _EVAL_826;
  assign _EVAL_2310 = _EVAL_900 & _EVAL_2941;
  assign _EVAL_2636 = _EVAL_757 & _EVAL_701;
  assign _EVAL_424 = _EVAL_1361[24];
  assign _EVAL_3768 = _EVAL_2339 & _EVAL_826;
  assign _EVAL_1362 = _EVAL_173 & _EVAL_2487;
  assign _EVAL_1091 = _EVAL_1927 & _EVAL_1850;
  assign _EVAL_3776 = _EVAL_2123 - 1'h1;
  assign _EVAL_397 = _EVAL_2869 & _EVAL_826;
  assign _EVAL_686 = _EVAL_1649 & _EVAL_2168;
  assign _EVAL_1186 = _EVAL_745 & _EVAL_2047;
  assign _EVAL_922 = _EVAL_3110 & _EVAL_701;
  assign _EVAL_3650 = _EVAL_1649 & _EVAL_1066;
  assign _EVAL_2330 = _EVAL_3705 & _EVAL_1004;
  assign _EVAL_3497 = _EVAL_2038[78];
  assign _EVAL_731 = |_EVAL_3187;
  assign _EVAL_3765 = _EVAL_2038[28];
  assign _EVAL_465 = _EVAL_1373 & _EVAL_2941;
  assign _EVAL_1161 = _EVAL_3301 & _EVAL_1004;
  assign _EVAL_1431 = _EVAL_2038[2];
  assign _EVAL_562 = _EVAL_1927 & _EVAL_659;
  assign _EVAL_3121 = _EVAL_2684 & _EVAL_3827;
  assign _EVAL_3631 = _EVAL_2038[115];
  assign _EVAL_1566 = _EVAL_2038[103];
  assign _EVAL_2886 = _EVAL_2840 & _EVAL_2941;
  assign _EVAL_2343 = _EVAL_2783 & _EVAL_2047;
  assign _EVAL_319 = _EVAL_3691 & _EVAL_2941;
  assign _EVAL_2901 = _EVAL_2771 & _EVAL_2047;
  assign _EVAL_229 = _EVAL_2532 & _EVAL_3207;
  assign _EVAL_611 = _EVAL_3585 & _EVAL_3300;
  assign _EVAL_2031 = _EVAL_1927 & _EVAL_3709;
  assign _EVAL_728 = _EVAL_2532 & _EVAL_3369;
  assign _EVAL_1326 = _EVAL_1403 & _EVAL_1004;
  assign _EVAL_2687 = _EVAL_1649 & _EVAL_1712;
  assign _EVAL_1836 = _EVAL_2850[20];
  assign _EVAL_2111 = _EVAL_84[2];
  assign _EVAL_1717 = _EVAL_1927 & _EVAL_3060;
  assign _EVAL_388 = _EVAL_1463 & _EVAL_2047;
  assign _EVAL_3163 = _EVAL_3125 & _EVAL_914;
  assign _EVAL_1759 = _EVAL_2993 & _EVAL_1478;
  assign _EVAL_2000 = _EVAL_1159 & _EVAL_3120;
  assign _EVAL_620 = _EVAL_3585 & _EVAL_1176;
  assign _EVAL_1898 = _EVAL_2532 & _EVAL_3630;
  assign _EVAL_1811 = |_EVAL_3038;
  assign _EVAL_984 = _EVAL_3239 & _EVAL_701;
  assign _EVAL_2365 = _EVAL_3511 & _EVAL_826;
  assign _EVAL_3181 = _EVAL_3125 & _EVAL_3224;
  assign _EVAL_1519 = _EVAL_1927 & _EVAL_399;
  assign _EVAL_3060 = _EVAL_2038[9];
  assign _EVAL_3042 = _EVAL_3583 & _EVAL_2047;
  assign _EVAL_3503 = _EVAL_1649 & _EVAL_1505;
  assign _EVAL_2824 = _EVAL_2591 & _EVAL_1004;
  assign _EVAL_2045 = _EVAL_577 & _EVAL_2047;
  assign _EVAL_3721 = _EVAL_1959 & _EVAL_2047;
  assign _EVAL_2714 = _EVAL_2775[4];
  assign _EVAL_2014 = _EVAL_1455 & _EVAL_2047;
  assign _EVAL_2500 = _EVAL_1179 & _EVAL_2047;
  assign _EVAL_3087 = |_EVAL_469;
  assign monitor__EVAL_3 = {{2'd0}, _EVAL_367};
  assign _EVAL_574 = _EVAL_2038[108];
  assign _EVAL_3699 = _EVAL_2529 & _EVAL_2941;
  assign _EVAL_941 = _EVAL_3188 & _EVAL_2941;
  assign _EVAL_2237 = _EVAL_2843 & _EVAL_2941;
  assign _EVAL_406 = _EVAL_1577 & _EVAL_1004;
  assign _EVAL_1226 = _EVAL_1927 & _EVAL_3698;
  assign _EVAL_3507 = _EVAL_2532 & _EVAL_1721;
  assign _EVAL_1993 = _EVAL_806 & _EVAL_2047;
  assign _EVAL_2771 = _EVAL_2532 & _EVAL_2407;
  assign _EVAL_2117 = _EVAL_2256 & _EVAL_1004;
  assign _EVAL_2092 = _EVAL_3021 & _EVAL_2047;
  assign _EVAL_315 = _EVAL_2850[3];
  assign _EVAL_1312 = _EVAL_163 & _EVAL_826;
  assign _EVAL_2851 = _EVAL_2634 & _EVAL_701;
  assign monitor__EVAL_0 = _EVAL_9;
  assign _EVAL_1149 = _EVAL_674 & _EVAL_2047;
  assign _EVAL_3604 = _EVAL_2532 & _EVAL_2223;
  assign _EVAL_3389 = _EVAL_1590 & _EVAL_2047;
  assign monitor__EVAL_13 = _EVAL_84;
  assign _EVAL_737 = _EVAL_397 & _EVAL_1930;
  assign _EVAL_2107 = _EVAL_332 & _EVAL_701;
  assign _EVAL_557 = _EVAL_1649 & _EVAL_903;
  assign _EVAL_1100 = _EVAL_173 & _EVAL_1583;
  assign _EVAL_2923 = _EVAL_3796 & _EVAL_826;
  assign _EVAL_3829 = _EVAL_2870 & _EVAL_2047;
  assign _EVAL_1277 = _EVAL_448 & _EVAL_2047;
  assign _EVAL_1728 = _EVAL_3816 & _EVAL_701;
  assign _EVAL_2246 = _EVAL_397 & _EVAL_3252;
  assign _EVAL_2267 = _EVAL_3125 & _EVAL_2194;
  assign _EVAL_1437 = _EVAL_2532 & _EVAL_790;
  assign _EVAL_3518 = _EVAL_1493 & _EVAL_701;
  assign _EVAL_249 = _EVAL_1514 & _EVAL_2047;
  assign _EVAL_2176 = _EVAL_2038[77];
  assign _EVAL_2287 = _EVAL_1927 & _EVAL_3428;
  assign _EVAL_2508 = _EVAL_2775[5];
  assign _EVAL_201 = _EVAL_2038[41];
  assign _EVAL_2139 = _EVAL_181 & _EVAL_826;
  assign _EVAL_2271 = _EVAL_3661 & _EVAL_1004;
  assign _EVAL_2993 = _EVAL_564 & _EVAL_2047;
  assign _EVAL_1671 = _EVAL_1106 & _EVAL_826;
  assign _EVAL_2643 = _EVAL_2038[45];
  assign _EVAL_2040 = _EVAL_397 & _EVAL_1275;
  assign _EVAL_226 = _EVAL_2038[74];
  assign _EVAL_2866 = _EVAL_3668 & _EVAL_701;
  assign _EVAL_1682 = _EVAL_2163 & _EVAL_2047;
  assign _EVAL_3070 = _EVAL_3585 & _EVAL_2908;
  assign _EVAL_1795 = _EVAL_1649 & _EVAL_1644;
  assign _EVAL_2551 = _EVAL_3731 & _EVAL_1004;
  assign _EVAL_2156 = _EVAL_1806 & _EVAL_2047;
  assign _EVAL_681 = _EVAL_3273 & _EVAL_2941;
  assign _EVAL_453 = _EVAL_2912 & _EVAL_1004;
  assign _EVAL_230 = _EVAL_1649 & _EVAL_3414;
  assign _EVAL_1546 = _EVAL_2709 & _EVAL_2047;
  assign _EVAL_2875 = _EVAL_3492 & _EVAL_826;
  assign _EVAL_882 = _EVAL_269 & _EVAL_2047;
  assign _EVAL_1730 = |_EVAL_1725;
  assign _EVAL_3688 = _EVAL_1927 & _EVAL_3821;
  assign _EVAL_2796 = _EVAL_2532 & _EVAL_3350;
  assign _EVAL_2823 = _EVAL_1941 & _EVAL_2047;
  assign _EVAL_2332 = ~_EVAL_1931;
  assign _EVAL_2212 = _EVAL_562 & _EVAL_2047;
  assign _EVAL_2359 = _EVAL_2038[20];
  assign _EVAL_650 = _EVAL_2038[120];
  assign _EVAL_3827 = |_EVAL_1016;
  assign _EVAL_1940 = _EVAL_2532 & _EVAL_3158;
  assign _EVAL_3854 = |_EVAL_2158;
  assign _EVAL_346 = _EVAL_2519 & _EVAL_1004;
  assign _EVAL_1640 = _EVAL_1437 & _EVAL_2047;
  assign _EVAL_1139 = _EVAL_1927 & _EVAL_2317;
  assign _EVAL_370 = |_EVAL_2166;
  assign _EVAL_1007 = _EVAL_3126 & _EVAL_1559;
  assign _EVAL_522 = _EVAL_261 & _EVAL_2047;
  assign _EVAL_3175 = _EVAL_3836 & _EVAL_826;
  assign _EVAL_3050 = _EVAL_1649 & _EVAL_2733;
  assign _EVAL_2940 = _EVAL_1649 & _EVAL_3588;
  assign _EVAL_1735 = _EVAL_2993 & _EVAL_2024;
  assign _EVAL_781 = _EVAL_2532 & _EVAL_204;
  assign _EVAL_831 = _EVAL_2806 & _EVAL_1004;
  assign _EVAL_786 = _EVAL_2993 & _EVAL_2447;
  assign _EVAL_2301 = _EVAL_2038[47];
  assign _EVAL_875 = _EVAL_1649 & _EVAL_1311;
  assign _EVAL_174 = _EVAL_3611 & _EVAL_2047;
  assign monitor__EVAL_12 = _EVAL_119;
  assign _EVAL_2024 = |_EVAL_1523;
  assign _EVAL_393 = _EVAL_3773 & _EVAL_2941;
  assign _EVAL_1077 = _EVAL_1027 & _EVAL_826;
  assign _EVAL_1929 = _EVAL_1361[12];
  assign _EVAL_491 = _EVAL_1649 & _EVAL_1956;
  assign _EVAL_192 = _EVAL_555 & _EVAL_2941;
  assign _EVAL_664 = _EVAL_1169 & _EVAL_2047;
  assign _EVAL_2648 = _EVAL_3292 & _EVAL_826;
  assign _EVAL_1934 = _EVAL_535 & _EVAL_2047;
  assign _EVAL_3547 = _EVAL_2481 & _EVAL_1004;
  assign _EVAL_2912 = _EVAL_401 & _EVAL_2047;
  assign _EVAL_2223 = _EVAL_2038[124];
  assign _EVAL_2843 = _EVAL_2037 & _EVAL_826;
  assign _EVAL_1165 = _EVAL_1910 & _EVAL_2047;
  assign _EVAL_2278 = _EVAL_3125 & _EVAL_3764;
  assign _EVAL_1070 = _EVAL_2850[0];
  assign _EVAL_2867 = _EVAL_2905 & _EVAL_2047;
  assign _EVAL_1474 = _EVAL_1649 & _EVAL_1094;
  assign _EVAL_2516 = _EVAL_788 & _EVAL_2047;
  assign _EVAL_200 = _EVAL_2848 & _EVAL_2047;
  assign _EVAL_649 = _EVAL_1312 & _EVAL_2941;
  assign _EVAL_1069 = _EVAL_255 & _EVAL_2047;
  assign _EVAL_1530 = _EVAL_3411 & _EVAL_701;
  assign _EVAL_1019 = _EVAL_2760 & _EVAL_701;
  assign _EVAL_1045 = _EVAL_1139 & _EVAL_2047;
  assign _EVAL_3670 = _EVAL_1048 & _EVAL_2941;
  assign _EVAL_1253 = _EVAL_2599 & _EVAL_2941;
  assign _EVAL_2414 = _EVAL_2449 & _EVAL_2047;
  assign _EVAL_568 = _EVAL_866 & _EVAL_2047;
  assign monitor__EVAL_9 = _EVAL_73;
  assign _EVAL_2547 = _EVAL_2120 & _EVAL_2971;
  assign _EVAL_836 = _EVAL_373 & _EVAL_826;
  assign _EVAL_207 = _EVAL_2532 & _EVAL_2422;
  assign _EVAL_914 = |_EVAL_2895;
  assign _EVAL_1790 = _EVAL_1391 & _EVAL_1004;
  assign _EVAL_3766 = _EVAL_2085 & _EVAL_826;
  assign _EVAL_3334 = _EVAL_173 & _EVAL_3423;
  assign _EVAL_1260 = _EVAL_1927 & _EVAL_969;
  assign _EVAL_1375 = _EVAL_1911 & _EVAL_826;
  assign _EVAL_746 = _EVAL_882 & _EVAL_154;
  assign _EVAL_952 = _EVAL_2532 & _EVAL_2317;
  assign _EVAL_2194 = |_EVAL_3323;
  assign _EVAL_2585 = _EVAL_3774 & _EVAL_3703;
  assign _EVAL_328 = _EVAL_1649 & _EVAL_295;
  assign _EVAL_893 = _EVAL_785 & _EVAL_2026;
  assign _EVAL_1331 = _EVAL_2112 & _EVAL_701;
  assign _EVAL_3195 = _EVAL_1914 & _EVAL_2941;
  assign _EVAL_2894 = _EVAL_1355 & _EVAL_2047;
  assign _EVAL_986 = _EVAL_1927 & _EVAL_3350;
  assign _EVAL_3525 = _EVAL_2181 & _EVAL_701;
  assign _EVAL_2047 = _EVAL_553 == 20'h0;
  assign _EVAL_198 = _EVAL_3126 & _EVAL_3423;
  assign _EVAL_1390 = _EVAL_1927 & _EVAL_3289;
  assign _EVAL_1425 = _EVAL_1649 & _EVAL_365;
  assign _EVAL_3135 = _EVAL_2290 & _EVAL_2047;
  assign _EVAL_2592 = _EVAL_760 & _EVAL_2941;
  assign _EVAL_897 = _EVAL_2532 & _EVAL_2185;
  assign _EVAL_497 = _EVAL_297 & _EVAL_2941;
  assign _EVAL_2393 = _EVAL_1361[6];
  assign _EVAL_2725 = _EVAL_3396 & _EVAL_1004;
  assign _EVAL_2065 = _EVAL_361 & _EVAL_2047;
  assign _EVAL_3231 = _EVAL_2972 & _EVAL_826;
  assign _EVAL_2039 = _EVAL_2949 & _EVAL_2047;
  assign _EVAL_2239 = _EVAL_2532 & _EVAL_950;
  assign _EVAL_1525 = _EVAL_1717 & _EVAL_2047;
  assign _EVAL_3411 = _EVAL_2003 & _EVAL_2047;
  assign _EVAL_3550 = _EVAL_2850[27];
  assign _EVAL_1639 = _EVAL_2830 & _EVAL_826;
  assign _EVAL_347 = _EVAL_3135 & _EVAL_701;
  assign _EVAL_1585 = _EVAL_2569 & _EVAL_2047;
  assign _EVAL_158 = _EVAL_3817 & _EVAL_2941;
  assign _EVAL_747 = _EVAL_1919 & _EVAL_2047;
  assign _EVAL_3051 = _EVAL_3585 & _EVAL_1275;
  assign _EVAL_3754 = _EVAL_1649 & _EVAL_1012;
  assign _EVAL_1742 = _EVAL_2398 & _EVAL_2941;
  assign _EVAL_494 = _EVAL_1265 & _EVAL_1004;
  assign _EVAL_3073 = _EVAL_1128 & _EVAL_701;
  assign _EVAL_2101 = _EVAL_1927 & _EVAL_2573;
  assign _EVAL_3398 = _EVAL_3125 & _EVAL_2436;
  assign _EVAL_1391 = _EVAL_761 & _EVAL_2047;
  assign _EVAL_2566 = _EVAL_2038[17];
  assign _EVAL_1656 = _EVAL_651[131];
  assign _EVAL_3795 = _EVAL_2173 & _EVAL_2941;
  assign _EVAL_2458 = _EVAL_1649 & _EVAL_2633;
  assign _EVAL_3188 = _EVAL_2857 & _EVAL_826;
  assign _EVAL_2545 = _EVAL_1166 & _EVAL_2941;
  assign _EVAL_3785 = _EVAL_2120 & _EVAL_3233;
  assign _EVAL_2553 = _EVAL_554 & _EVAL_1004;
  assign _EVAL_1965 = _EVAL_591 & _EVAL_2047;
  assign _EVAL_1725 = _EVAL_1361[11];
  assign _EVAL_486 = _EVAL_1927 & _EVAL_271;
  assign _EVAL_923 = _EVAL_1077 & _EVAL_2941;
  assign _EVAL_2108 = _EVAL_2041 & _EVAL_826;
  assign _EVAL_448 = _EVAL_2532 & _EVAL_3823;
  assign _EVAL_864 = _EVAL_2429 & _EVAL_701;
  assign _EVAL_757 = _EVAL_260 & _EVAL_2047;
  assign _EVAL_2412 = _EVAL_2007 & _EVAL_701;
  assign _EVAL_2971 = &_EVAL_3499;
  assign _EVAL_2729 = _EVAL_1649 & _EVAL_2945;
  assign _EVAL_3405 = _EVAL_2038[60];
  assign _EVAL_2955 = _EVAL_1361[5];
  assign _EVAL_3664 = _EVAL_1649 & _EVAL_2233;
  assign _EVAL_2802 = _EVAL_237 & _EVAL_826;
  assign _EVAL_234 = _EVAL_2038[116];
  assign _EVAL_3098 = _EVAL_2532 & _EVAL_2731;
  assign _EVAL_559 = _EVAL_397 & _EVAL_846;
  assign _EVAL_1420 = _EVAL_470 & _EVAL_2047;
  assign _EVAL_2596 = _EVAL_2356 & _EVAL_1429;
  assign _EVAL_2210 = _EVAL_3126 & _EVAL_2780;
  assign _EVAL_1760 = _EVAL_1611 & _EVAL_2941;
  assign _EVAL_1142 = _EVAL_2699[0];
  assign _EVAL_943 = _EVAL_1648 & _EVAL_2047;
  assign _EVAL_3058 = _EVAL_3054 & _EVAL_701;
  assign _EVAL_1865 = _EVAL_3853 & _EVAL_701;
  assign _EVAL_3194 = _EVAL_3774 & _EVAL_1470;
  assign _EVAL_2154 = _EVAL_397 & _EVAL_481;
  assign _EVAL_1955 = _EVAL_2850[15];
  assign _EVAL_1378 = _EVAL_2038[36];
  assign _EVAL_2893 = _EVAL_1361[30];
  assign _EVAL_3522 = _EVAL_682 & _EVAL_701;
  assign _EVAL_3783 = _EVAL_1361[13];
  assign _EVAL_2859 = _EVAL_1427 & _EVAL_1004;
  assign _EVAL_3448 = _EVAL_2532 & _EVAL_635;
  assign _EVAL_2743 = _EVAL_3009 & _EVAL_2941;
  assign _EVAL_2409 = _EVAL_2644 & _EVAL_701;
  assign _EVAL_2172 = _EVAL_3750 & _EVAL_2047;
  assign _EVAL_3582 = _EVAL_1927 & _EVAL_698;
  assign _EVAL_1971 = _EVAL_1479 & _EVAL_2941;
  assign _EVAL_1163 = _EVAL_2532 & _EVAL_271;
  assign _EVAL_3144 = _EVAL_501 & _EVAL_2047;
  assign _EVAL_3833 = _EVAL_2850[9];
  assign _EVAL_1679 = _EVAL_1926 & _EVAL_2047;
  assign _EVAL_2273 = _EVAL_2038[40];
  assign _EVAL_2953 = _EVAL_1649 & _EVAL_3681;
  assign _EVAL_3372 = _EVAL_1159 & _EVAL_154;
  assign _EVAL_662 = _EVAL_3562 & _EVAL_3232;
  assign _EVAL_3344 = _EVAL_2532 & _EVAL_263;
  assign _EVAL_3310 = _EVAL_2993 & _EVAL_2678;
  assign _EVAL_1296 = _EVAL_1927 & _EVAL_2176;
  assign _EVAL_2994 = _EVAL_2850[10];
  assign _EVAL_2025 = _EVAL_2984 & _EVAL_2941;
  assign _EVAL_825 = _EVAL_1915 & _EVAL_2047;
  assign _EVAL_2538 = _EVAL_2038[19];
  assign _EVAL_2883 = _EVAL_1649 & _EVAL_3732;
  assign _EVAL_438 = _EVAL_2532 & _EVAL_3808;
  assign _EVAL_3499 = _EVAL_1361[7:0];
  assign _EVAL_2937 = _EVAL_2532 & _EVAL_187;
  assign _EVAL_1291 = _EVAL_1649 & _EVAL_3852;
  assign _EVAL_3698 = _EVAL_2038[93];
  assign _EVAL_3365 = _EVAL_2038[126];
  assign _EVAL_1653 = _EVAL_2532 & _EVAL_1475;
  assign _EVAL_2162 = |_EVAL_315;
  assign _EVAL_3203 = _EVAL_2993 & _EVAL_1868;
  assign _EVAL_3004 = _EVAL_173 & _EVAL_370;
  assign _EVAL_1629 = _EVAL_1649 & _EVAL_3622;
  assign _EVAL_1974 = _EVAL_1284 & _EVAL_701;
  assign _EVAL_932 = _EVAL_3066 & _EVAL_701;
  assign _EVAL_2690 = _EVAL_229 & _EVAL_2047;
  assign _EVAL_656 = _EVAL_1927 & _EVAL_2301;
  assign _EVAL_2470 = _EVAL_2302 & _EVAL_2047;
  assign _EVAL_1602 = _EVAL_2850[21];
  assign _EVAL_1834 = _EVAL_2993 & _EVAL_2541;
  assign _EVAL_2200 = _EVAL_2924 & _EVAL_2047;
  assign _EVAL_3812 = _EVAL_2414 & _EVAL_1004;
  assign _EVAL_950 = _EVAL_2038[34];
  assign _EVAL_3694 = _EVAL_3562 & _EVAL_1111;
  assign _EVAL_1734 = _EVAL_2850[31];
  assign _EVAL_3491 = out_back__EVAL_2;
  assign _EVAL_705 = _EVAL_397 & _EVAL_1176;
  assign _EVAL_2684 = _EVAL_1131 & _EVAL_826;
  assign _EVAL_3581 = _EVAL_1639 & _EVAL_2941;
  assign _EVAL_1870 = _EVAL_1649 & _EVAL_625;
  assign _EVAL_1701 = _EVAL_2038[91];
  assign _EVAL_1567 = _EVAL_1924 & _EVAL_701;
  assign _EVAL_2574 = _EVAL_397 & _EVAL_3761;
  assign _EVAL_1572 = _EVAL_2993 & _EVAL_370;
  assign _EVAL_2183 = _EVAL_2749 & _EVAL_2047;
  assign _EVAL_960 = _EVAL_2038[84];
  assign _EVAL_3233 = &_EVAL_3805;
  assign _EVAL_2908 = |_EVAL_3413;
  assign _EVAL_3764 = |_EVAL_2994;
  assign _EVAL_3019 = _EVAL_200 & _EVAL_1004;
  assign _EVAL_626 = _EVAL_2105 & _EVAL_1004;
  assign _EVAL_1669 = _EVAL_397 & _EVAL_3300;
  assign _EVAL_2085 = _EVAL_1649 & _EVAL_1731;
  assign _EVAL_1287 = _EVAL_3727 & _EVAL_701;
  assign _EVAL_1319 = _EVAL_2674 & _EVAL_2941;
  assign _EVAL_1897 = _EVAL_1519 & _EVAL_2047;
  assign _EVAL_3549 = |_EVAL_1003;
  assign _EVAL_2036 = _EVAL_839 & _EVAL_2941;
  assign _EVAL_1198 = _EVAL_174 & _EVAL_701;
  assign _EVAL_3269 = _EVAL_3585 & _EVAL_1930;
  assign _EVAL_3666 = _EVAL_1649 & _EVAL_3148;
  assign _EVAL_3003 = _EVAL_1649 & _EVAL_2879;
  assign _EVAL_823 = _EVAL_2532 & _EVAL_3631;
  assign _EVAL_2539 = _EVAL_3126 & _EVAL_3498;
  assign _EVAL_2086 = _EVAL_3464 & _EVAL_2941;
  assign _EVAL_1632 = _EVAL_2532 & _EVAL_1318;
  assign _EVAL_1914 = _EVAL_926 & _EVAL_826;
  assign _EVAL_389 = _EVAL_706 & _EVAL_1004;
  assign _EVAL_3544 = _EVAL_1115 & _EVAL_2047;
  assign _EVAL_2299 = _EVAL_3660 & _EVAL_2941;
  assign _EVAL_2960 = _EVAL_3774 & _EVAL_1708;
  assign _EVAL_1732 = _EVAL_3570 & _EVAL_1004;
  assign _EVAL_3562 = _EVAL_1888 & _EVAL_826;
  assign _EVAL_659 = _EVAL_2038[8];
  assign _EVAL_1345 = _EVAL_1649 & _EVAL_693;
  assign _EVAL_1082 = _EVAL_1649 & _EVAL_3572;
  assign _EVAL_1616 = _EVAL_2625 & _EVAL_2941;
  assign _EVAL_767 = _EVAL_1649 & _EVAL_3249;
  assign _EVAL_558 = _EVAL_357 & _EVAL_826;
  assign _EVAL_2192 = _EVAL_3774 & _EVAL_3423;
  assign _EVAL_2544 = _EVAL_1649 & _EVAL_3672;
  assign _EVAL_2662 = _EVAL_1851 & _EVAL_2941;
  assign _EVAL_475 = _EVAL_2038[38];
  assign _EVAL_2184 = _EVAL_1649 & _EVAL_3456;
  assign _EVAL_711 = _EVAL_1332 & _EVAL_2047;
  assign _EVAL_1290 = _EVAL_1390 & _EVAL_2047;
  assign _EVAL_255 = _EVAL_1927 & _EVAL_3631;
  assign _EVAL_1092 = _EVAL_3843 & _EVAL_2047;
  assign _EVAL_186 = _EVAL_2323 & _EVAL_826;
  assign _EVAL_1927 = _EVAL_159 & _EVAL_3846;
  assign _EVAL_3478 = _EVAL_3585 & _EVAL_3224;
  assign _EVAL_1606 = _EVAL_3562 & _EVAL_1245;
  assign _EVAL_1495 = _EVAL_3774 & _EVAL_1868;
  assign _EVAL_1035 = _EVAL_1361[1];
  assign _EVAL_634 = _EVAL_1149 & _EVAL_1004;
  assign _EVAL_1911 = _EVAL_1649 & _EVAL_1248;
  assign _EVAL_1128 = _EVAL_242 & _EVAL_2047;
  assign _EVAL_1995 = _EVAL_2854 & _EVAL_2047;
  assign _EVAL_2037 = _EVAL_1649 & _EVAL_3462;
  assign _EVAL_761 = _EVAL_1927 & _EVAL_2764;
  assign _EVAL_2854 = _EVAL_1927 & _EVAL_329;
  assign _EVAL_2587 = _EVAL_1927 & _EVAL_1685;
  assign _EVAL_459 = _EVAL_1649 & _EVAL_1787;
  assign _EVAL_2434 = _EVAL_3580 & _EVAL_2047;
  assign _EVAL_830 = _EVAL_1849 & _EVAL_1004;
  assign _EVAL_931 = _EVAL_1649 & _EVAL_403;
  assign _EVAL_938 = _EVAL_558 & _EVAL_2941;
  assign _EVAL_1126 = _EVAL_1649 & _EVAL_2103;
  assign _EVAL_3841 = _EVAL_2757 > 7'h0;
  assign _EVAL_2467 = _EVAL_742 & _EVAL_2941;
  assign _EVAL_618 = _EVAL_1045 & _EVAL_1004;
  assign _EVAL_2816 = _EVAL_3826 & _EVAL_826;
  assign _EVAL_3472 = _EVAL_1649 & _EVAL_463;
  assign _EVAL_1945 = _EVAL_2850[6];
  assign _EVAL_806 = _EVAL_1927 & _EVAL_2962;
  assign _EVAL_2423 = _EVAL_2172 & _EVAL_1004;
  assign _EVAL_157 = _EVAL_3688 & _EVAL_2047;
  assign _EVAL_878 = _EVAL_1927 & _EVAL_2411;
  assign _EVAL_2680 = _EVAL_1649 & _EVAL_369;
  assign _EVAL_1104 = _EVAL_173 & _EVAL_2540;
  assign _EVAL_3678 = _EVAL_397 & _EVAL_3606;
  assign _EVAL_2076 = _EVAL_2244 & _EVAL_701;
  assign _EVAL_3640 = _EVAL_2365 & _EVAL_2941;
  assign _EVAL_2764 = _EVAL_2038[52];
  assign _EVAL_1154 = _EVAL_3126 & _EVAL_2540;
  assign _EVAL_474 = _EVAL_3774 & _EVAL_2096;
  assign _EVAL_942 = |_EVAL_2735;
  assign _EVAL_2644 = _EVAL_3578 & _EVAL_2047;
  assign _EVAL_3136 = _EVAL_2684 & _EVAL_3087;
  assign _EVAL_1177 = |_EVAL_1006;
  assign _EVAL_1470 = |_EVAL_1233;
  assign _EVAL_542 = _EVAL_2775[3];
  assign _EVAL_636 = _EVAL_717 & _EVAL_2971;
  assign _EVAL_3407 = |_EVAL_3250;
  assign _EVAL_2016 = _EVAL_2993 & _EVAL_2635;
  assign _EVAL_2116 = _EVAL_363 | _EVAL_110;
  assign _EVAL_2540 = |_EVAL_3689;
  assign _EVAL_2947 = _EVAL_2038[50];
  assign _EVAL_155 = _EVAL_2610 & _EVAL_197;
  assign _EVAL_2746 = _EVAL_3012 & _EVAL_2047;
  assign _EVAL_3295 = _EVAL_235 & _EVAL_2047;
  assign _EVAL_197 = _EVAL_3093[126:0];
  assign _EVAL_1858 = _EVAL_1406 & _EVAL_826;
  assign _EVAL_791 = _EVAL_2532 & _EVAL_201;
  assign _EVAL_3083 = _EVAL_3042 & _EVAL_701;
  assign _EVAL_1716 = _EVAL_3164 & _EVAL_2047;
  assign _EVAL_1410 = _EVAL_1927 & _EVAL_1775;
  assign _EVAL_1580 = _EVAL_3664 & _EVAL_826;
  assign _EVAL_460 = _EVAL_805 ? 8'hff : 8'h0;
  assign _EVAL_1827 = _EVAL_3125 & _EVAL_1930;
  assign _EVAL_1798 = _EVAL_2532 & _EVAL_3365;
  assign _EVAL_2606 = _EVAL_2532 & _EVAL_2947;
  assign _EVAL_1737 = _EVAL_3561 & _EVAL_1004;
  assign _EVAL_1714 = _EVAL_756 & _EVAL_701;
  assign _EVAL_675 = _EVAL_1474 & _EVAL_826;
  assign _EVAL_3532 = _EVAL_2183 & _EVAL_1004;
  assign _EVAL_3178 = _EVAL_587 & _EVAL_2047;
  assign _EVAL_3477 = _EVAL_1927 & _EVAL_188;
  assign _EVAL_250 = _EVAL_1819 & _EVAL_2047;
  assign _EVAL_3170 = _EVAL_882 & _EVAL_802;
  assign _EVAL_2304 = _EVAL_818 & _EVAL_2941;
  assign _EVAL_3470 = _EVAL_1927 & _EVAL_2359;
  assign _EVAL_934 = _EVAL_1840 & _EVAL_1004;
  assign _EVAL_2699 = _EVAL_1560 - 1'h1;
  assign _EVAL_2272 = _EVAL_2038[125];
  assign _EVAL_2718 = _EVAL_2038[65];
  assign _EVAL_2400 = _EVAL_2669 & _EVAL_2047;
  assign _EVAL_1908 = _EVAL_946 & _EVAL_2047;
  assign _EVAL_2164 = _EVAL_491 & _EVAL_826;
  assign _EVAL_1259 = _EVAL_767 & _EVAL_826;
  assign _EVAL_981 = _EVAL_2058 & _EVAL_2941;
  assign _EVAL_3044 = _EVAL_84[0];
  assign _EVAL_2806 = _EVAL_2353 & _EVAL_2047;
  assign _EVAL_145 = _EVAL_1633 & _EVAL_2941;
  always @(posedge _EVAL_9) begin
    if (_EVAL_110) begin
      _EVAL_1581 <= 1'h0;
    end else if (_EVAL_3439) begin
      _EVAL_1581 <= _EVAL_1917;
    end
    _EVAL_1777 <= _EVAL_2296 & _EVAL_304;
    if (_EVAL_110) begin
      _EVAL_2890 <= 1'h0;
    end else if (_EVAL_3439) begin
      _EVAL_2890 <= _EVAL_1560;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3163 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ba5dc84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1861 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4962830)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1938 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac41f6b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3555 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84a4413d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3838 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8968dbbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3662 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9fad6f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1399 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c8cab05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3281 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bfa7ecf6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3314 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1c970ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1728 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e3fdef3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3026 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22fb967e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_901 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dbd356e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3517 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9942b0d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1769 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d876c4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_831 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2406136)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2100 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be588fa5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_233 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a5459)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3839 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1a6aa78f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1047 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(893ea67e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3478 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a07728f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3592 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d1725d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2259 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b5699b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3598 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8214f66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_426 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62fa06de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2328 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72a2c568)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_898 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88db11a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_754 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1456666e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_835 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85266753)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2368 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dadcc87e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_961 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ac6023d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3351 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72eb2289)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2526 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7c9a7bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3785 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f650f9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1164 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ccfcd32c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_599 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(624e6115)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1228 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ac5933b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_888 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa8d1607)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3814 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9f5ae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2630 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cec1fdb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3509 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3cdb0fb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1476 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfec98fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1747 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77c51635)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1616 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21ce864)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3088 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(945b7585)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1521 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a6615f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_863 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20d77b7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1531 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf97423c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3658 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(14e2b4ce)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_541 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60b442e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3190 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50c9ee69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_769 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(783846da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2651 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acb6db03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3228 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5f4d3f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1121 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(59a11683)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2688 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f101045a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2432 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76bb409e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_684 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19307a1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2958 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1dc30742)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3673 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25cc4205)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3629 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35ea82c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2457 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95c10267)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1462 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(114340b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3621 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d04fa58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1216 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0b6b74)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2208 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1522e782)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1154 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ddc55aeb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_613 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d23a3117)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3779 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ebf52532)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1686 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6355783b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1719 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d30da542)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1038 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65d6cab8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1484 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c8d41d7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2382 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba7499b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3230 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a688f897)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2546 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26d602c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_868 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4993c71)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2142 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bb09f0ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2916 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7c03595)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2022 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ebd219b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2499 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3bae3e7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2866 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b4cca59)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2756 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c54819e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2237 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24270004)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1150 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af017c60)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3141 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(881a7417)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_580 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b997b4a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_932 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(445ce47a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2015 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(acc61884)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2299 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c3739bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1584 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5b6b3cb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_662 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3dd2ead)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_777 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be1fffd5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2829 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7cab0bd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2006 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd81f83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2443 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(289e0935)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3445 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91e32072)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2578 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b9e74e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1013 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f463cc9a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1054 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(112d2e05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_319 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb34ec42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1715 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be9b128)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3309 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98e562c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1958 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3506ade0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3500 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca3398fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3553 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4a5f604)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_447 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1104dcb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2744 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6757642)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1068 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38985a4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1772 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62fde11b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_786 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26ea769d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2774 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(177b4784)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2785 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b91c3018)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_545 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b91dc28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2990 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(adc61929)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3208 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e92746ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_799 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df4118e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2886 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c3799db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2511 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e2ebd86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2504 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0be939c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1305 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16d291d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2952 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c7298049)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1961 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62071bd5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1204 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(546fe1a5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2412 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d3f1179)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3192 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd3dd7ea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_908 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1350915f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3443 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36251c15)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1972 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d521ddbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3563 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dadc6a47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1735 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c759992)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3693 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ae87d1a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2539 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(346ff6ef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1227 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe687838)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_923 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e22095)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2790 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df99a5fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2583 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f03b7f8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1324 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(390479e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3740 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(263d43f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3031 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4859365c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2097 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80377a7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_444 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(232efff2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_551 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b2776d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_604 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b41a8a04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3269 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(425b5862)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1363 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94dfeaf1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3552 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7bf139d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2475 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b059656d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_537 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(be61e589)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3286 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65259a6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3179 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65544ba1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2497 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(467bea5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2016 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92e87396)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_634 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c115f4b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3025 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(939d0e79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_618 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2b244be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1105 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8acb27b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2265 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4965040e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3601 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b28d853)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_563 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1211349)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1513 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(999c8ee7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2522 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1aad0bf6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1563 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f57eeb6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2773 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a0ae69a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1401 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bef156a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3813 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90961da7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2964 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1572d597)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3379 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(850dd615)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1279 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6cb2f4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2960 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bb18dcb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1755 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(55dbd948)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_816 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d95e016a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3348 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76b08020)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2401 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87a0eb87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1234 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c4add68)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1108 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(437562df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_772 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1deba7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1469 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6721b48b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_984 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad7d692f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2501 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8baa80e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3356 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2b4fcdf5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2658 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7f24da2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2657 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd8ff769)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2545 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9458305)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3078 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e9a2c4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2611 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6977dbd4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3665 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f173c00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1939 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9975f7a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3522 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9323ee72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2190 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe4461be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2959 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1379530)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1377 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1949b89a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2310 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a68e6639)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1953 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4c5c71a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_704 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73a35d3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3380 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4022e3c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3789 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ad9ffdc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1502 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5037d4dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_264 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96fbfab2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2046 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc220dca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2374 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdb1e4b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1744 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1baa3c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2736 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af628d4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3028 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79b71d98)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_572 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e36b2f3d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2567 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1c906a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3730 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e550f7c7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2117 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6065183)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1614 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9ba16f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3173 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c861b44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3733 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ee423a3c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3136 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac55abca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3117 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4c5278e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2560 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a19c515)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2582 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7481bbe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2000 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d65448e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3722 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e97254f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1445 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3202bf56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1724 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57a01d48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1207 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7a69598)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1458 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d0901dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2642 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab9b2d22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3677 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6a16ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_335 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(33c8f9dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1980 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e259dcef)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1230 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ee5e746)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2032 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(183bdd5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2876 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45b637fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2210 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48500e40)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3325 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e0321c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_708 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ddaae7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_884 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d0d8639)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1748 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba22dccf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_528 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29afa792)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3227 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c509f48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3738 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fbc344a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_205 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7c4ad13)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_620 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fb1c8f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2270 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba6b020e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1253 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a558f030)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3494 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f715f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1231 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7da976ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2480 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6d9e706)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3181 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6f3071a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_764 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76a9b512)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1720 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d0e5451)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3720 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(adda4547)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2954 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70bd0360)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1790 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af641ea1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2673 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfa2456e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_837 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4e0e7d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_871 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(743876bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3056 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(728e5185)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2577 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35e782cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1845 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(76fce6a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_244 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27162a8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_947) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1574 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cebc098)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2372 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dcc369f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1309 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8e19b65)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2574 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5909f3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_431 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ab59dfe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1423 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a6883bf2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1662 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(137c2ffa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2087 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(698488f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3482 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9cb23be2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2846 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f07d50e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3032 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d9ef94a7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3008 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5d4398d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3023 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eaa31402)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2454 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27d02c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2271 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3744487)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2280 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f9f283e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_387 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5dad36d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2093 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4468e83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1188 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c1def70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3771 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a887739d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1132 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ffc28ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3594 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(75444f8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1596 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6439cd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2752 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bcd0ade7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1491 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(232efbe9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_407 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6866d2e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1808 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5beb6f8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_579 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d7e1971f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1778 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f9db4f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2664 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb4cc22d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2510 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92307ccb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3614 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce71a5e2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2859 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e738eb16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2242 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3add280)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_730 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(918934de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1331 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e26ef66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2818 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e52d1dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1161 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(278af90b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3581 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(915f6739)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3347 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e06cfd3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3645 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(977a3267)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_158 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ae6aad1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1654 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9720f1f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2040 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a872b008)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3719 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8e0c941)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1992 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(601133c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2327 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea0be704)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_485 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82086431)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2266 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(896d2dae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_857 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9adb27)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1301 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df775c46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1874 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d77ec1af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3518 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eadefb19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_977 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd106275)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_654 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c261e01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2547 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9ffaab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1825 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fce3a773)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2409 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cfef426)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1249 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ffa3e19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2931 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0a5695d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1097 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bcc91241)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2291 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d52395f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2010 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3824a881)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3113 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(301c72c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1820 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(192fda56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2044 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3163058e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2358 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c718caf2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3515 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49817b42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2666 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e652e2d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1971 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66ed3ded)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1022 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fabcf24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1538 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7428950)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1362 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44004d22)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_372 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa98f806)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3487 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efe484ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_864 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e446e271)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1007 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68570232)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2402 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6317f86)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_830 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a9cc734)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2403 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f95eebd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_972 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9b2f11f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_162 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db684ea9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2329 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(daad96b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3371 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b7720c06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_928 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(46256b5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3466 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5261fb9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2269 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8188993)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1055 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51dfcfb4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3670 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6733887d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_715 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(581a1383)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_968 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(103e8c1f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1816 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab9b5030)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_441 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8262f95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2318 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(381156fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1904 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9de1540)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3634 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac044f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1328 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(863d1d7a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2330 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(762b6ce6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1951 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3165769b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2513 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1214e7dc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1261 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5529c5ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_649 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95e7ae3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_637 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5404d12f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1913 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b992a151)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1652 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(409e2cb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_418 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65a16ea9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2073 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a0d0f717)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_453 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5840bbd1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1916 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b62c4df5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2025 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af17b35c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1388 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f002e884)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1389 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d317f47e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3641 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4d699e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_800 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c12784d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3197 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61cc2438)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1287 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62426c6e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_180 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b3ee62f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2590 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f133c178)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1344 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d03285d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2278 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a31e7f9c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1609 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a66c11ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3694 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5ecca4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3787 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4de5c009)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3282 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db188c38)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3097 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fc09333)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_283 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d0b2c4d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2351 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb6af9f5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2887 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c845d50)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a7230f2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2362 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35809459)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3094d605)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3229 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e297ba55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2689 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef3541eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_934 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fcf32652)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1552 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(841ff229)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1759 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74e3cfd3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_389 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(229ed2ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3194 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4bd3b2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_798 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f8fa5723)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2229 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(99525b90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3390 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(812795f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1426 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d97838e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2170 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(105180f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3547 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3cf46fd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_658 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6834d03f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1cd50cf9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2307 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2417750)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3022 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ce0bf02e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2219 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7293e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2336 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb84f95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2815 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e1bb8697)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1906 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4694dba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3277 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f172c32c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_619 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aeeda00f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2609 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cf4978b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3083 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21f6f7fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_377 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c9e6a24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2751 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d451605)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1782 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d5863c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2594 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e23b63f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2425 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2d3d5c01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1726 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c21d0cd0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_629 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43a050)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3248 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9082049b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2066 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7435ee48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1240 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4ab8071)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2919 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d820ab8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1107 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7418d0a4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2882 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e3cea9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3091 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4139dd8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3170 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(85707950)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3452 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd617728)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2076 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(61265115)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2036 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b727370)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_626 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c0c6426e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3160 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab03540b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1613 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4305d651)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_519 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e11a5bdd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_305 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2596741e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1676 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8401514)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2858 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7149b034)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1263 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2542308b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_896 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f91641f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_347 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d2f6b85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_833 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f712186)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2489 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9b4d53d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1737 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97bbb839)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_885 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c7a0ecf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1664 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b471899)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1922 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3f7f1475)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3052 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f4485a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_509 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cba7d75e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2189 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b02e7a45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_192 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e0005db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1080 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2dd39bf0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_746 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9219b106)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2963 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(249035c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1494 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9dc5e1b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1570 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e817dd21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2740 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba3dde56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2819 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42762d5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_862 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9640ee9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2154 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed5a5a5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_636 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(648d7e93)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2973 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfa2456e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_705 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b5168e0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_348 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ca6efbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1615 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(918934de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_861 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f9ffef11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_533 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca9802b8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_2332) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2734 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2c0f05b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2052 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7d54de3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1146 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d422188d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2430 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1f0cc8e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1709 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(646b0468)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3809 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42272e42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3359 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc5e29b5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3676 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e170fbe7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_262 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2426d6a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2089 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40088174)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1742 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(897f5412)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_327 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c84a7ba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1213 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ad2d7804)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1522 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(521b08ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2123 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5792e62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1746 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a30624)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_893 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c8ae2cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_687 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9069fe3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_680 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e45c9967)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1235 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1b84099)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_239 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f5b56fad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3382 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3bae136)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2113 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2e1aedc8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3064 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2027b4c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2367 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34d0a90b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_765 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(609d7826)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1823 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(551660d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3372 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a2b6c138)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_971 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3bd5b5d8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3609 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aabcb82a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2930 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7a23123)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_494 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6cf665fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3745 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(907547dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_891 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45a6e53f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_666 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(233991e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_259 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfd56710)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2072 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74a32a81)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2585 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c0a5135)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1729 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c867d8f1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3139 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3dcd164)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1353 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a0c3dee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2119 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6ae8e255)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1050 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca0dda36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2636 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ffebe49e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1136 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e03cc0e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3131 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f2201ff7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_924 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c582ce99)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1357 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a6a71cb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_676 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1c836f82)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1098 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ec571fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1572 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9fa663a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3713 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c23bd25)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2304 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(43ed51fb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1387 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fedcd08e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3159 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf029759)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1863 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(779db55e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1975 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bb015d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_530 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cb45272)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3180 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e0bf383)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2750 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7df843e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3608 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b67b11db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2588 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd63f984)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1567 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9024cc03)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_821 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2eab5180)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_814 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(39612b88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3334 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89b27769)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1409 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(853fd3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2851 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e7906408)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3408 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aa6d091f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_622 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b116e33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_291 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d68c2f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2899 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db8cd8d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3532 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3396285d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1196 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e826bb6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2596 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c034e8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2001 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(295f56cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_947) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b098f87)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3296 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(27faa01)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1206 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(275787af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_941 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94f60929)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1044 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1156d55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_221 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2997df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1383 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb65b693)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2177 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(492c96f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_275 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15b5f41)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2371 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d8b1e86b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_912 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a3b8e4f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3137 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f33b3dec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3519 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b114f228)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_681 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bef6f315)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2494 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4648114e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3820 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af4370ed)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3068 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(91fce163)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1974 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37ef5e0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2283 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(517eb870)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2786 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b5deae14)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_358 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c10ad29)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_442 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4620a25f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2333 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ef99f79d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3149 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1842321d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1991 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c20ad62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2741 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca84beff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_395 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25e02161)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3586 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5a6bef8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1215 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f52d457)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_633 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e434a6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3079 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a70a3806)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1319 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(51325f47)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2602 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb7a08b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1042 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e6d3a6d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1829 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(38da8270)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1750 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d03cffc3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3203 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87042743)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1545 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35089ca0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3364 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2e080c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2435 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31b55575)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1575 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b61ba943)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2410 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d40a9a1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3019 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(40c712da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2334 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6af1eda)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3424 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4a18d16)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1198 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7db9ddb2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2054 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c66ab3a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1109 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c23d078)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2225 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0176641)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1037 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84c38459)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2766 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32937171)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3812 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57d8f18a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1896 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d67713d1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1266 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c2599b6a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3678 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c18c276)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1079 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9ef12104)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_311 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a0b68f0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1100 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2968aff0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3339 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ff8c485)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3447 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe795697)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3525 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(68dcb78e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_737 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21cb7a48)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_749 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(724cb412)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1817 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25751bad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2267 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b6f8742)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_333 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df70b364)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_958 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3081f069)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3321 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(600bb397)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2661 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b528e78)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1386 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82c659fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_489 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25cb79eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3121 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c638c978)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3049 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(efca4cde)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1376 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8135577a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1019 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c5e18e9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1539 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f38a436e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3212 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(124a70a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1168 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d41730ca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2662 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e31d75c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1905 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(688217a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1827 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(469a9f5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1933 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3ad7ec8c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_917 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ccc5d37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3707 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(197f47da)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_851 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(42b18f72)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3090 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6f83c97)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1218 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6057eea)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1110 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ec0623a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3415 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b6909cd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3728 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a8836804)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2665 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(391f61b1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1620 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79a9ffa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2058b962)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1352 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(66ce89de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2631 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4b425d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3283 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5808c3c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1834 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3d83c5e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1160 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cdd707fc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2864 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5d9d82fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1075 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b665eac7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1326 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3b7ae180)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1591 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c02c2ee0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2553 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8673aa6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1104 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e95e051d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_493 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6b49f53)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2420 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f93e256c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_750 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e8d339bc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2232 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b8e98ab)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2647 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1090f588)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2807 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba772983)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1321 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(832d5aae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3419 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78565376)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2620 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(411d7de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1841 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b462c85a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3640 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa28108f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2338 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e792d337)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1051 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e7a2588)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_432 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ea40e43e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1714 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9daaecfc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2141 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3a6b5e62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_741 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eefa8a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_497 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(500d1133)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_346 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3b69555)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2247 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ec043f5a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1477 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e742121b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3539 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(747379d3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_521 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(962e6a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1606 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4c9109f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3752 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52dc363)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_198 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41adc566)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3623 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba6d7bad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2086 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78135d3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_734 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(29391964)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2824 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21bdd613)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2967 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2aec3436)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1865 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d9e04a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_312 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41ccd030)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3058 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e61b6dcc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_796 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50839510)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_300 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48cb5b7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3602 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e115af1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_611 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f7f0f113)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1831 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aeb61f9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2110 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73923af3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3410 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(643588ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2467 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3a7d2c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1642 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(52eb643b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_439 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74e67941)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2638 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(92f91a2e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3542 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9e144f62)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3453 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f01c6ccf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3574 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16be7395)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_550 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d34f1b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2506 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3b8955b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1297 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(82e5fc45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1250 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2db14a0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3070 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19b7e506)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2976 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5832d936)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_561 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1b7b991)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_191 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(faee1a58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1573 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f6670166)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1756 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(845d30d4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_252 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80d73272)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1705 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(80b05edd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_716 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30f4108f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2762 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2616fc2a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2107 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6799c025)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2725 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(defb8f11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_393 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5db822cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1327 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c180aec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3004 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5657098)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3196 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4d584761)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3541 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e05d670)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_714 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9960e371)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_406 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b38fd55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2390 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de00b5a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_145 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c32b2579)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1202 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(96c34936)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_606 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d632c425)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_474 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de51b964)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1273 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(313b7235)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_652 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c0f3612)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2743 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7ac5bd7b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1669 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c40f534c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1402 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20acaa1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3010 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6bda8fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1225 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d84785b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1837 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f4ffd68a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1217 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b09395ff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_575 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(10b4f14f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2201 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e38a8ea7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3795 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(35e66492)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_151 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f93740f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1256 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(918934de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2825 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74bdb460)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_725 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4c23d784)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_887 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86777a0f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1885 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(90f3632a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_590 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbfc8354)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1152 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca8f493)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_286 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(854a4d94)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2151 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8614073)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2198 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1fc3c75)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_420 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(32d39ac2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_559 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88dd098d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2884 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(903c98c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1267 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74b52ed9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2646 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d4655d4e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3735 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3b99ec3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3338 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(49512aa6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1628 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d206504b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3045 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d6fd9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2357 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2484a0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3617 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f2821c3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2592 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8e53adaa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_690 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9fb34f4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3484 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6518becd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1103 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58a945ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1049 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2ba9b80)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3784 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c9655b91)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2683 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60d77b84)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1672 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(202cb54f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3715 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ecb503e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_452 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9250318f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_508 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(754aa716)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1860 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2c3f2a09)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3195 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4e8ab9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2939 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(71f7421b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_596 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de7319fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3073 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(df203fa3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_632 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb1e4b06)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2920 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(caecac2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2192 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(207525c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3543 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36d1380)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3176 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a022eae)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1320 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a7121de)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_822 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b1febd1d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1535 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(adefd03a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3053 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9beb42c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3182 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(747c4997)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1530 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2b0faa2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3065 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(440d912d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2206 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(25067d83)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1753 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2fc1cd21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_981 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a15d8d28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_723 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(adc4ecbb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3048 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f0ecb36)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1797 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbb4cd3f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1490 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(88db4f2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_803 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4982c0df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1495 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(eb9dfe4a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_938 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d6cca93b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_510 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8493d4c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2246 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dee983f3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2600 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e09b7733)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2820 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6bd2e854)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3062 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edda6ae6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_922 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7899c19b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2180 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2ae8c79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2925 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1420597e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1818 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(87ae8a69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2305 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(72e42947)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2615 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(31f35cba)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_867 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(97ce6a0a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2068 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dfa2456e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_503 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c97c5e95)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1663 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7554040e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2011 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ee927be)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1397 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1808627c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1760 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(57a7d15d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1699 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ca5fc8f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1468 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0dc7b5f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2360 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a19ee0e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2082 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f006d96f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3051 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b8a815b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1864 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b1444e5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1586 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3e3acc9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1691 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3aedfe4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3799 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(98054e23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2551 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1dfd7960)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2042 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4db3ab7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3146 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9b34d20)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3168 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73b34e6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_795 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(54cd5b8b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1886 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(81f35739)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_548 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e22783c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1791 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bbdfeb27)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_223 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(22d3194e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_320 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c7a6b07)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_465 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e328dc88)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1651 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(30291c2c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb53378f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3398 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2dafac9f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2423 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8a490907)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1155 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fda0655c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2536 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4ab9374f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3310 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6718bfc3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1727 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f08466c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_2837 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34267dc6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3699 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd733f56)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3763 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cce39718)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1394 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf43dcf6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_3840 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(466bb9db)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_1732 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b179dd27)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_356 & _EVAL_3332) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4a4c6aa4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_1581 = _RAND_0[0:0];
  _RAND_1 = {4{`RANDOM}};
  _EVAL_1777 = _RAND_1[126:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_2890 = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
