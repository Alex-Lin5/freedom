//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_150_assert(
  input         _EVAL,
  input  [1:0]  _EVAL_0,
  input  [9:0]  _EVAL_1,
  input  [2:0]  _EVAL_2,
  input         _EVAL_3,
  input  [25:0] _EVAL_4,
  input  [2:0]  _EVAL_5,
  input         _EVAL_6,
  input         _EVAL_7,
  input         _EVAL_8,
  input  [9:0]  _EVAL_9,
  input         _EVAL_10,
  input  [3:0]  _EVAL_11,
  input  [2:0]  _EVAL_12,
  input  [1:0]  _EVAL_13,
  input         _EVAL_14
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [575:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_15;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire [575:0] _EVAL_21;
  wire  _EVAL_22;
  reg  _EVAL_23;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  reg [1:0] _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire [3:0] _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire [1:0] _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire [25:0] _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire [26:0] _EVAL_64;
  wire  _EVAL_65;
  wire [1:0] _EVAL_66;
  wire  _EVAL_67;
  reg [9:0] _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  reg [25:0] _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  reg  _EVAL_75;
  wire  _EVAL_76;
  wire [575:0] _EVAL_77;
  wire  _EVAL_78;
  wire [1:0] _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  reg [2:0] _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_85;
  wire  _EVAL_86;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_87;
  wire [575:0] _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire [26:0] _EVAL_92;
  wire  _EVAL_93;
  wire [1:0] _EVAL_95;
  wire  _EVAL_96;
  wire [4:0] _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire [1023:0] _EVAL_108;
  wire  _EVAL_110;
  wire [1:0] _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire [31:0] _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_123;
  wire [25:0] _EVAL_124;
  reg  _EVAL_125;
  wire  _EVAL_127;
  wire [3:0] _EVAL_128;
  wire [1023:0] _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire [3:0] _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire [26:0] _EVAL_137;
  wire  _EVAL_138;
  reg [31:0] _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire [575:0] _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire [575:0] _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire [575:0] _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire [32:0] _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire [3:0] _EVAL_166;
  wire  _EVAL_167;
  wire [1:0] _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire [25:0] _EVAL_176;
  wire  _EVAL_177;
  reg [9:0] _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  wire  _EVAL_187;
  reg  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  reg [575:0] _EVAL_194;
  wire  _EVAL_196;
  reg [2:0] _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire [575:0] _EVAL_220;
  wire  _EVAL_221;
  wire [1:0] _EVAL_222;
  wire  _EVAL_223;
  wire [1023:0] _EVAL_224;
  wire  _EVAL_225;
  reg [2:0] _EVAL_226;
  wire [575:0] _EVAL_227;
  reg [1:0] _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire [1:0] _EVAL_232;
  wire [1023:0] _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire  _EVAL_237;
  wire  _EVAL_238;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_205 = _EVAL_2 == 3'h6;
  assign _EVAL_32 = _EVAL_119 & _EVAL_46;
  assign _EVAL_208 = ~_EVAL_70;
  assign _EVAL_162 = _EVAL_0 <= 2'h2;
  assign _EVAL_176 = _EVAL_4 ^ 26'h2000000;
  assign _EVAL_123 = _EVAL_158 & _EVAL_189;
  assign _EVAL_164 = _EVAL_9 == _EVAL_69;
  assign _EVAL_190 = ~_EVAL_160;
  assign _EVAL_18 = _EVAL_5 == _EVAL_197;
  assign _EVAL_16 = _EVAL_7 & _EVAL_49;
  assign _EVAL_149 = _EVAL_194 >> _EVAL_1;
  assign _EVAL_170 = ~_EVAL_198;
  assign _EVAL_173 = _EVAL_91 | _EVAL_14;
  assign _EVAL_15 = _EVAL_1 <= 10'h23f;
  assign _EVAL_104 = _EVAL_6 & _EVAL_130;
  assign _EVAL_202 = _EVAL_158 & _EVAL_229;
  assign _EVAL_234 = _EVAL_5 <= 3'h3;
  assign _EVAL_56 = _EVAL_0[0];
  assign _EVAL_64 = _EVAL_92;
  assign _EVAL_53 = 2'h1 << _EVAL_56;
  assign _EVAL_40 = ~_EVAL_166;
  assign _EVAL_112 = _EVAL_116 & _EVAL_110;
  assign _EVAL_111 = _EVAL_97[1:0];
  assign _EVAL_97 = 5'h3 << _EVAL_0;
  assign _EVAL_43 = ~_EVAL_173;
  assign _EVAL_142 = ~_EVAL;
  assign _EVAL_27 = _EVAL_116 & _EVAL_123;
  assign _EVAL_157 = _EVAL_52 & _EVAL_132;
  assign _EVAL_33 = _EVAL_7 & _EVAL_212;
  assign _EVAL_209 = ~_EVAL_186;
  assign _EVAL_218 = _EVAL_7 & _EVAL_106;
  assign _EVAL_174 = _EVAL_171 | _EVAL_204;
  assign _EVAL_221 = _EVAL_200 | _EVAL_14;
  assign _EVAL_73 = _EVAL_11 == _EVAL_166;
  assign _EVAL_91 = _EVAL_15 & _EVAL_127;
  assign _EVAL_116 = _EVAL_66[0];
  assign _EVAL_76 = ~_EVAL_59;
  assign _EVAL_67 = _EVAL_12 == 3'h7;
  assign _EVAL_90 = _EVAL_217 | _EVAL_14;
  assign _EVAL_95 = ~_EVAL_111;
  assign _EVAL_89 = ~_EVAL_145;
  assign _EVAL_34 = _EVAL_85 | _EVAL_14;
  assign _EVAL_171 = _EVAL_93 | _EVAL_161;
  assign _EVAL_105 = _EVAL_134 == 4'h0;
  assign _EVAL_106 = _EVAL_12 == 3'h6;
  assign _EVAL_219 = ~_EVAL_14;
  assign _EVAL_50 = _EVAL_7 & _EVAL_199;
  assign _EVAL_212 = ~_EVAL_230;
  assign _EVAL_179 = _EVAL_151 | _EVAL_14;
  assign _EVAL_133 = ~_EVAL_37;
  assign _EVAL_124 = _EVAL_4 & _EVAL_61;
  assign _EVAL_99 = _EVAL_215 | _EVAL_214;
  assign _EVAL_193 = _EVAL_32 & _EVAL_216;
  assign _EVAL_163 = ~_EVAL_125;
  assign _EVAL_46 = ~_EVAL_23;
  assign _EVAL_216 = ~_EVAL_205;
  assign _EVAL_63 = _EVAL_149[0];
  assign _EVAL_214 = _EVAL_116 & _EVAL_184;
  assign _EVAL_21 = _EVAL_224[575:0];
  assign _EVAL_37 = _EVAL_15 | _EVAL_14;
  assign _EVAL_107 = _EVAL_168[0];
  assign _EVAL_54 = ~_EVAL_144;
  assign _EVAL_19 = _EVAL_12 == _EVAL_82;
  assign _EVAL_25 = _EVAL_6 & _EVAL_87;
  assign _EVAL_156 = _EVAL_7 & _EVAL_81;
  assign _EVAL_45 = _EVAL_177 | _EVAL_14;
  assign _EVAL_128 = _EVAL_11 & _EVAL_40;
  assign _EVAL_52 = _EVAL_66[1];
  assign _EVAL_155 = _EVAL_139 + 32'h1;
  assign _EVAL_29 = _EVAL_6 & _EVAL_205;
  assign _EVAL_84 = _EVAL_98 | _EVAL_14;
  assign _EVAL_38 = $signed(_EVAL_64) == 27'sh0;
  assign _EVAL_136 = _EVAL_211 | _EVAL_14;
  assign _EVAL_98 = _EVAL_0 == _EVAL_228;
  assign _EVAL_210 = ~_EVAL_179;
  assign _EVAL_114 = _EVAL_155[31:0];
  assign _EVAL_143 = _EVAL_152 & _EVAL_220;
  assign _EVAL_204 = _EVAL_139 < plusarg_reader_out;
  assign _EVAL_225 = ~_EVAL_20;
  assign _EVAL_119 = _EVAL_10 & _EVAL_6;
  assign _EVAL_222 = _EVAL_23 - 1'h1;
  assign _EVAL_113 = _EVAL_4 == _EVAL_72;
  assign _EVAL_121 = ~_EVAL_60;
  assign _EVAL_70 = ~_EVAL_75;
  assign _EVAL_57 = _EVAL_73 | _EVAL_14;
  assign _EVAL_80 = _EVAL_2 == _EVAL_226;
  assign _EVAL_184 = _EVAL_132 & _EVAL_229;
  assign _EVAL_66 = _EVAL_53 | 2'h1;
  assign _EVAL_93 = ~_EVAL_169;
  assign _EVAL_196 = _EVAL_167 & _EVAL_230;
  assign _EVAL_238 = _EVAL_7 & _EVAL_183;
  assign _EVAL_217 = _EVAL_13 == _EVAL_31;
  assign _EVAL_22 = ~_EVAL_35;
  assign _EVAL_153 = _EVAL_5 <= 3'h4;
  assign _EVAL_203 = _EVAL_19 | _EVAL_14;
  assign _EVAL_131 = ~_EVAL_45;
  assign _EVAL_189 = _EVAL_4[0];
  assign _EVAL_231 = ~_EVAL_71;
  assign _EVAL_39 = ~_EVAL_203;
  assign _EVAL_232 = _EVAL_188 - 1'h1;
  assign _EVAL_44 = ~_EVAL_221;
  assign _EVAL_103 = ~_EVAL_150;
  assign _EVAL_92 = $signed(_EVAL_137) & -27'sh10000;
  assign _EVAL_135 = _EVAL_192 | _EVAL_27;
  assign _EVAL_42 = _EVAL_52 & _EVAL_158;
  assign _EVAL_20 = _EVAL_78 | _EVAL_14;
  assign _EVAL_30 = _EVAL_5 <= 3'h1;
  assign _EVAL_167 = _EVAL_8 & _EVAL_7;
  assign _EVAL_159 = _EVAL_6 & _EVAL_180;
  assign _EVAL_168 = _EVAL_75 - 1'h1;
  assign _EVAL_224 = _EVAL_193 ? _EVAL_108 : 1024'h0;
  assign _EVAL_81 = _EVAL_12 == 3'h3;
  assign _EVAL_154 = _EVAL_167 & _EVAL_163;
  assign _EVAL_74 = _EVAL_6 & _EVAL_146;
  assign _EVAL_166 = {_EVAL_135,_EVAL_141,_EVAL_17,_EVAL_99};
  assign _EVAL_59 = _EVAL_55 | _EVAL_14;
  assign _EVAL_148 = ~_EVAL_62;
  assign _EVAL_145 = _EVAL_153 | _EVAL_14;
  assign _EVAL_185 = _EVAL_234 | _EVAL_14;
  assign _EVAL_83 = _EVAL_13 >= 2'h2;
  assign _EVAL_187 = ~_EVAL_136;
  assign _EVAL_71 = _EVAL_101 | _EVAL_14;
  assign _EVAL_199 = _EVAL_12 == 3'h1;
  assign _EVAL_129 = 1024'h1 << _EVAL_1;
  assign _EVAL_102 = _EVAL_116 & _EVAL_202;
  assign _EVAL_141 = _EVAL_192 | _EVAL_102;
  assign _EVAL_236 = _EVAL_7 & _EVAL_67;
  assign _EVAL_213 = _EVAL_222[0];
  assign _EVAL_130 = _EVAL_2 == 3'h0;
  assign _EVAL_144 = _EVAL_83 | _EVAL_14;
  assign _EVAL_165 = ~_EVAL_235;
  assign _EVAL_211 = _EVAL_128 == 4'h0;
  assign _EVAL_134 = ~_EVAL_11;
  assign _EVAL_227 = _EVAL_88 | _EVAL_194;
  assign _EVAL_58 = _EVAL_9 <= 10'h23f;
  assign _EVAL_65 = _EVAL_12 == 3'h2;
  assign _EVAL_100 = _EVAL_174 | _EVAL_14;
  assign _EVAL_77 = _EVAL_227 >> _EVAL_9;
  assign _EVAL_51 = ~_EVAL_96;
  assign _EVAL_132 = ~_EVAL_158;
  assign _EVAL_96 = _EVAL_105 | _EVAL_14;
  assign _EVAL_233 = _EVAL_154 ? _EVAL_129 : 1024'h0;
  assign _EVAL_140 = ~_EVAL_84;
  assign _EVAL_41 = ~_EVAL_57;
  assign _EVAL_215 = _EVAL_85 | _EVAL_157;
  assign _EVAL_169 = |_EVAL_194;
  assign _EVAL_191 = _EVAL_232[0];
  assign _EVAL_78 = _EVAL_1 == _EVAL_178;
  assign _EVAL_146 = _EVAL_2 == 3'h2;
  assign _EVAL_28 = _EVAL_7 & _EVAL_65;
  assign _EVAL_138 = _EVAL_7 & _EVAL_201;
  assign _EVAL_230 = ~_EVAL_188;
  assign _EVAL_223 = ~_EVAL_185;
  assign _EVAL_117 = _EVAL_6 & _EVAL_208;
  assign _EVAL_61 = {{24'd0}, _EVAL_95};
  assign _EVAL_198 = _EVAL_113 | _EVAL_14;
  assign _EVAL_118 = _EVAL_119 & _EVAL_70;
  assign _EVAL_201 = _EVAL_12 == 3'h5;
  assign _EVAL_55 = _EVAL_5 == 3'h0;
  assign _EVAL_160 = _EVAL_30 | _EVAL_14;
  assign _EVAL_172 = ~_EVAL_63;
  assign _EVAL_180 = _EVAL_2 == 3'h1;
  assign _EVAL_150 = _EVAL_18 | _EVAL_14;
  assign _EVAL_47 = ~_EVAL_90;
  assign _EVAL_110 = _EVAL_132 & _EVAL_189;
  assign _EVAL_237 = _EVAL_120 | _EVAL_14;
  assign _EVAL_151 = _EVAL_5 != 3'h0;
  assign _EVAL_183 = _EVAL_12 == 3'h4;
  assign _EVAL_161 = plusarg_reader_out == 32'h0;
  assign _EVAL_175 = _EVAL_79[0];
  assign _EVAL_115 = ~_EVAL_34;
  assign _EVAL_88 = _EVAL_233[575:0];
  assign _EVAL_87 = _EVAL_2 == 3'h4;
  assign _EVAL_62 = _EVAL_142 | _EVAL_14;
  assign _EVAL_200 = _EVAL_124 == 26'h0;
  assign _EVAL_181 = _EVAL_6 & _EVAL_147;
  assign _EVAL_35 = _EVAL_80 | _EVAL_14;
  assign _EVAL_158 = _EVAL_4[1];
  assign _EVAL_147 = _EVAL_2 == 3'h5;
  assign _EVAL_26 = _EVAL_167 | _EVAL_119;
  assign _EVAL_49 = _EVAL_12 == 3'h0;
  assign _EVAL_101 = _EVAL_77[0];
  assign _EVAL_152 = _EVAL_194 | _EVAL_88;
  assign _EVAL_192 = _EVAL_85 | _EVAL_42;
  assign _EVAL_85 = _EVAL_0 >= 2'h2;
  assign _EVAL_206 = ~_EVAL_237;
  assign _EVAL_186 = _EVAL_127 | _EVAL_14;
  assign _EVAL_79 = _EVAL_125 - 1'h1;
  assign _EVAL_177 = _EVAL_2 <= 3'h6;
  assign _EVAL_60 = _EVAL_172 | _EVAL_14;
  assign _EVAL_120 = _EVAL_5 <= 3'h2;
  assign _EVAL_36 = ~_EVAL_100;
  assign _EVAL_17 = _EVAL_215 | _EVAL_112;
  assign _EVAL_182 = ~_EVAL_86;
  assign _EVAL_220 = ~_EVAL_21;
  assign _EVAL_229 = ~_EVAL_189;
  assign _EVAL_235 = _EVAL_58 | _EVAL_14;
  assign _EVAL_86 = _EVAL_164 | _EVAL_14;
  assign _EVAL_127 = _EVAL_162 & _EVAL_38;
  assign _EVAL_137 = {1'b0,$signed(_EVAL_176)};
  assign _EVAL_108 = 1024'h1 << _EVAL_9;
  always @(posedge _EVAL_3) begin
    if (_EVAL_14) begin
      _EVAL_23 <= 1'h0;
    end else if (_EVAL_119) begin
      if (_EVAL_46) begin
        _EVAL_23 <= 1'h0;
      end else begin
        _EVAL_23 <= _EVAL_213;
      end
    end
    if (_EVAL_118) begin
      _EVAL_31 <= _EVAL_13;
    end
    if (_EVAL_118) begin
      _EVAL_69 <= _EVAL_9;
    end
    if (_EVAL_196) begin
      _EVAL_72 <= _EVAL_4;
    end
    if (_EVAL_14) begin
      _EVAL_75 <= 1'h0;
    end else if (_EVAL_119) begin
      if (_EVAL_70) begin
        _EVAL_75 <= 1'h0;
      end else begin
        _EVAL_75 <= _EVAL_107;
      end
    end
    if (_EVAL_196) begin
      _EVAL_82 <= _EVAL_12;
    end
    if (_EVAL_14) begin
      _EVAL_125 <= 1'h0;
    end else if (_EVAL_167) begin
      if (_EVAL_163) begin
        _EVAL_125 <= 1'h0;
      end else begin
        _EVAL_125 <= _EVAL_175;
      end
    end
    if (_EVAL_14) begin
      _EVAL_139 <= 32'h0;
    end else if (_EVAL_26) begin
      _EVAL_139 <= 32'h0;
    end else begin
      _EVAL_139 <= _EVAL_114;
    end
    if (_EVAL_196) begin
      _EVAL_178 <= _EVAL_1;
    end
    if (_EVAL_14) begin
      _EVAL_188 <= 1'h0;
    end else if (_EVAL_167) begin
      if (_EVAL_230) begin
        _EVAL_188 <= 1'h0;
      end else begin
        _EVAL_188 <= _EVAL_191;
      end
    end
    if (_EVAL_14) begin
      _EVAL_194 <= 576'h0;
    end else begin
      _EVAL_194 <= _EVAL_143;
    end
    if (_EVAL_196) begin
      _EVAL_197 <= _EVAL_5;
    end
    if (_EVAL_118) begin
      _EVAL_226 <= _EVAL_2;
    end
    if (_EVAL_196) begin
      _EVAL_228 <= _EVAL_0;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff03b96d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67393d85)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_36) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12bb7e04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c1c62f90)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_223) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6391a00d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44cd83b4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_187) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_182) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f0c87bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fc625f7c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_225) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6472ab5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(712963c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(11b2514a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_36) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(900d76f6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_131) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b348c45f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_187) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e0c19a2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(44291095)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_140) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dbc96655)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0feae33)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c3a8ca7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_43) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c93adc3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1509da2b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(460cf432)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(615992a3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45d3ef8d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_210) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3ffa5b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(73ddfdb5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(942bd67f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(abc3a8aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2119dca1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(709394b6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_89) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f8e107b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fbdee4e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8ff2157e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8832ba21)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_29 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_206) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8d7cf8e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4b4905af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1c11fdf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7f44432c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd28062c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_51) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(311cfd24)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20ebc132)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(67e7e8f9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(36f7126d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_47) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(711ffd6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7575cbe0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3bd7eca)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_210) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_22) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_43) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6309e185)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e3a8052)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_115) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_121) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(37c7b0e4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a42d0fe6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_51) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_206) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5dbea378)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_6 & _EVAL_131) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62f58504)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_22) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6a48f487)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2148839)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_133) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8954e04)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_140) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(79a6686)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_74 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2c0dcc0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_182) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_25 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(febb75af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6d4030cc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f1c11fdf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9d82fee1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_159 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7aad7aa0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(778771ec)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_39) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_170) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_104 & _EVAL_165) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_16 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_121) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_209) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edd25195)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_148) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3530c6ee)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e4986459)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_115) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(19544ee7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_76) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f7ec811)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_165) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c5d0a05)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_133) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_89) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_47) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f14e9299)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_156 & _EVAL_219) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_181 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fe97f546)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_138 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_44) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2f123877)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_236 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_28 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_39) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(95f85006)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_218 & _EVAL_148) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_33 & _EVAL_170) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fa4afa00)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_44) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(13e67033)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_219) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20439fdc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_50 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_76) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_238 & _EVAL_209) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_23 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_31 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_69 = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_72 = _RAND_3[25:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_75 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_82 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_125 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_139 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_178 = _RAND_8[9:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_188 = _RAND_9[0:0];
  _RAND_10 = {18{`RANDOM}};
  _EVAL_194 = _RAND_10[575:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_197 = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_226 = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_228 = _RAND_13[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
