//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_155_assert(
  input        _EVAL,
  input        _EVAL_0,
  input  [2:0] _EVAL_1,
  input        _EVAL_2,
  input        _EVAL_3,
  input        _EVAL_4,
  input  [6:0] _EVAL_5,
  input        _EVAL_6,
  input  [2:0] _EVAL_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_8;
  wire  _EVAL_9;
  reg [6:0] _EVAL_10;
  wire  _EVAL_11;
  wire  _EVAL_12;
  wire  _EVAL_13;
  wire  _EVAL_14;
  wire  _EVAL_15;
  wire  _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire [1:0] _EVAL_19;
  wire  _EVAL_21;
  reg  _EVAL_22;
  reg [2:0] _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire  _EVAL_26;
  wire  _EVAL_27;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire  _EVAL_31;
  wire  _EVAL_32;
  reg  _EVAL_33;
  wire  _EVAL_34;
  wire [7:0] _EVAL_35;
  wire  _EVAL_36;
  wire [1:0] _EVAL_37;
  reg  _EVAL_38;
  wire [7:0] _EVAL_39;
  wire [32:0] _EVAL_40;
  wire  _EVAL_41;
  reg  _EVAL_42;
  wire  _EVAL_43;
  reg [2:0] _EVAL_44;
  wire [6:0] _EVAL_45;
  wire [7:0] _EVAL_46;
  wire  _EVAL_47;
  wire [1:0] _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire [6:0] _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire [7:0] _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire  _EVAL_63;
  wire [31:0] _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire [1:0] _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  reg  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  reg [31:0] _EVAL_83;
  wire  _EVAL_84;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire [7:0] _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire [1:0] _EVAL_96;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire  _EVAL_103;
  wire [7:0] _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire [1:0] _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire [6:0] _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_118;
  wire  _EVAL_119;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_106 = ~_EVAL_42;
  assign _EVAL_48 = _EVAL_42 - 1'h1;
  assign _EVAL_114 = _EVAL_6 & _EVAL_66;
  assign _EVAL_80 = _EVAL_7 == _EVAL_23;
  assign _EVAL_12 = _EVAL_6 & _EVAL_21;
  assign _EVAL_118 = ~_EVAL_34;
  assign _EVAL_18 = _EVAL_83 < plusarg_reader_out;
  assign _EVAL_24 = _EVAL_7 == 3'h1;
  assign _EVAL_93 = $signed(_EVAL_104) == 8'sh0;
  assign _EVAL_65 = _EVAL & _EVAL_61;
  assign _EVAL_36 = _EVAL_7 == 3'h0;
  assign _EVAL_81 = _EVAL_96[0];
  assign _EVAL_110 = _EVAL_33 - 1'h1;
  assign _EVAL_98 = _EVAL_102 & _EVAL_47;
  assign _EVAL_79 = _EVAL_108 | _EVAL_11;
  assign _EVAL_108 = ~_EVAL_38;
  assign _EVAL_96 = _EVAL_98 ? 2'h1 : 2'h0;
  assign _EVAL_69 = _EVAL_6 & _EVAL_13;
  assign _EVAL_26 = ~_EVAL_106;
  assign _EVAL_32 = _EVAL_6 & _EVAL_36;
  assign _EVAL_102 = _EVAL_2 & _EVAL_6;
  assign _EVAL_45 = _EVAL_5 & 7'h3;
  assign _EVAL_54 = ~_EVAL_86;
  assign _EVAL_21 = _EVAL_7 == 3'h4;
  assign _EVAL_105 = _EVAL_6 & _EVAL_26;
  assign _EVAL_107 = _EVAL_6 & _EVAL_76;
  assign _EVAL_13 = _EVAL_7 == 3'h3;
  assign _EVAL_100 = ~_EVAL_33;
  assign _EVAL_75 = _EVAL_5 == _EVAL_10;
  assign _EVAL_82 = _EVAL_89 | _EVAL_11;
  assign _EVAL_109 = plusarg_reader_out == 32'h0;
  assign _EVAL_112 = _EVAL_52 | _EVAL_11;
  assign _EVAL_99 = _EVAL_6 & _EVAL_24;
  assign _EVAL_119 = _EVAL_19[0];
  assign _EVAL_11 = _EVAL_0;
  assign _EVAL_14 = _EVAL_1 == 3'h6;
  assign _EVAL_19 = _EVAL_72 - 1'h1;
  assign _EVAL_71 = ~_EVAL_111;
  assign _EVAL_39 = $signed(_EVAL_91) & -8'sh8;
  assign _EVAL_111 = _EVAL_80 | _EVAL_11;
  assign _EVAL_31 = _EVAL_38 | _EVAL_81;
  assign _EVAL_17 = ~_EVAL_97;
  assign _EVAL_84 = $signed(_EVAL_58) == 8'sh0;
  assign _EVAL_15 = _EVAL_95 & _EVAL_92;
  assign _EVAL_90 = _EVAL_6 & _EVAL_57;
  assign _EVAL_41 = _EVAL_110[0];
  assign _EVAL_16 = ~_EVAL_79;
  assign _EVAL_49 = _EVAL_4 & _EVAL;
  assign _EVAL_73 = _EVAL & _EVAL_62;
  assign _EVAL_101 = ~_EVAL_55;
  assign _EVAL_76 = _EVAL_7 == 3'h5;
  assign _EVAL_59 = _EVAL_50 | _EVAL_11;
  assign _EVAL_34 = _EVAL_75 | _EVAL_11;
  assign _EVAL_77 = ~_EVAL_8;
  assign _EVAL_64 = _EVAL_40[31:0];
  assign _EVAL_35 = {1'b0,$signed(_EVAL_51)};
  assign _EVAL_62 = _EVAL_1 == 3'h5;
  assign _EVAL_88 = _EVAL_1 == _EVAL_44;
  assign _EVAL_68 = _EVAL_22 - 1'h1;
  assign _EVAL_37 = _EVAL_15 ? 2'h1 : 2'h0;
  assign _EVAL_87 = _EVAL_60 | _EVAL_11;
  assign _EVAL_116 = ~_EVAL_59;
  assign _EVAL_53 = _EVAL_6 & _EVAL_30;
  assign _EVAL_67 = _EVAL_48[0];
  assign _EVAL_74 = _EVAL_102 & _EVAL_106;
  assign _EVAL_55 = ~_EVAL_22;
  assign _EVAL_63 = _EVAL_1 <= 3'h6;
  assign _EVAL_46 = $signed(_EVAL_35) & -8'shc;
  assign _EVAL_104 = _EVAL_46;
  assign _EVAL_89 = _EVAL_81 | _EVAL_38;
  assign _EVAL_78 = _EVAL_115 | _EVAL_109;
  assign _EVAL_40 = _EVAL_83 + 32'h1;
  assign _EVAL_115 = ~_EVAL_70;
  assign _EVAL_25 = _EVAL_68[0];
  assign _EVAL_50 = _EVAL_93 | _EVAL_84;
  assign _EVAL_29 = ~_EVAL_11;
  assign _EVAL_94 = ~_EVAL_87;
  assign _EVAL_47 = ~_EVAL_72;
  assign _EVAL_103 = ~_EVAL_112;
  assign _EVAL_95 = _EVAL_49 & _EVAL_100;
  assign _EVAL_66 = _EVAL_7 == 3'h6;
  assign _EVAL_56 = ~_EVAL_82;
  assign _EVAL_30 = _EVAL_7 == 3'h7;
  assign _EVAL_43 = _EVAL_49 & _EVAL_55;
  assign _EVAL_61 = _EVAL_1 == 3'h4;
  assign _EVAL_97 = _EVAL_37[0];
  assign _EVAL_86 = _EVAL_88 | _EVAL_11;
  assign _EVAL_58 = _EVAL_39;
  assign _EVAL_60 = _EVAL_78 | _EVAL_18;
  assign _EVAL_70 = |_EVAL_38;
  assign _EVAL_9 = _EVAL_102 | _EVAL_49;
  assign _EVAL_91 = {1'b0,$signed(_EVAL_113)};
  assign _EVAL_8 = _EVAL_63 | _EVAL_11;
  assign _EVAL_113 = _EVAL_5 ^ 7'h50;
  assign _EVAL_51 = _EVAL_5 ^ 7'h40;
  assign _EVAL_92 = ~_EVAL_14;
  assign _EVAL_27 = _EVAL & _EVAL_101;
  assign _EVAL_52 = _EVAL_45 == 7'h0;
  assign _EVAL_57 = _EVAL_7 == 3'h2;
  always @(posedge _EVAL_3) begin
    if (_EVAL_74) begin
      _EVAL_10 <= _EVAL_5;
    end
    if (_EVAL_74) begin
      _EVAL_23 <= _EVAL_7;
    end
    if (_EVAL_43) begin
      _EVAL_44 <= _EVAL_1;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_54) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7226c730)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f70a43d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(312625c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_16) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c3795348)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e12bfcdb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2f93b23)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fdfff19a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_27 & _EVAL_54) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8e12b9e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL & _EVAL_77) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c6c6e0c9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(de5b8fa9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_12 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a052a45)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c19b3e1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_73 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1ee44c89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c8b27308)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(58edd98d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(17d44d08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_71) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(566611c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_98 & _EVAL_16) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_15 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_12 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(94e7109)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6dfeb592)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_118) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(89213bde)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_90 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ff4c92fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac81bc9b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4f70a43d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(18b7f5b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_12 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_12 & _EVAL_116) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_99 & _EVAL_116) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cad3381e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_118) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b2927a7d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(84e2aca9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9844c3df)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_114 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_105 & _EVAL_71) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ab7b37c8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL & _EVAL_77) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_53 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_69 & _EVAL_103) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_32 & _EVAL_103) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a4ec6ef4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge _EVAL_3 or posedge _EVAL_0) begin
    if (_EVAL_0) begin
      _EVAL_22 <= 1'h0;
    end else if (_EVAL_49) begin
      if (_EVAL_55) begin
        _EVAL_22 <= 1'h0;
      end else begin
        _EVAL_22 <= _EVAL_25;
      end
    end
  end
  always @(posedge _EVAL_3 or posedge _EVAL_0) begin
    if (_EVAL_0) begin
      _EVAL_33 <= 1'h0;
    end else if (_EVAL_49) begin
      if (_EVAL_100) begin
        _EVAL_33 <= 1'h0;
      end else begin
        _EVAL_33 <= _EVAL_41;
      end
    end
  end
  always @(posedge _EVAL_3 or posedge _EVAL_0) begin
    if (_EVAL_0) begin
      _EVAL_38 <= 1'h0;
    end else begin
      _EVAL_38 <= _EVAL_31 & _EVAL_17;
    end
  end
  always @(posedge _EVAL_3 or posedge _EVAL_0) begin
    if (_EVAL_0) begin
      _EVAL_42 <= 1'h0;
    end else if (_EVAL_102) begin
      if (_EVAL_106) begin
        _EVAL_42 <= 1'h0;
      end else begin
        _EVAL_42 <= _EVAL_67;
      end
    end
  end
  always @(posedge _EVAL_3 or posedge _EVAL_0) begin
    if (_EVAL_0) begin
      _EVAL_72 <= 1'h0;
    end else if (_EVAL_102) begin
      if (_EVAL_47) begin
        _EVAL_72 <= 1'h0;
      end else begin
        _EVAL_72 <= _EVAL_119;
      end
    end
  end
  always @(posedge _EVAL_3 or posedge _EVAL_0) begin
    if (_EVAL_0) begin
      _EVAL_83 <= 32'h0;
    end else if (_EVAL_9) begin
      _EVAL_83 <= 32'h0;
    end else begin
      _EVAL_83 <= _EVAL_64;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_10 = _RAND_0[6:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_22 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_23 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_33 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_38 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_42 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_44 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_72 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_83 = _RAND_8[31:0];
`endif // RANDOMIZE_REG_INIT
  if (_EVAL_0) begin
    _EVAL_22 = 1'h0;
  end
  if (_EVAL_0) begin
    _EVAL_33 = 1'h0;
  end
  if (_EVAL_0) begin
    _EVAL_38 = 1'h0;
  end
  if (_EVAL_0) begin
    _EVAL_42 = 1'h0;
  end
  if (_EVAL_0) begin
    _EVAL_72 = 1'h0;
  end
  if (_EVAL_0) begin
    _EVAL_83 = 32'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
