//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_88(
  output [2:0]  _EVAL,
  input         _EVAL_0,
  output        _EVAL_1,
  input         _EVAL_2,
  output [2:0]  _EVAL_3,
  input  [2:0]  _EVAL_4,
  input  [31:0] _EVAL_5,
  input  [2:0]  _EVAL_6,
  output [3:0]  _EVAL_7,
  input  [29:0] _EVAL_8,
  input         _EVAL_9,
  output        _EVAL_10,
  output [29:0] _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  output        _EVAL_15,
  output        _EVAL_16,
  input         _EVAL_17,
  output [31:0] _EVAL_18,
  output        _EVAL_19,
  output [2:0]  _EVAL_20,
  input  [3:0]  _EVAL_21,
  input  [4:0]  _EVAL_22,
  input  [31:0] _EVAL_23,
  input         _EVAL_24,
  input         _EVAL_25,
  output [4:0]  _EVAL_26,
  output        _EVAL_27,
  output [1:0]  _EVAL_28,
  output [31:0] _EVAL_29,
  input         _EVAL_30,
  output [1:0]  _EVAL_31,
  input  [2:0]  _EVAL_32,
  input         _EVAL_33
);
  wire [2:0] _EVAL_34;
  wire  _EVAL_35;
  wire  _EVAL_36;
  wire [31:0] _EVAL_37;
  wire  _EVAL_38;
  wire [31:0] _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire [2:0] _EVAL_42;
  wire  _EVAL_43;
  wire [2:0] _EVAL_44;
  wire [2:0] _EVAL_45;
  wire  _EVAL_46;
  wire [2:0] _EVAL_47;
  wire [4:0] _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  wire [1:0] _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire [2:0] _EVAL_55;
  wire [2:0] _EVAL_56;
  wire  _EVAL_57;
  wire [2:0] _EVAL_58;
  wire [31:0] _EVAL_59;
  wire [2:0] _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire [3:0] _EVAL_63;
  wire [2:0] _EVAL_64;
  wire  _EVAL_65;
  wire [4:0] _EVAL_66;
  wire  _EVAL_67;
  wire [2:0] _EVAL_68;
  wire [29:0] _EVAL_69;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire [4:0] _EVAL_72;
  wire [1:0] _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire [29:0] _EVAL_77;
  wire  _EVAL_78;
  wire [31:0] _EVAL_79;
  wire  fragmenter__EVAL;
  wire  fragmenter__EVAL_0;
  wire  fragmenter__EVAL_1;
  wire [1:0] fragmenter__EVAL_2;
  wire  fragmenter__EVAL_3;
  wire  fragmenter__EVAL_4;
  wire [2:0] fragmenter__EVAL_5;
  wire  fragmenter__EVAL_6;
  wire [31:0] fragmenter__EVAL_7;
  wire [4:0] fragmenter__EVAL_8;
  wire [29:0] fragmenter__EVAL_9;
  wire  fragmenter__EVAL_10;
  wire [2:0] fragmenter__EVAL_11;
  wire [3:0] fragmenter__EVAL_12;
  wire [3:0] fragmenter__EVAL_13;
  wire [29:0] fragmenter__EVAL_14;
  wire [31:0] fragmenter__EVAL_15;
  wire  fragmenter__EVAL_16;
  wire [1:0] fragmenter__EVAL_17;
  wire  fragmenter__EVAL_18;
  wire  fragmenter__EVAL_19;
  wire [9:0] fragmenter__EVAL_20;
  wire [2:0] fragmenter__EVAL_21;
  wire [2:0] fragmenter__EVAL_22;
  wire [9:0] fragmenter__EVAL_23;
  wire  fragmenter__EVAL_24;
  wire  fragmenter__EVAL_25;
  wire  fragmenter__EVAL_26;
  wire [4:0] fragmenter__EVAL_27;
  wire  fragmenter__EVAL_28;
  wire  fragmenter__EVAL_29;
  wire  fragmenter__EVAL_30;
  wire [1:0] fragmenter__EVAL_31;
  wire  fragmenter__EVAL_32;
  wire [1:0] fragmenter__EVAL_33;
  wire [2:0] fragmenter__EVAL_34;
  wire  fragmenter__EVAL_35;
  wire [31:0] fragmenter__EVAL_36;
  wire [2:0] fragmenter__EVAL_37;
  wire  fragmenter__EVAL_38;
  wire  fragmenter__EVAL_39;
  wire  fragmenter__EVAL_40;
  wire [31:0] fragmenter__EVAL_41;
  wire  fragmenter__EVAL_42;
  wire [2:0] fragmenter__EVAL_43;
  wire  fragmenter__EVAL_44;
  wire [2:0] fragmenter__EVAL_45;
  wire  fragmenter__EVAL_46;
  wire  fragmenter__EVAL_47;
  wire  fragmenter__EVAL_48;
  wire  _EVAL_80;
  wire [4:0] _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire [4:0] _EVAL_85;
  wire [3:0] _EVAL_86;
  wire [31:0] _EVAL_87;
  wire [1:0] _EVAL_88;
  wire [29:0] _EVAL_89;
  wire  _EVAL_90;
  wire [1:0] _EVAL_91;
  wire [2:0] _EVAL_92;
  wire [31:0] _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire [9:0] buffer__EVAL;
  wire  buffer__EVAL_0;
  wire [1:0] buffer__EVAL_1;
  wire  buffer__EVAL_2;
  wire  buffer__EVAL_3;
  wire [1:0] buffer__EVAL_4;
  wire  buffer__EVAL_5;
  wire  buffer__EVAL_6;
  wire  buffer__EVAL_7;
  wire [2:0] buffer__EVAL_8;
  wire [2:0] buffer__EVAL_9;
  wire [2:0] buffer__EVAL_10;
  wire [9:0] buffer__EVAL_11;
  wire  buffer__EVAL_12;
  wire [1:0] buffer__EVAL_13;
  wire  buffer__EVAL_14;
  wire  buffer__EVAL_15;
  wire [2:0] buffer__EVAL_16;
  wire [31:0] buffer__EVAL_17;
  wire [31:0] buffer__EVAL_18;
  wire [1:0] buffer__EVAL_19;
  wire [2:0] buffer__EVAL_20;
  wire  buffer__EVAL_21;
  wire [3:0] buffer__EVAL_22;
  wire  buffer__EVAL_23;
  wire [9:0] buffer__EVAL_24;
  wire [29:0] buffer__EVAL_25;
  wire [31:0] buffer__EVAL_26;
  wire  buffer__EVAL_27;
  wire  buffer__EVAL_28;
  wire  buffer__EVAL_29;
  wire  buffer__EVAL_30;
  wire [3:0] buffer__EVAL_31;
  wire  buffer__EVAL_32;
  wire  buffer__EVAL_33;
  wire  buffer__EVAL_34;
  wire [31:0] buffer__EVAL_35;
  wire  buffer__EVAL_36;
  wire [1:0] buffer__EVAL_37;
  wire [2:0] buffer__EVAL_38;
  wire  buffer__EVAL_39;
  wire [1:0] buffer__EVAL_40;
  wire  buffer__EVAL_41;
  wire  buffer__EVAL_42;
  wire [29:0] buffer__EVAL_43;
  wire [9:0] buffer__EVAL_44;
  wire  buffer__EVAL_45;
  wire  buffer__EVAL_46;
  wire  buffer__EVAL_47;
  wire  buffer__EVAL_48;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire [31:0] tl2ahb__EVAL;
  wire  tl2ahb__EVAL_0;
  wire [9:0] tl2ahb__EVAL_1;
  wire  tl2ahb__EVAL_2;
  wire [31:0] tl2ahb__EVAL_3;
  wire  tl2ahb__EVAL_4;
  wire  tl2ahb__EVAL_5;
  wire  tl2ahb__EVAL_6;
  wire  tl2ahb__EVAL_7;
  wire [1:0] tl2ahb__EVAL_8;
  wire  tl2ahb__EVAL_9;
  wire  tl2ahb__EVAL_10;
  wire [9:0] tl2ahb__EVAL_11;
  wire [29:0] tl2ahb__EVAL_12;
  wire [1:0] tl2ahb__EVAL_13;
  wire  tl2ahb__EVAL_14;
  wire  tl2ahb__EVAL_15;
  wire [2:0] tl2ahb__EVAL_16;
  wire [1:0] tl2ahb__EVAL_17;
  wire [31:0] tl2ahb__EVAL_18;
  wire [3:0] tl2ahb__EVAL_19;
  wire [2:0] tl2ahb__EVAL_20;
  wire [1:0] tl2ahb__EVAL_21;
  wire  tl2ahb__EVAL_22;
  wire [3:0] tl2ahb__EVAL_23;
  wire  tl2ahb__EVAL_24;
  wire  tl2ahb__EVAL_25;
  wire [31:0] tl2ahb__EVAL_26;
  wire [29:0] tl2ahb__EVAL_27;
  wire  tl2ahb__EVAL_28;
  wire  tl2ahb__EVAL_29;
  wire [2:0] tl2ahb__EVAL_30;
  wire  tl2ahb__EVAL_31;
  wire  tl2ahb__EVAL_32;
  wire [2:0] tl2ahb__EVAL_33;
  wire [2:0] _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire [29:0] _EVAL_103;
  wire [3:0] _EVAL_104;
  wire [31:0] _EVAL_105;
  wire [3:0] _EVAL_106;
  wire [2:0] _EVAL_107;
  wire [4:0] _EVAL_108;
  wire [2:0] _EVAL_109;
  wire [4:0] _EVAL_110;
  wire [4:0] _EVAL_111;
  wire  _EVAL_112;
  wire [2:0] _EVAL_113;
  wire [31:0] _EVAL_114;
  wire  _EVAL_115;
  wire [2:0] _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire [2:0] _EVAL_123;
  wire [2:0] _EVAL_124;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire [2:0] _EVAL_129;
  _EVAL_87 fragmenter (
    ._EVAL(fragmenter__EVAL),
    ._EVAL_0(fragmenter__EVAL_0),
    ._EVAL_1(fragmenter__EVAL_1),
    ._EVAL_2(fragmenter__EVAL_2),
    ._EVAL_3(fragmenter__EVAL_3),
    ._EVAL_4(fragmenter__EVAL_4),
    ._EVAL_5(fragmenter__EVAL_5),
    ._EVAL_6(fragmenter__EVAL_6),
    ._EVAL_7(fragmenter__EVAL_7),
    ._EVAL_8(fragmenter__EVAL_8),
    ._EVAL_9(fragmenter__EVAL_9),
    ._EVAL_10(fragmenter__EVAL_10),
    ._EVAL_11(fragmenter__EVAL_11),
    ._EVAL_12(fragmenter__EVAL_12),
    ._EVAL_13(fragmenter__EVAL_13),
    ._EVAL_14(fragmenter__EVAL_14),
    ._EVAL_15(fragmenter__EVAL_15),
    ._EVAL_16(fragmenter__EVAL_16),
    ._EVAL_17(fragmenter__EVAL_17),
    ._EVAL_18(fragmenter__EVAL_18),
    ._EVAL_19(fragmenter__EVAL_19),
    ._EVAL_20(fragmenter__EVAL_20),
    ._EVAL_21(fragmenter__EVAL_21),
    ._EVAL_22(fragmenter__EVAL_22),
    ._EVAL_23(fragmenter__EVAL_23),
    ._EVAL_24(fragmenter__EVAL_24),
    ._EVAL_25(fragmenter__EVAL_25),
    ._EVAL_26(fragmenter__EVAL_26),
    ._EVAL_27(fragmenter__EVAL_27),
    ._EVAL_28(fragmenter__EVAL_28),
    ._EVAL_29(fragmenter__EVAL_29),
    ._EVAL_30(fragmenter__EVAL_30),
    ._EVAL_31(fragmenter__EVAL_31),
    ._EVAL_32(fragmenter__EVAL_32),
    ._EVAL_33(fragmenter__EVAL_33),
    ._EVAL_34(fragmenter__EVAL_34),
    ._EVAL_35(fragmenter__EVAL_35),
    ._EVAL_36(fragmenter__EVAL_36),
    ._EVAL_37(fragmenter__EVAL_37),
    ._EVAL_38(fragmenter__EVAL_38),
    ._EVAL_39(fragmenter__EVAL_39),
    ._EVAL_40(fragmenter__EVAL_40),
    ._EVAL_41(fragmenter__EVAL_41),
    ._EVAL_42(fragmenter__EVAL_42),
    ._EVAL_43(fragmenter__EVAL_43),
    ._EVAL_44(fragmenter__EVAL_44),
    ._EVAL_45(fragmenter__EVAL_45),
    ._EVAL_46(fragmenter__EVAL_46),
    ._EVAL_47(fragmenter__EVAL_47),
    ._EVAL_48(fragmenter__EVAL_48)
  );
  _EVAL_84 buffer (
    ._EVAL(buffer__EVAL),
    ._EVAL_0(buffer__EVAL_0),
    ._EVAL_1(buffer__EVAL_1),
    ._EVAL_2(buffer__EVAL_2),
    ._EVAL_3(buffer__EVAL_3),
    ._EVAL_4(buffer__EVAL_4),
    ._EVAL_5(buffer__EVAL_5),
    ._EVAL_6(buffer__EVAL_6),
    ._EVAL_7(buffer__EVAL_7),
    ._EVAL_8(buffer__EVAL_8),
    ._EVAL_9(buffer__EVAL_9),
    ._EVAL_10(buffer__EVAL_10),
    ._EVAL_11(buffer__EVAL_11),
    ._EVAL_12(buffer__EVAL_12),
    ._EVAL_13(buffer__EVAL_13),
    ._EVAL_14(buffer__EVAL_14),
    ._EVAL_15(buffer__EVAL_15),
    ._EVAL_16(buffer__EVAL_16),
    ._EVAL_17(buffer__EVAL_17),
    ._EVAL_18(buffer__EVAL_18),
    ._EVAL_19(buffer__EVAL_19),
    ._EVAL_20(buffer__EVAL_20),
    ._EVAL_21(buffer__EVAL_21),
    ._EVAL_22(buffer__EVAL_22),
    ._EVAL_23(buffer__EVAL_23),
    ._EVAL_24(buffer__EVAL_24),
    ._EVAL_25(buffer__EVAL_25),
    ._EVAL_26(buffer__EVAL_26),
    ._EVAL_27(buffer__EVAL_27),
    ._EVAL_28(buffer__EVAL_28),
    ._EVAL_29(buffer__EVAL_29),
    ._EVAL_30(buffer__EVAL_30),
    ._EVAL_31(buffer__EVAL_31),
    ._EVAL_32(buffer__EVAL_32),
    ._EVAL_33(buffer__EVAL_33),
    ._EVAL_34(buffer__EVAL_34),
    ._EVAL_35(buffer__EVAL_35),
    ._EVAL_36(buffer__EVAL_36),
    ._EVAL_37(buffer__EVAL_37),
    ._EVAL_38(buffer__EVAL_38),
    ._EVAL_39(buffer__EVAL_39),
    ._EVAL_40(buffer__EVAL_40),
    ._EVAL_41(buffer__EVAL_41),
    ._EVAL_42(buffer__EVAL_42),
    ._EVAL_43(buffer__EVAL_43),
    ._EVAL_44(buffer__EVAL_44),
    ._EVAL_45(buffer__EVAL_45),
    ._EVAL_46(buffer__EVAL_46),
    ._EVAL_47(buffer__EVAL_47),
    ._EVAL_48(buffer__EVAL_48)
  );
  _EVAL_80 tl2ahb (
    ._EVAL(tl2ahb__EVAL),
    ._EVAL_0(tl2ahb__EVAL_0),
    ._EVAL_1(tl2ahb__EVAL_1),
    ._EVAL_2(tl2ahb__EVAL_2),
    ._EVAL_3(tl2ahb__EVAL_3),
    ._EVAL_4(tl2ahb__EVAL_4),
    ._EVAL_5(tl2ahb__EVAL_5),
    ._EVAL_6(tl2ahb__EVAL_6),
    ._EVAL_7(tl2ahb__EVAL_7),
    ._EVAL_8(tl2ahb__EVAL_8),
    ._EVAL_9(tl2ahb__EVAL_9),
    ._EVAL_10(tl2ahb__EVAL_10),
    ._EVAL_11(tl2ahb__EVAL_11),
    ._EVAL_12(tl2ahb__EVAL_12),
    ._EVAL_13(tl2ahb__EVAL_13),
    ._EVAL_14(tl2ahb__EVAL_14),
    ._EVAL_15(tl2ahb__EVAL_15),
    ._EVAL_16(tl2ahb__EVAL_16),
    ._EVAL_17(tl2ahb__EVAL_17),
    ._EVAL_18(tl2ahb__EVAL_18),
    ._EVAL_19(tl2ahb__EVAL_19),
    ._EVAL_20(tl2ahb__EVAL_20),
    ._EVAL_21(tl2ahb__EVAL_21),
    ._EVAL_22(tl2ahb__EVAL_22),
    ._EVAL_23(tl2ahb__EVAL_23),
    ._EVAL_24(tl2ahb__EVAL_24),
    ._EVAL_25(tl2ahb__EVAL_25),
    ._EVAL_26(tl2ahb__EVAL_26),
    ._EVAL_27(tl2ahb__EVAL_27),
    ._EVAL_28(tl2ahb__EVAL_28),
    ._EVAL_29(tl2ahb__EVAL_29),
    ._EVAL_30(tl2ahb__EVAL_30),
    ._EVAL_31(tl2ahb__EVAL_31),
    ._EVAL_32(tl2ahb__EVAL_32),
    ._EVAL_33(tl2ahb__EVAL_33)
  );
  assign _EVAL_45 = fragmenter__EVAL_11;
  assign _EVAL_76 = fragmenter__EVAL_32;
  assign _EVAL_106 = _EVAL_63;
  assign _EVAL_71 = _EVAL_127;
  assign fragmenter__EVAL_24 = _EVAL_36;
  assign fragmenter__EVAL_8 = _EVAL_108;
  assign _EVAL_52 = _EVAL_88;
  assign _EVAL_53 = fragmenter__EVAL_4;
  assign _EVAL_35 = _EVAL_40;
  assign _EVAL_43 = _EVAL_95;
  assign fragmenter__EVAL_33 = buffer__EVAL_4;
  assign _EVAL_123 = _EVAL_92;
  assign _EVAL_63 = _EVAL_21;
  assign _EVAL_119 = _EVAL_38;
  assign _EVAL_129 = _EVAL_55;
  assign _EVAL_29 = tl2ahb__EVAL_3;
  assign _EVAL_117 = _EVAL_112;
  assign fragmenter__EVAL_48 = _EVAL_67;
  assign tl2ahb__EVAL_28 = buffer__EVAL_23;
  assign tl2ahb__EVAL_32 = buffer__EVAL_46;
  assign tl2ahb__EVAL_15 = _EVAL_13;
  assign fragmenter__EVAL_10 = _EVAL_33;
  assign _EVAL_16 = _EVAL_94;
  assign buffer__EVAL_2 = tl2ahb__EVAL_24;
  assign buffer__EVAL_30 = _EVAL_2;
  assign _EVAL_125 = _EVAL_51;
  assign _EVAL_103 = _EVAL_89;
  assign tl2ahb__EVAL_27 = buffer__EVAL_43;
  assign buffer__EVAL_3 = tl2ahb__EVAL_4;
  assign fragmenter__EVAL_0 = buffer__EVAL_21;
  assign _EVAL_91 = _EVAL_73;
  assign _EVAL_105 = _EVAL_114;
  assign _EVAL_127 = _EVAL_12;
  assign fragmenter__EVAL_40 = buffer__EVAL_28;
  assign buffer__EVAL_15 = fragmenter__EVAL_1;
  assign _EVAL_48 = _EVAL_110;
  assign _EVAL_89 = _EVAL_77;
  assign _EVAL_93 = _EVAL_79;
  assign fragmenter__EVAL_19 = buffer__EVAL_32;
  assign _EVAL_95 = _EVAL_53;
  assign fragmenter__EVAL_45 = _EVAL_64;
  assign _EVAL_1 = _EVAL_70;
  assign fragmenter__EVAL_44 = _EVAL_2;
  assign tl2ahb__EVAL_19 = buffer__EVAL_31;
  assign _EVAL_42 = _EVAL_123;
  assign _EVAL_46 = _EVAL_71;
  assign _EVAL_118 = _EVAL_43;
  assign _EVAL_82 = _EVAL_125;
  assign _EVAL_44 = _EVAL_6;
  assign _EVAL_61 = _EVAL_101;
  assign tl2ahb__EVAL_30 = buffer__EVAL_8;
  assign tl2ahb__EVAL_22 = buffer__EVAL_12;
  assign _EVAL_88 = _EVAL_91;
  assign fragmenter__EVAL_17 = buffer__EVAL_19;
  assign _EVAL_67 = _EVAL_46;
  assign fragmenter__EVAL_30 = _EVAL_57;
  assign fragmenter__EVAL_39 = buffer__EVAL_48;
  assign _EVAL_108 = _EVAL_48;
  assign fragmenter__EVAL_29 = buffer__EVAL_29;
  assign _EVAL_73 = fragmenter__EVAL_2;
  assign fragmenter__EVAL_42 = _EVAL_49;
  assign _EVAL_85 = _EVAL_72;
  assign _EVAL_39 = _EVAL_105;
  assign _EVAL_87 = _EVAL_93;
  assign buffer__EVAL_37 = fragmenter__EVAL_31;
  assign buffer__EVAL_22 = fragmenter__EVAL_13;
  assign _EVAL_124 = _EVAL_98;
  assign fragmenter__EVAL_9 = _EVAL_69;
  assign _EVAL_3 = _EVAL_68;
  assign _EVAL_15 = _EVAL_84;
  assign _EVAL_126 = _EVAL_119;
  assign _EVAL_62 = fragmenter__EVAL_25;
  assign tl2ahb__EVAL_11 = buffer__EVAL_44;
  assign _EVAL_100 = _EVAL_102;
  assign _EVAL_69 = _EVAL_103;
  assign fragmenter__EVAL_35 = _EVAL_97;
  assign buffer__EVAL_24 = fragmenter__EVAL_23;
  assign tl2ahb__EVAL_29 = _EVAL_2;
  assign _EVAL_50 = _EVAL_62;
  assign _EVAL_80 = _EVAL_90;
  assign _EVAL_75 = _EVAL_65;
  assign _EVAL_83 = _EVAL_80;
  assign _EVAL_92 = _EVAL_107;
  assign _EVAL_27 = _EVAL_126;
  assign _EVAL_81 = _EVAL_85;
  assign _EVAL_70 = _EVAL_99;
  assign _EVAL_90 = _EVAL_14;
  assign _EVAL_84 = _EVAL_78;
  assign _EVAL_121 = _EVAL_128;
  assign _EVAL_86 = _EVAL_104;
  assign _EVAL_107 = _EVAL_4;
  assign fragmenter__EVAL_15 = buffer__EVAL_17;
  assign tl2ahb__EVAL_21 = buffer__EVAL_13;
  assign fragmenter__EVAL_12 = _EVAL_86;
  assign _EVAL_101 = fragmenter__EVAL_6;
  assign buffer__EVAL_5 = tl2ahb__EVAL_31;
  assign buffer__EVAL_1 = tl2ahb__EVAL_8;
  assign _EVAL_110 = _EVAL_111;
  assign _EVAL_7 = tl2ahb__EVAL_23;
  assign buffer__EVAL_47 = fragmenter__EVAL;
  assign _EVAL_57 = _EVAL_41;
  assign _EVAL_78 = _EVAL_50;
  assign _EVAL_64 = _EVAL_124;
  assign buffer__EVAL_38 = fragmenter__EVAL_22;
  assign tl2ahb__EVAL_5 = buffer__EVAL_0;
  assign _EVAL_11 = tl2ahb__EVAL_12;
  assign tl2ahb__EVAL_18 = buffer__EVAL_35;
  assign _EVAL_36 = _EVAL_75;
  assign _EVAL_122 = _EVAL_96;
  assign buffer__EVAL_25 = fragmenter__EVAL_14;
  assign tl2ahb__EVAL_7 = _EVAL_33;
  assign buffer__EVAL_18 = tl2ahb__EVAL;
  assign buffer__EVAL = tl2ahb__EVAL_1;
  assign _EVAL_109 = _EVAL_113;
  assign _EVAL_120 = _EVAL_117;
  assign _EVAL_31 = _EVAL_52;
  assign _EVAL_59 = _EVAL_87;
  assign fragmenter__EVAL_26 = _EVAL_35;
  assign _EVAL_114 = _EVAL_23;
  assign _EVAL_47 = _EVAL_116;
  assign _EVAL_49 = _EVAL_122;
  assign _EVAL_116 = _EVAL_34;
  assign buffer__EVAL_33 = tl2ahb__EVAL_25;
  assign _EVAL_55 = fragmenter__EVAL_5;
  assign _EVAL_104 = _EVAL_106;
  assign _EVAL_98 = _EVAL_44;
  assign buffer__EVAL_36 = _EVAL_33;
  assign tl2ahb__EVAL_26 = _EVAL_5;
  assign _EVAL_96 = _EVAL_74;
  assign tl2ahb__EVAL_6 = buffer__EVAL_45;
  assign _EVAL_28 = tl2ahb__EVAL_13;
  assign fragmenter__EVAL_38 = _EVAL_115;
  assign _EVAL_99 = _EVAL_61;
  assign fragmenter__EVAL_20 = buffer__EVAL_11;
  assign tl2ahb__EVAL_2 = buffer__EVAL_6;
  assign _EVAL_68 = _EVAL_56;
  assign _EVAL_20 = tl2ahb__EVAL_20;
  assign buffer__EVAL_14 = fragmenter__EVAL_3;
  assign fragmenter__EVAL_43 = _EVAL_42;
  assign buffer__EVAL_41 = fragmenter__EVAL_18;
  assign _EVAL_40 = _EVAL_121;
  assign _EVAL_56 = _EVAL_129;
  assign _EVAL_112 = _EVAL_25;
  assign _EVAL_72 = _EVAL_66;
  assign _EVAL_77 = _EVAL_8;
  assign _EVAL_19 = _EVAL_118;
  assign buffer__EVAL_39 = fragmenter__EVAL_16;
  assign _EVAL_41 = _EVAL_100;
  assign _EVAL_128 = _EVAL_24;
  assign _EVAL_51 = fragmenter__EVAL_28;
  assign _EVAL_97 = _EVAL_120;
  assign buffer__EVAL_7 = tl2ahb__EVAL_0;
  assign _EVAL_37 = _EVAL_39;
  assign _EVAL = _EVAL_47;
  assign buffer__EVAL_34 = fragmenter__EVAL_46;
  assign _EVAL_38 = _EVAL_76;
  assign _EVAL_10 = tl2ahb__EVAL_10;
  assign _EVAL_113 = _EVAL_58;
  assign _EVAL_65 = _EVAL_54;
  assign _EVAL_66 = fragmenter__EVAL_27;
  assign buffer__EVAL_20 = fragmenter__EVAL_34;
  assign _EVAL_111 = _EVAL_22;
  assign _EVAL_18 = _EVAL_59;
  assign _EVAL_115 = _EVAL_83;
  assign buffer__EVAL_26 = fragmenter__EVAL_7;
  assign _EVAL_102 = _EVAL_30;
  assign buffer__EVAL_27 = fragmenter__EVAL_47;
  assign buffer__EVAL_9 = tl2ahb__EVAL_33;
  assign tl2ahb__EVAL_16 = buffer__EVAL_10;
  assign fragmenter__EVAL_36 = _EVAL_37;
  assign tl2ahb__EVAL_9 = buffer__EVAL_42;
  assign _EVAL_58 = _EVAL_32;
  assign _EVAL_54 = _EVAL_9;
  assign fragmenter__EVAL_21 = buffer__EVAL_16;
  assign tl2ahb__EVAL_14 = _EVAL_0;
  assign buffer__EVAL_40 = tl2ahb__EVAL_17;
  assign _EVAL_79 = fragmenter__EVAL_41;
  assign _EVAL_34 = _EVAL_45;
  assign fragmenter__EVAL_37 = _EVAL_60;
  assign _EVAL_74 = _EVAL_17;
  assign _EVAL_60 = _EVAL_109;
  assign _EVAL_26 = _EVAL_81;
  assign _EVAL_94 = _EVAL_82;
endmodule
