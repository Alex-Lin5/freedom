//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_111(
  output        _EVAL,
  input         _EVAL_0,
  output        _EVAL_1,
  input         _EVAL_2,
  output        _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  output        _EVAL_6,
  input  [31:0] _EVAL_7,
  input  [3:0]  _EVAL_8,
  output [1:0]  _EVAL_9,
  input         _EVAL_10,
  input  [10:0] _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  output [31:0] _EVAL_14,
  output [31:0] _EVAL_15,
  output        _EVAL_16,
  input         _EVAL_17,
  input         _EVAL_18,
  input         _EVAL_19,
  input  [1:0]  _EVAL_20,
  output        _EVAL_21,
  input         _EVAL_22,
  output        _EVAL_23,
  input  [24:0] _EVAL_24,
  output        _EVAL_25,
  input  [3:0]  _EVAL_26,
  output [31:0] _EVAL_27,
  input  [2:0]  _EVAL_28,
  output [10:0] _EVAL_29,
  input  [31:0] _EVAL_30,
  input  [2:0]  _EVAL_31,
  input  [31:0] _EVAL_32,
  input  [31:0] _EVAL_33,
  input         _EVAL_34,
  output        _EVAL_35,
  input  [31:0] _EVAL_36,
  output [2:0]  _EVAL_37
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [255:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
`endif // RANDOMIZE_REG_INIT
  reg  _EVAL_38;
  reg  _EVAL_41;
  wire [255:0] _EVAL_43;
  reg  _EVAL_44;
  wire  _EVAL_45;
  wire [7:0] _EVAL_46;
  wire [255:0] _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_51;
  wire  _EVAL_52;
  wire [31:0] _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_58;
  wire [31:0] _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_62;
  wire [6:0] _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire [7:0] _EVAL_68;
  wire  _EVAL_70;
  wire  _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire [7:0] _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_83;
  wire  _EVAL_84;
  reg  _EVAL_85;
  wire [10:0] _EVAL_86;
  wire  _EVAL_87;
  wire [31:0] _EVAL_90;
  reg  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire [10:0] _EVAL_95;
  wire [255:0] _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  reg  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_103;
  wire [10:0] _EVAL_104;
  wire  _EVAL_105;
  wire [255:0] _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_109;
  reg [31:0] _EVAL_111;
  reg  _EVAL_112;
  wire  _EVAL_113;
  wire [6:0] tag_array__EVAL;
  wire  tag_array__EVAL_0;
  wire [19:0] tag_array__EVAL_1;
  wire [19:0] tag_array__EVAL_2;
  wire [19:0] tag_array__EVAL_3;
  wire  tag_array__EVAL_4;
  wire [19:0] tag_array__EVAL_5;
  wire  tag_array__EVAL_6;
  wire  tag_array__EVAL_7;
  wire  tag_array__EVAL_8;
  wire  _EVAL_114;
  wire [7:0] _EVAL_116;
  wire  _EVAL_117;
  wire [10:0] _EVAL_119;
  wire [7:0] _EVAL_121;
  wire  _EVAL_122;
  wire [31:0] _EVAL_123;
  wire  _EVAL_125;
  wire  _EVAL_126;
  wire  _EVAL_130;
  reg [5:0] _EVAL_132;
  wire  _EVAL_133;
  wire [7:0] _EVAL_137;
  wire  _EVAL_138;
  wire [10:0] _EVAL_140;
  wire  _EVAL_142;
  wire [31:0] _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_147;
  wire [7:0] _EVAL_151;
  reg  _EVAL_153;
  wire [5:0] _EVAL_154;
  wire [7:0] _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_161;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire [7:0] _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  reg  _EVAL_168;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire [7:0] _EVAL_172;
  wire  _EVAL_173;
  reg [31:0] _EVAL_174;
  wire [7:0] _EVAL_176;
  wire  _EVAL_177;
  reg  _EVAL_178;
  wire [7:0] _EVAL_179;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire  _EVAL_184;
  wire [18:0] _EVAL_185;
  wire [1:0] _EVAL_186;
  wire [31:0] _EVAL_187;
  wire  _EVAL_188;
  wire [7:0] _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire  _EVAL_192;
  wire  _EVAL_193;
  wire [31:0] _EVAL_194;
  reg [31:0] _EVAL_195;
  wire [7:0] _EVAL_196;
  wire  _EVAL_197;
  wire [255:0] _EVAL_198;
  wire  _EVAL_200;
  wire [18:0] _EVAL_202;
  reg [2:0] _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  reg [10:0] _EVAL_206;
  wire [31:0] _EVAL_207;
  wire [10:0] _EVAL_208;
  wire  _EVAL_211;
  reg  _EVAL_212;
  reg  _EVAL_214;
  reg [255:0] _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  reg [3:0] _EVAL_218;
  wire [18:0] _EVAL_220;
  wire  _EVAL_221;
  wire  _EVAL_224;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire [6:0] _EVAL_230;
  wire  _EVAL_231;
  wire [6:0] _EVAL_232;
  wire  _EVAL_233;
  wire [7:0] _EVAL_234;
  wire  _EVAL_235;
  wire  _EVAL_236;
  wire [5:0] _EVAL_237;
  wire [10:0] _EVAL_238;
  wire [31:0] data_arrays_0__EVAL;
  wire  data_arrays_0__EVAL_0;
  wire [31:0] data_arrays_0__EVAL_1;
  wire [10:0] data_arrays_0__EVAL_2;
  wire  data_arrays_0__EVAL_3;
  wire  data_arrays_0__EVAL_4;
  wire [31:0] data_arrays_0__EVAL_5;
  wire [31:0] data_arrays_0__EVAL_6;
  wire  data_arrays_0__EVAL_7;
  wire  data_arrays_0__EVAL_8;
  wire [31:0] _EVAL_241;
  wire  _EVAL_242;
  wire [25:0] _EVAL_243;
  wire [255:0] _EVAL_244;
  reg  _EVAL_246;
  wire  _EVAL_247;
  wire [10:0] _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire [24:0] _EVAL_254;
  wire  _EVAL_256;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire [18:0] _EVAL_260;
  reg  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire [5:0] _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire [7:0] _EVAL_270;
  wire  _EVAL_272;
  wire [5:0] _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire [15:0] _EVAL_276;
  wire  _EVAL_278;
  reg  _EVAL_279;
  wire  _EVAL_281;
  wire  _EVAL_282;
  reg [31:0] _EVAL_285;
  wire  _EVAL_286;
  wire [255:0] _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  wire  _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_293;
  reg [13:0] _EVAL_294;
  wire [7:0] _EVAL_296;
  wire  _EVAL_298;
  wire  _EVAL_302;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_307;
  wire  _EVAL_308;
  wire  repl_way_v0_prng__EVAL;
  wire  repl_way_v0_prng__EVAL_0;
  wire  repl_way_v0_prng__EVAL_1;
  wire  repl_way_v0_prng__EVAL_2;
  wire  repl_way_v0_prng__EVAL_3;
  wire  repl_way_v0_prng__EVAL_4;
  wire  repl_way_v0_prng__EVAL_5;
  wire  repl_way_v0_prng__EVAL_6;
  wire  repl_way_v0_prng__EVAL_7;
  wire  repl_way_v0_prng__EVAL_8;
  wire  repl_way_v0_prng__EVAL_9;
  wire  repl_way_v0_prng__EVAL_10;
  wire  repl_way_v0_prng__EVAL_11;
  wire  repl_way_v0_prng__EVAL_12;
  wire  repl_way_v0_prng__EVAL_13;
  wire  repl_way_v0_prng__EVAL_14;
  wire  repl_way_v0_prng__EVAL_15;
  wire  repl_way_v0_prng__EVAL_16;
  wire  repl_way_v0_prng__EVAL_17;
  wire [7:0] _EVAL_309;
  wire [5:0] _EVAL_310;
  wire  _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_313;
  reg [1:0] _EVAL_314;
  reg [6:0] _EVAL_315;
  wire [22:0] _EVAL_317;
  wire  _EVAL_318;
  wire [6:0] _EVAL_319;
  wire [31:0] _EVAL_320;
  wire  _EVAL_321;
  _EVAL_208 tag_array (
    ._EVAL(tag_array__EVAL),
    ._EVAL_0(tag_array__EVAL_0),
    ._EVAL_1(tag_array__EVAL_1),
    ._EVAL_2(tag_array__EVAL_2),
    ._EVAL_3(tag_array__EVAL_3),
    ._EVAL_4(tag_array__EVAL_4),
    ._EVAL_5(tag_array__EVAL_5),
    ._EVAL_6(tag_array__EVAL_6),
    ._EVAL_7(tag_array__EVAL_7),
    ._EVAL_8(tag_array__EVAL_8)
  );
  _EVAL_209 data_arrays_0 (
    ._EVAL(data_arrays_0__EVAL),
    ._EVAL_0(data_arrays_0__EVAL_0),
    ._EVAL_1(data_arrays_0__EVAL_1),
    ._EVAL_2(data_arrays_0__EVAL_2),
    ._EVAL_3(data_arrays_0__EVAL_3),
    ._EVAL_4(data_arrays_0__EVAL_4),
    ._EVAL_5(data_arrays_0__EVAL_5),
    ._EVAL_6(data_arrays_0__EVAL_6),
    ._EVAL_7(data_arrays_0__EVAL_7),
    ._EVAL_8(data_arrays_0__EVAL_8)
  );
  _EVAL_106 repl_way_v0_prng (
    ._EVAL(repl_way_v0_prng__EVAL),
    ._EVAL_0(repl_way_v0_prng__EVAL_0),
    ._EVAL_1(repl_way_v0_prng__EVAL_1),
    ._EVAL_2(repl_way_v0_prng__EVAL_2),
    ._EVAL_3(repl_way_v0_prng__EVAL_3),
    ._EVAL_4(repl_way_v0_prng__EVAL_4),
    ._EVAL_5(repl_way_v0_prng__EVAL_5),
    ._EVAL_6(repl_way_v0_prng__EVAL_6),
    ._EVAL_7(repl_way_v0_prng__EVAL_7),
    ._EVAL_8(repl_way_v0_prng__EVAL_8),
    ._EVAL_9(repl_way_v0_prng__EVAL_9),
    ._EVAL_10(repl_way_v0_prng__EVAL_10),
    ._EVAL_11(repl_way_v0_prng__EVAL_11),
    ._EVAL_12(repl_way_v0_prng__EVAL_12),
    ._EVAL_13(repl_way_v0_prng__EVAL_13),
    ._EVAL_14(repl_way_v0_prng__EVAL_14),
    ._EVAL_15(repl_way_v0_prng__EVAL_15),
    ._EVAL_16(repl_way_v0_prng__EVAL_16),
    ._EVAL_17(repl_way_v0_prng__EVAL_17)
  );
  assign repl_way_v0_prng__EVAL_14 = _EVAL_34;
  assign _EVAL_144 = _EVAL_191 & _EVAL_91;
  assign _EVAL_302 = ~_EVAL_308;
  assign repl_way_v0_prng__EVAL_11 = _EVAL_17;
  assign _EVAL_211 = _EVAL_74 < 1'h1;
  assign _EVAL_250 = _EVAL_105 & _EVAL_109;
  assign _EVAL_259 = _EVAL_217 | _EVAL_72;
  assign _EVAL_97 = ~_EVAL_198;
  assign _EVAL_37 = _EVAL_51 ? 3'h0 : 3'h1;
  assign _EVAL_52 = _EVAL_41 & _EVAL_278;
  assign _EVAL_59 = data_arrays_0__EVAL_6;
  assign _EVAL_233 = _EVAL_66 | _EVAL_214;
  assign _EVAL_228 = _EVAL_18 | _EVAL_144;
  assign _EVAL_217 = _EVAL_132 == 6'h1;
  assign _EVAL_234 = _EVAL_143[23:16];
  assign _EVAL_104 = _EVAL_204 ? _EVAL_208 : _EVAL_249;
  assign _EVAL_196 = _EVAL_90[15:8];
  assign _EVAL_188 = _EVAL_235 & _EVAL_58;
  assign _EVAL_166 = _EVAL_30[13];
  assign _EVAL_142 = _EVAL_30 < 32'h1804000;
  assign _EVAL_133 = _EVAL_85 ? _EVAL_264 : _EVAL_321;
  assign _EVAL_272 = _EVAL_12 & _EVAL_161;
  assign _EVAL_198 = _EVAL_43 | _EVAL_287;
  assign _EVAL_235 = _EVAL_197 & _EVAL_117;
  assign _EVAL_101 = ~_EVAL_188;
  assign _EVAL_55 = ~_EVAL_288;
  assign _EVAL_47 = _EVAL_215 | _EVAL_287;
  assign _EVAL_87 = ~_EVAL_13;
  assign _EVAL_113 = _EVAL_262 & _EVAL_125;
  assign _EVAL_312 = tag_array__EVAL_3[19];
  assign _EVAL_173 = _EVAL_41 | _EVAL_85;
  assign _EVAL_35 = ~_EVAL_313;
  assign _EVAL_3 = ~_EVAL_214;
  assign _EVAL_290 = _EVAL_93 ? _EVAL_304 : _EVAL_22;
  assign _EVAL_177 = ~_EVAL_214;
  assign _EVAL_291 = _EVAL_77 <= _EVAL_296;
  assign _EVAL_296 = {{1'd0}, _EVAL_315};
  assign _EVAL_189 = {1'h1,_EVAL_232};
  assign _EVAL_90 = _EVAL_55 ? _EVAL_194 : _EVAL_174;
  assign data_arrays_0__EVAL_5 = _EVAL_214 ? _EVAL_174 : _EVAL_7;
  assign _EVAL_125 = _EVAL_165 <= _EVAL_296;
  assign _EVAL_140 = {_EVAL_230, 4'h0};
  assign _EVAL_267 = _EVAL_311 & _EVAL_60;
  assign _EVAL_220 = _EVAL_30[31:13];
  assign _EVAL_163 = _EVAL_256 | _EVAL_153;
  assign _EVAL_98 = _EVAL_214 ? _EVAL_49 : _EVAL_268;
  assign _EVAL_307 = ~_EVAL_166;
  assign _EVAL_319 = _EVAL_32[12:6];
  assign tag_array__EVAL_7 = ~_EVAL_268;
  assign _EVAL_170 = _EVAL_51 & _EVAL_164;
  assign _EVAL_54 = _EVAL_101 & _EVAL_200;
  assign _EVAL_172 = _EVAL_93 ? _EVAL_156 : {{1'd0}, _EVAL_315};
  assign tag_array__EVAL_2 = {_EVAL_228,_EVAL_260};
  assign _EVAL_182 = _EVAL_235 | _EVAL_204;
  assign _EVAL_70 = _EVAL_258 | _EVAL_269;
  assign _EVAL_254 = _EVAL_204 ? _EVAL_24 : {{11'd0}, _EVAL_294};
  assign _EVAL_186 = {_EVAL_250,_EVAL_114};
  assign _EVAL_158 = |_EVAL_186;
  assign _EVAL_64 = _EVAL_132 == 6'h0;
  assign _EVAL_145 = _EVAL_262 & _EVAL_226;
  assign _EVAL_230 = _EVAL_111[12:6];
  assign _EVAL_119 = _EVAL_214 ? _EVAL_86 : _EVAL_104;
  assign _EVAL_256 = _EVAL_227 | _EVAL_85;
  assign _EVAL_236 = ~_EVAL_170;
  assign _EVAL_273 = _EVAL_63[5:0];
  assign _EVAL_23 = ~_EVAL_308;
  assign _EVAL_260 = _EVAL_111[31:13];
  assign _EVAL_298 = _EVAL_188 & _EVAL_281;
  assign _EVAL_251 = &_EVAL_218;
  assign tag_array__EVAL_0 = _EVAL_54 | _EVAL_188;
  assign _EVAL_187 = _EVAL_178 ? _EVAL_285 : 32'h0;
  assign _EVAL_242 = _EVAL_203[2];
  assign _EVAL_231 = _EVAL_212 & _EVAL_84;
  assign _EVAL_252 = _EVAL_38 & _EVAL_79;
  assign _EVAL_317 = 23'hff << _EVAL_26;
  assign _EVAL_194 = _EVAL_187 | _EVAL_207;
  assign _EVAL_244 = _EVAL_215 >> _EVAL_189;
  assign _EVAL_275 = _EVAL_41 & _EVAL_305;
  assign _EVAL_126 = _EVAL_30 >= 32'h1800000;
  assign _EVAL_79 = ~_EVAL_19;
  assign _EVAL_25 = _EVAL_279;
  assign _EVAL_65 = _EVAL_262 & _EVAL_45;
  assign _EVAL_93 = ~_EVAL_130;
  assign _EVAL_83 = _EVAL_147 | _EVAL_212;
  assign _EVAL_321 = _EVAL_73 & _EVAL_307;
  assign tag_array__EVAL_6 = _EVAL_235 & _EVAL_58;
  assign _EVAL_311 = ~_EVAL_233;
  assign _EVAL_48 = _EVAL_202 == _EVAL_220;
  assign _EVAL_207 = _EVAL_100 ? _EVAL_195 : 32'h0;
  assign _EVAL_282 = _EVAL_107 | _EVAL_44;
  assign _EVAL_265 = _EVAL_270[7:2];
  assign _EVAL_86 = _EVAL_294[12:2];
  assign _EVAL_241 = {_EVAL_176,_EVAL_234,_EVAL_196,_EVAL_46};
  assign _EVAL_232 = _EVAL_30[12:6];
  assign _EVAL_258 = _EVAL_71 | _EVAL_105;
  assign _EVAL_289 = _EVAL_51 & _EVAL_263;
  assign _EVAL_45 = _EVAL_151 <= _EVAL_296;
  assign _EVAL_67 = _EVAL_106[0];
  assign _EVAL_109 = tag_array__EVAL_1[19];
  assign _EVAL_278 = ~_EVAL_2;
  assign _EVAL_72 = _EVAL_154 == 6'h0;
  assign _EVAL_95 = {{5'd0}, _EVAL_237};
  assign _EVAL_190 = ~_EVAL_10;
  assign _EVAL_270 = ~_EVAL_121;
  assign _EVAL_238 = _EVAL_140 | _EVAL_95;
  assign _EVAL_286 = _EVAL_218[1];
  assign data_arrays_0__EVAL_4 = _EVAL_214 ? _EVAL_49 : _EVAL_268;
  assign _EVAL_264 = _EVAL_145 & _EVAL_266;
  assign _EVAL_122 = _EVAL_221 | _EVAL_168;
  assign _EVAL_263 = _EVAL_218[2];
  assign _EVAL_84 = ~_EVAL_112;
  assign _EVAL_287 = 256'h1 << _EVAL_309;
  assign _EVAL_281 = ~_EVAL_44;
  assign _EVAL_58 = _EVAL_259 & _EVAL_197;
  assign _EVAL_114 = _EVAL_193 & _EVAL_312;
  assign _EVAL_60 = _EVAL_200 | _EVAL_204;
  assign _EVAL_1 = _EVAL_12 & _EVAL_161;
  assign _EVAL_164 = _EVAL_218[0];
  assign _EVAL_14 = {_EVAL_243, 6'h0};
  assign _EVAL_151 = _EVAL_24[13:6];
  assign _EVAL_221 = _EVAL_231 & _EVAL_87;
  assign _EVAL_9 = _EVAL_314;
  assign _EVAL_156 = _EVAL_80 ? _EVAL_151 : {{1'd0}, _EVAL_315};
  assign _EVAL_185 = tag_array__EVAL_1[18:0];
  assign tag_array__EVAL_8 = _EVAL_17;
  assign _EVAL_143 = _EVAL_184 ? _EVAL_194 : _EVAL_174;
  assign _EVAL_202 = tag_array__EVAL_3[18:0];
  assign _EVAL_107 = _EVAL_204 ? _EVAL_290 : _EVAL_22;
  assign _EVAL = _EVAL_221 & _EVAL_246;
  assign _EVAL_227 = _EVAL_4 | _EVAL_38;
  assign data_arrays_0__EVAL_8 = _EVAL_267 | _EVAL_233;
  assign _EVAL_293 = _EVAL_185 == _EVAL_220;
  assign _EVAL_208 = _EVAL_24[12:2];
  assign _EVAL_197 = _EVAL_177 & _EVAL_0;
  assign _EVAL_191 = _EVAL_237 > 6'h0;
  assign _EVAL_92 = _EVAL_138 & _EVAL_181;
  assign _EVAL_305 = ~_EVAL_122;
  assign _EVAL_117 = _EVAL_31[0];
  assign _EVAL_56 = _EVAL_218[3];
  assign _EVAL_266 = ~_EVAL_49;
  assign _EVAL_106 = _EVAL_215 >> _EVAL_116;
  assign data_arrays_0__EVAL = _EVAL_214 ? _EVAL_174 : _EVAL_7;
  assign _EVAL_205 = _EVAL_51 & _EVAL_56;
  assign data_arrays_0__EVAL_2 = _EVAL_235 ? _EVAL_238 : _EVAL_119;
  assign _EVAL_103 = _EVAL_94 | _EVAL_214;
  assign _EVAL_268 = _EVAL_274 | _EVAL_247;
  assign _EVAL_46 = _EVAL_53[7:0];
  assign _EVAL_247 = _EVAL_262 & _EVAL_291;
  assign _EVAL_94 = _EVAL_99 | _EVAL_153;
  assign _EVAL_15 = _EVAL_187 | _EVAL_207;
  assign _EVAL_276 = {repl_way_v0_prng__EVAL_6,repl_way_v0_prng__EVAL_8,repl_way_v0_prng__EVAL_13,repl_way_v0_prng__EVAL
    ,repl_way_v0_prng__EVAL_4,repl_way_v0_prng__EVAL_10,repl_way_v0_prng__EVAL_7,repl_way_v0_prng__EVAL_0,_EVAL_68};
  assign _EVAL_27 = _EVAL_174;
  assign _EVAL_29 = _EVAL_206;
  assign _EVAL_137 = _EVAL_294[13:6];
  assign _EVAL_161 = _EVAL_221 & _EVAL_246;
  assign _EVAL_81 = ~_EVAL_205;
  assign _EVAL_16 = _EVAL_83 | _EVAL_168;
  assign _EVAL_304 = _EVAL_80 | _EVAL_22;
  assign _EVAL_320 = data_arrays_0__EVAL_1;
  assign _EVAL_147 = _EVAL_318 | _EVAL_41;
  assign repl_way_v0_prng__EVAL_2 = _EVAL_12 & _EVAL_161;
  assign _EVAL_171 = _EVAL_272 | _EVAL_168;
  assign _EVAL_130 = _EVAL_28[2];
  assign _EVAL_192 = _EVAL_103 | _EVAL_38;
  assign _EVAL_116 = {1'h0,_EVAL_232};
  assign _EVAL_274 = _EVAL_276[0];
  assign _EVAL_237 = _EVAL_154 & _EVAL_310;
  assign _EVAL_62 = _EVAL_85 & _EVAL_167;
  assign _EVAL_51 = ~_EVAL_242;
  assign _EVAL_249 = _EVAL_32[12:2];
  assign data_arrays_0__EVAL_3 = _EVAL_17;
  assign _EVAL_309 = {_EVAL_268,_EVAL_230};
  assign tag_array__EVAL_5 = {_EVAL_228,_EVAL_260};
  assign data_arrays_0__EVAL_0 = _EVAL_66 | _EVAL_214;
  assign _EVAL_74 = _EVAL_24[13];
  assign _EVAL_71 = _EVAL_193 | _EVAL_133;
  assign _EVAL_105 = _EVAL_92 & _EVAL_293;
  assign _EVAL_165 = _EVAL_30[13:6];
  assign _EVAL_193 = _EVAL_78 & _EVAL_48;
  assign _EVAL_318 = _EVAL_163 | _EVAL_214;
  assign _EVAL_226 = _EVAL_137 <= _EVAL_296;
  assign _EVAL_68 = {repl_way_v0_prng__EVAL_15,repl_way_v0_prng__EVAL_17,repl_way_v0_prng__EVAL_16,
    repl_way_v0_prng__EVAL_3,repl_way_v0_prng__EVAL_12,repl_way_v0_prng__EVAL_1,repl_way_v0_prng__EVAL_5,
    repl_way_v0_prng__EVAL_9};
  assign _EVAL_204 = _EVAL_302 & _EVAL_4;
  assign _EVAL_216 = ~_EVAL_168;
  assign _EVAL_200 = _EVAL_35 & _EVAL_5;
  assign _EVAL_184 = ~_EVAL_289;
  assign _EVAL_78 = _EVAL_67 & _EVAL_181;
  assign _EVAL_49 = _EVAL_294[13];
  assign _EVAL_181 = ~_EVAL_85;
  assign data_arrays_0__EVAL_7 = ~_EVAL_98;
  assign _EVAL_138 = _EVAL_244[0];
  assign tag_array__EVAL = _EVAL_188 ? _EVAL_230 : _EVAL_319;
  assign _EVAL_99 = _EVAL_0 | _EVAL_85;
  assign _EVAL_73 = _EVAL_224 & _EVAL_113;
  assign _EVAL_243 = _EVAL_111[31:6];
  assign _EVAL_157 = _EVAL_153 | _EVAL_252;
  assign _EVAL_123 = _EVAL_81 ? _EVAL_194 : _EVAL_174;
  assign _EVAL_154 = _EVAL_117 ? _EVAL_265 : 6'h0;
  assign _EVAL_269 = _EVAL_85 | _EVAL_224;
  assign _EVAL_176 = _EVAL_123[31:24];
  assign _EVAL_313 = _EVAL_182 | _EVAL_214;
  assign _EVAL_308 = _EVAL_192 | _EVAL_190;
  assign _EVAL_121 = _EVAL_317[7:0];
  assign _EVAL_66 = _EVAL_235 & _EVAL_281;
  assign _EVAL_43 = ~_EVAL_215;
  assign _EVAL_179 = _EVAL_204 ? _EVAL_172 : {{1'd0}, _EVAL_315};
  assign _EVAL_224 = _EVAL_126 & _EVAL_142;
  assign _EVAL_167 = _EVAL_51 & _EVAL_251;
  assign _EVAL_53 = _EVAL_236 ? _EVAL_194 : _EVAL_174;
  assign tag_array__EVAL_4 = _EVAL_274 | _EVAL_247;
  assign _EVAL_63 = _EVAL_132 - 6'h1;
  assign _EVAL_80 = ~_EVAL_65;
  assign _EVAL_6 = _EVAL_38;
  assign _EVAL_77 = {_EVAL_274,_EVAL_230};
  assign _EVAL_288 = _EVAL_51 & _EVAL_286;
  assign _EVAL_21 = _EVAL_212 & _EVAL_112;
  assign _EVAL_310 = ~_EVAL_273;
  always @(posedge _EVAL_17) begin
    if (_EVAL_34) begin
      _EVAL_38 <= 1'h0;
    end else begin
      _EVAL_38 <= _EVAL_157;
    end
    if (_EVAL_34) begin
      _EVAL_41 <= 1'h0;
    end else begin
      _EVAL_41 <= _EVAL_200;
    end
    if (_EVAL_216) begin
      _EVAL_44 <= 1'h0;
    end else begin
      _EVAL_44 <= _EVAL_282;
    end
    if (_EVAL_34) begin
      _EVAL_85 <= 1'h0;
    end else begin
      _EVAL_85 <= _EVAL_204;
    end
    if (_EVAL_235) begin
      _EVAL_91 <= _EVAL_228;
    end
    if (_EVAL_173) begin
      if (_EVAL_62) begin
        _EVAL_100 <= 1'h0;
      end else begin
        _EVAL_100 <= _EVAL_105;
      end
    end
    if (_EVAL_275) begin
      _EVAL_111 <= _EVAL_30;
    end
    _EVAL_112 <= _EVAL_70;
    if (_EVAL_34) begin
      _EVAL_132 <= 6'h0;
    end else if (_EVAL_197) begin
      if (_EVAL_64) begin
        if (_EVAL_117) begin
          _EVAL_132 <= _EVAL_265;
        end else begin
          _EVAL_132 <= 6'h0;
        end
      end else begin
        _EVAL_132 <= _EVAL_273;
      end
    end
    if (_EVAL_34) begin
      _EVAL_153 <= 1'h0;
    end else begin
      _EVAL_153 <= _EVAL_85;
    end
    if (_EVAL_34) begin
      _EVAL_168 <= 1'h0;
    end else if (_EVAL_188) begin
      _EVAL_168 <= 1'h0;
    end else begin
      _EVAL_168 <= _EVAL_171;
    end
    if (_EVAL_153) begin
      _EVAL_174 <= _EVAL_241;
    end else if (_EVAL_204) begin
      _EVAL_174 <= _EVAL_33;
    end
    if (_EVAL_173) begin
      if (_EVAL_62) begin
        _EVAL_178 <= 1'h0;
      end else begin
        _EVAL_178 <= _EVAL_71;
      end
    end
    if (_EVAL_173) begin
      _EVAL_195 <= _EVAL_320;
    end
    if (_EVAL_204) begin
      _EVAL_203 <= _EVAL_28;
    end
    if (_EVAL_204) begin
      _EVAL_206 <= _EVAL_11;
    end
    if (_EVAL_34) begin
      _EVAL_212 <= 1'h0;
    end else begin
      _EVAL_212 <= _EVAL_52;
    end
    _EVAL_214 <= _EVAL_153 & _EVAL_51;
    if (_EVAL_34) begin
      _EVAL_215 <= 256'h0;
    end else if (_EVAL_107) begin
      _EVAL_215 <= 256'h0;
    end else if (_EVAL_235) begin
      if (_EVAL_298) begin
        _EVAL_215 <= _EVAL_47;
      end else begin
        _EVAL_215 <= _EVAL_97;
      end
    end
    if (_EVAL_204) begin
      _EVAL_218 <= _EVAL_8;
    end
    _EVAL_246 <= ~_EVAL_122;
    if (_EVAL_34) begin
      _EVAL_262 <= 1'h0;
    end else if (_EVAL_204) begin
      if (_EVAL_93) begin
        _EVAL_262 <= _EVAL_211;
      end
    end
    if (_EVAL_173) begin
      _EVAL_279 <= _EVAL_158;
    end
    if (_EVAL_173) begin
      _EVAL_285 <= _EVAL_59;
    end
    _EVAL_294 <= _EVAL_254[13:0];
    if (_EVAL_204) begin
      _EVAL_314 <= _EVAL_20;
    end
    _EVAL_315 <= _EVAL_179[6:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_38 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_41 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_44 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_85 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_91 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_100 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_111 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_112 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_132 = _RAND_8[5:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_153 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_168 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_174 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_178 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_195 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_203 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_206 = _RAND_15[10:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_212 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _EVAL_214 = _RAND_17[0:0];
  _RAND_18 = {8{`RANDOM}};
  _EVAL_215 = _RAND_18[255:0];
  _RAND_19 = {1{`RANDOM}};
  _EVAL_218 = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  _EVAL_246 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _EVAL_262 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  _EVAL_279 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  _EVAL_285 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  _EVAL_294 = _RAND_24[13:0];
  _RAND_25 = {1{`RANDOM}};
  _EVAL_314 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  _EVAL_315 = _RAND_26[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
