//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_36_assert(
  input         _EVAL,
  input  [2:0]  _EVAL_0,
  input         _EVAL_1,
  input  [3:0]  _EVAL_2,
  input  [3:0]  _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  input  [1:0]  _EVAL_6,
  input  [3:0]  _EVAL_7,
  input  [2:0]  _EVAL_8,
  input         _EVAL_9,
  input  [31:0] _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  wire [1:0] _EVAL_16;
  wire  _EVAL_17;
  wire  _EVAL_18;
  wire  _EVAL_19;
  wire  _EVAL_20;
  wire [32:0] _EVAL_21;
  wire  _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire  _EVAL_25;
  wire [32:0] _EVAL_26;
  wire  _EVAL_27;
  wire [3:0] _EVAL_28;
  wire  _EVAL_29;
  wire [32:0] _EVAL_30;
  wire  _EVAL_31;
  reg [1:0] _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  wire [32:0] _EVAL_35;
  wire [31:0] _EVAL_36;
  wire [32:0] _EVAL_37;
  wire  _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire  _EVAL_43;
  wire [32:0] _EVAL_44;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  reg  _EVAL_51;
  wire  _EVAL_52;
  wire [5:0] _EVAL_53;
  wire [32:0] _EVAL_54;
  wire [22:0] _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire [5:0] _EVAL_61;
  wire  _EVAL_63;
  wire  _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  reg [5:0] _EVAL_71;
  wire [6:0] _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire [6:0] _EVAL_75;
  wire  _EVAL_76;
  wire [31:0] _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire [32:0] _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire [7:0] _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire [32:0] _EVAL_88;
  wire  _EVAL_89;
  wire [22:0] _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  reg  _EVAL_100;
  wire  _EVAL_101;
  wire [32:0] _EVAL_102;
  wire  _EVAL_103;
  reg [5:0] _EVAL_104;
  wire [1:0] _EVAL_105;
  wire [31:0] _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  reg [31:0] _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire  _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  reg [2:0] _EVAL_125;
  wire  _EVAL_126;
  wire [32:0] _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  reg [2:0] _EVAL_132;
  wire  _EVAL_133;
  wire [5:0] _EVAL_134;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire  _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  reg [5:0] _EVAL_142;
  reg [31:0] _EVAL_143;
  wire [7:0] _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire [31:0] _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_151;
  wire [7:0] _EVAL_152;
  wire [31:0] _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire [5:0] _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire [6:0] _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire [32:0] _EVAL_170;
  wire  _EVAL_171;
  wire [32:0] _EVAL_172;
  reg [3:0] _EVAL_173;
  wire [32:0] _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire [7:0] _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire [32:0] _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire [32:0] _EVAL_186;
  wire  _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire [32:0] _EVAL_192;
  wire  _EVAL_193;
  wire  _EVAL_194;
  wire  _EVAL_195;
  wire  _EVAL_196;
  wire [31:0] _EVAL_197;
  wire  _EVAL_198;
  wire [31:0] _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire [3:0] _EVAL_208;
  wire [32:0] _EVAL_209;
  wire [31:0] _EVAL_210;
  wire [31:0] _EVAL_211;
  wire  _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  reg [3:0] _EVAL_219;
  reg [5:0] _EVAL_220;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire [1:0] _EVAL_227;
  wire [32:0] _EVAL_228;
  wire  _EVAL_229;
  wire  _EVAL_230;
  wire  _EVAL_231;
  wire  _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire [1:0] _EVAL_236;
  wire  _EVAL_237;
  wire [32:0] _EVAL_238;
  wire [32:0] _EVAL_239;
  wire  _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_243;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_248;
  wire  _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire [32:0] _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  reg  _EVAL_255;
  wire  _EVAL_256;
  wire  _EVAL_257;
  wire  _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_262;
  wire  _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  reg  _EVAL_270;
  wire [5:0] _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire  _EVAL_277;
  wire  _EVAL_278;
  wire  _EVAL_279;
  wire [3:0] _EVAL_280;
  wire [6:0] _EVAL_281;
  wire [3:0] _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  wire  _EVAL_285;
  wire  _EVAL_286;
  wire  _EVAL_287;
  wire  _EVAL_288;
  wire [31:0] _EVAL_289;
  wire  _EVAL_290;
  wire [1:0] _EVAL_291;
  wire  _EVAL_292;
  wire [32:0] _EVAL_293;
  wire [32:0] _EVAL_294;
  wire [5:0] _EVAL_295;
  wire  _EVAL_296;
  wire  _EVAL_297;
  wire [32:0] _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  wire  _EVAL_302;
  wire  _EVAL_304;
  wire  _EVAL_305;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_94 = _EVAL_260 | _EVAL_4;
  assign _EVAL_87 = ~_EVAL_86;
  assign _EVAL_154 = _EVAL_49 | _EVAL_118;
  assign _EVAL_101 = ~_EVAL_272;
  assign _EVAL_203 = _EVAL_0 == 3'h6;
  assign _EVAL_281 = _EVAL_71 - 6'h1;
  assign _EVAL_175 = $signed(_EVAL_170) & -33'sh2000;
  assign _EVAL_222 = _EVAL_300 & _EVAL_249;
  assign _EVAL_78 = ~_EVAL_4;
  assign _EVAL_52 = _EVAL_11 & _EVAL_141;
  assign _EVAL_304 = ~_EVAL_305;
  assign _EVAL_120 = _EVAL_97 | _EVAL_4;
  assign _EVAL_40 = _EVAL_169 & _EVAL_176;
  assign _EVAL_290 = ~_EVAL_155;
  assign _EVAL_107 = _EVAL_5 & _EVAL_121;
  assign _EVAL_246 = _EVAL_5 & _EVAL_226;
  assign _EVAL_30 = _EVAL_110 + 32'h1;
  assign _EVAL_230 = ~_EVAL_9;
  assign _EVAL_291 = _EVAL_105 | 2'h1;
  assign _EVAL_192 = _EVAL_81;
  assign _EVAL_28 = {_EVAL_23,_EVAL_189,_EVAL_278,_EVAL_301};
  assign _EVAL_258 = _EVAL_11 & _EVAL_114;
  assign _EVAL_103 = _EVAL_46 & _EVAL_145;
  assign _EVAL_225 = _EVAL_24 & _EVAL_233;
  assign _EVAL_119 = ~_EVAL_120;
  assign _EVAL_300 = _EVAL_17 & _EVAL_244;
  assign _EVAL_139 = _EVAL_5 & _EVAL_203;
  assign _EVAL_248 = _EVAL_6 == 2'h0;
  assign _EVAL_274 = _EVAL_89 | _EVAL_147;
  assign _EVAL_102 = $signed(_EVAL_54) & -33'sh400000;
  assign _EVAL_244 = _EVAL_142 == 6'h0;
  assign _EVAL_21 = {1'b0,$signed(_EVAL_200)};
  assign _EVAL_17 = _EVAL_13 & _EVAL_11;
  assign _EVAL_33 = ~_EVAL_22;
  assign _EVAL_49 = _EVAL_19 | _EVAL_245;
  assign _EVAL_187 = _EVAL_103 | _EVAL_225;
  assign _EVAL_172 = _EVAL_175;
  assign _EVAL_106 = {{24'd0}, _EVAL_180};
  assign _EVAL_116 = _EVAL_74 & _EVAL_151;
  assign _EVAL_235 = _EVAL_103 | _EVAL_232;
  assign _EVAL_122 = _EVAL_297 | _EVAL_4;
  assign _EVAL_193 = ~_EVAL_224;
  assign _EVAL_83 = ~_EVAL_284;
  assign _EVAL_253 = _EVAL_158 | _EVAL_9;
  assign _EVAL_65 = _EVAL_5 & _EVAL_137;
  assign _EVAL_223 = _EVAL_2[0];
  assign _EVAL_286 = _EVAL_66 != _EVAL_250;
  assign _EVAL_214 = _EVAL_237 | _EVAL_4;
  assign _EVAL_302 = _EVAL_103 | _EVAL_202;
  assign _EVAL_39 = _EVAL_71 == 6'h0;
  assign _EVAL_190 = ~_EVAL_159;
  assign _EVAL_76 = _EVAL_0 == 3'h7;
  assign _EVAL_228 = $signed(_EVAL_44) & -33'sh5000;
  assign _EVAL_22 = _EVAL_235 | _EVAL_4;
  assign _EVAL_84 = ~_EVAL_167;
  assign _EVAL_191 = _EVAL_245 | _EVAL_118;
  assign _EVAL_163 = _EVAL_0[2];
  assign _EVAL_245 = $signed(_EVAL_172) == 33'sh0;
  assign _EVAL_99 = _EVAL_230 | _EVAL_4;
  assign _EVAL_212 = _EVAL_151 & _EVAL_79;
  assign _EVAL_53 = _EVAL_72[5:0];
  assign _EVAL_60 = _EVAL_153 == 32'h0;
  assign _EVAL_305 = _EVAL_96 | _EVAL_4;
  assign _EVAL_213 = _EVAL_168 & _EVAL_136;
  assign _EVAL_250 = _EVAL_16[0];
  assign _EVAL_82 = ~_EVAL_163;
  assign _EVAL_57 = ~_EVAL_206;
  assign _EVAL_243 = _EVAL_0 == 3'h3;
  assign _EVAL_128 = _EVAL_43 | _EVAL_4;
  assign _EVAL_79 = ~_EVAL_205;
  assign _EVAL_206 = _EVAL_264 | _EVAL_4;
  assign _EVAL_59 = ~_EVAL_268;
  assign _EVAL_63 = _EVAL_292 & _EVAL_256;
  assign _EVAL_141 = _EVAL_8 == 3'h4;
  assign _EVAL_68 = _EVAL_12 == _EVAL_51;
  assign _EVAL_168 = _EVAL_291[0];
  assign _EVAL_179 = _EVAL_2 == _EVAL_219;
  assign _EVAL_257 = _EVAL_3 >= 4'h2;
  assign _EVAL_211 = _EVAL_10 ^ 32'h3000;
  assign _EVAL_287 = _EVAL_11 & _EVAL_188;
  assign _EVAL_185 = _EVAL_2 <= 4'hb;
  assign _EVAL_178 = _EVAL_5 & _EVAL_216;
  assign _EVAL_285 = _EVAL_185 & _EVAL_235;
  assign _EVAL_151 = _EVAL_10[1];
  assign _EVAL_176 = ~_EVAL_250;
  assign _EVAL_121 = ~_EVAL_256;
  assign _EVAL_200 = _EVAL_10 ^ 32'h40000000;
  assign _EVAL_159 = _EVAL_253 | _EVAL_4;
  assign _EVAL_262 = ~_EVAL_38;
  assign _EVAL_240 = _EVAL_5 & _EVAL_76;
  assign _EVAL_92 = _EVAL_201 >> _EVAL_14;
  assign _EVAL_204 = ~_EVAL_166;
  assign _EVAL_146 = _EVAL_0 == 3'h5;
  assign _EVAL_138 = _EVAL_274 | _EVAL_157;
  assign _EVAL_263 = ~_EVAL_69;
  assign _EVAL_169 = _EVAL_100 | _EVAL_66;
  assign _EVAL_269 = _EVAL_185 | _EVAL_4;
  assign _EVAL_294 = _EVAL_102;
  assign _EVAL_259 = _EVAL_168 & _EVAL_212;
  assign _EVAL_295 = _EVAL_180[7:2];
  assign _EVAL_229 = ~_EVAL_99;
  assign _EVAL_232 = _EVAL_24 & _EVAL_266;
  assign _EVAL_237 = _EVAL_2 >= 4'h2;
  assign _EVAL_254 = _EVAL_237 | _EVAL_116;
  assign _EVAL_70 = _EVAL_0 == 3'h2;
  assign _EVAL_161 = ~_EVAL_80;
  assign _EVAL_108 = _EVAL_280 == 4'h0;
  assign _EVAL_162 = |_EVAL_100;
  assign _EVAL_42 = ~_EVAL_162;
  assign _EVAL_236 = 2'h1 << _EVAL_14;
  assign _EVAL_208 = ~_EVAL_7;
  assign _EVAL_77 = _EVAL_10 ^ 32'hc000000;
  assign _EVAL_109 = _EVAL_74 & _EVAL_131;
  assign _EVAL_69 = _EVAL_242 | _EVAL_4;
  assign _EVAL_105 = 2'h1 << _EVAL_223;
  assign _EVAL_186 = _EVAL_88;
  assign _EVAL_164 = _EVAL_142 - 6'h1;
  assign _EVAL_124 = _EVAL_8 == 3'h1;
  assign _EVAL_249 = ~_EVAL_31;
  assign _EVAL_98 = ~_EVAL_133;
  assign _EVAL_123 = _EVAL_8[0];
  assign _EVAL_227 = _EVAL_113 ? 2'h1 : 2'h0;
  assign _EVAL_31 = _EVAL_8 == 3'h6;
  assign _EVAL_160 = _EVAL_281[5:0];
  assign _EVAL_46 = _EVAL_2 <= 4'h8;
  assign _EVAL_27 = ~_EVAL_181;
  assign _EVAL_111 = ~_EVAL_94;
  assign _EVAL_231 = _EVAL_3 == _EVAL_173;
  assign _EVAL_54 = {1'b0,$signed(_EVAL_77)};
  assign _EVAL_90 = 23'hff << _EVAL_2;
  assign _EVAL_96 = ~_EVAL_100;
  assign _EVAL_239 = _EVAL_238;
  assign _EVAL_126 = ~_EVAL_214;
  assign _EVAL_18 = _EVAL_179 | _EVAL_4;
  assign _EVAL_210 = _EVAL_30[31:0];
  assign _EVAL_36 = _EVAL_10 ^ 32'h2000000;
  assign _EVAL_272 = _EVAL_187 | _EVAL_4;
  assign _EVAL_207 = _EVAL_42 | _EVAL_41;
  assign _EVAL_153 = _EVAL_10 & _EVAL_106;
  assign _EVAL_149 = _EVAL_7 == _EVAL_28;
  assign _EVAL_215 = _EVAL_110 < plusarg_reader_out;
  assign _EVAL_260 = _EVAL_10 == _EVAL_143;
  assign _EVAL_182 = _EVAL_5 & _EVAL_70;
  assign _EVAL_97 = ~_EVAL_14;
  assign _EVAL_140 = _EVAL_91 | _EVAL_4;
  assign _EVAL_195 = _EVAL_14 == _EVAL_270;
  assign _EVAL_155 = _EVAL_158 | _EVAL_4;
  assign _EVAL_217 = _EVAL_11 & _EVAL_124;
  assign _EVAL_242 = _EVAL_8 == _EVAL_125;
  assign _EVAL_266 = _EVAL_154 | _EVAL_198;
  assign _EVAL_34 = _EVAL_285 | _EVAL_4;
  assign _EVAL_66 = _EVAL_227[0];
  assign _EVAL_280 = _EVAL_7 & _EVAL_282;
  assign _EVAL_256 = _EVAL_104 == 6'h0;
  assign _EVAL_73 = _EVAL_149 | _EVAL_4;
  assign _EVAL_115 = $signed(_EVAL_294) == 33'sh0;
  assign _EVAL_44 = {1'b0,$signed(_EVAL_10)};
  assign _EVAL_171 = |_EVAL_66;
  assign _EVAL_64 = _EVAL_220 == 6'h0;
  assign _EVAL_147 = $signed(_EVAL_192) == 33'sh0;
  assign _EVAL_29 = ~_EVAL_34;
  assign _EVAL_275 = _EVAL_248 | _EVAL_4;
  assign _EVAL_72 = _EVAL_220 - 6'h1;
  assign _EVAL_188 = _EVAL_8 == 3'h0;
  assign _EVAL_268 = _EVAL_60 | _EVAL_4;
  assign _EVAL_145 = $signed(_EVAL_239) == 33'sh0;
  assign _EVAL_35 = {1'b0,$signed(_EVAL_289)};
  assign _EVAL_201 = _EVAL_66 | _EVAL_100;
  assign _EVAL_166 = _EVAL_196 | _EVAL_4;
  assign _EVAL_118 = $signed(_EVAL_186) == 33'sh0;
  assign _EVAL_19 = _EVAL_138 | _EVAL_115;
  assign _EVAL_89 = $signed(_EVAL_293) == 33'sh0;
  assign _EVAL_279 = ~_EVAL_64;
  assign _EVAL_273 = _EVAL_286 | _EVAL_67;
  assign _EVAL_209 = _EVAL_298;
  assign _EVAL_234 = ~_EVAL_50;
  assign _EVAL_271 = _EVAL_75[5:0];
  assign _EVAL_284 = _EVAL_231 | _EVAL_4;
  assign _EVAL_216 = _EVAL_0 == 3'h1;
  assign _EVAL_194 = _EVAL_5 & _EVAL_146;
  assign _EVAL_67 = ~_EVAL_171;
  assign _EVAL_85 = _EVAL_55[7:0];
  assign _EVAL_74 = _EVAL_291[1];
  assign _EVAL_197 = _EVAL_10 ^ 32'h20000000;
  assign _EVAL_226 = _EVAL_0 == 3'h0;
  assign _EVAL_276 = _EVAL_168 & _EVAL_165;
  assign _EVAL_158 = ~_EVAL_15;
  assign _EVAL_20 = _EVAL_5 & _EVAL_243;
  assign _EVAL_55 = 23'hff << _EVAL_3;
  assign _EVAL_282 = ~_EVAL_28;
  assign _EVAL_61 = _EVAL_152[7:2];
  assign _EVAL_16 = _EVAL_222 ? _EVAL_236 : 2'h0;
  assign _EVAL_148 = _EVAL_10 ^ 32'h80000000;
  assign _EVAL_218 = _EVAL_8 == 3'h2;
  assign _EVAL_165 = _EVAL_131 & _EVAL_79;
  assign _EVAL_167 = _EVAL_302 | _EVAL_4;
  assign _EVAL_81 = $signed(_EVAL_35) & -33'sh4000;
  assign _EVAL_297 = _EVAL_15 == _EVAL_255;
  assign _EVAL_130 = _EVAL_8 <= 3'h6;
  assign _EVAL_113 = _EVAL_292 & _EVAL_39;
  assign _EVAL_58 = ~_EVAL_128;
  assign _EVAL_292 = _EVAL & _EVAL_5;
  assign _EVAL_241 = _EVAL_207 | _EVAL_215;
  assign _EVAL_180 = ~_EVAL_144;
  assign _EVAL_88 = $signed(_EVAL_21) & -33'sh2000;
  assign _EVAL_91 = _EVAL_208 == 4'h0;
  assign _EVAL_224 = _EVAL_273 | _EVAL_4;
  assign _EVAL_24 = _EVAL_2 <= 4'h6;
  assign _EVAL_95 = _EVAL_241 | _EVAL_4;
  assign _EVAL_296 = ~_EVAL_269;
  assign _EVAL_93 = ~_EVAL_95;
  assign _EVAL_289 = _EVAL_10 ^ 32'h1800000;
  assign _EVAL_183 = {1'b0,$signed(_EVAL_211)};
  assign _EVAL_117 = _EVAL_11 & _EVAL_218;
  assign _EVAL_80 = _EVAL_257 | _EVAL_4;
  assign _EVAL_86 = _EVAL_195 | _EVAL_4;
  assign _EVAL_50 = _EVAL_108 | _EVAL_4;
  assign _EVAL_131 = ~_EVAL_151;
  assign _EVAL_288 = _EVAL_11 & _EVAL_279;
  assign _EVAL_75 = _EVAL_104 - 6'h1;
  assign _EVAL_299 = _EVAL_6 != 2'h2;
  assign _EVAL_41 = plusarg_reader_out == 32'h0;
  assign _EVAL_277 = ~_EVAL_275;
  assign _EVAL_233 = _EVAL_19 | _EVAL_198;
  assign _EVAL_278 = _EVAL_25 | _EVAL_184;
  assign _EVAL_26 = {1'b0,$signed(_EVAL_148)};
  assign _EVAL_112 = ~_EVAL_18;
  assign _EVAL_202 = _EVAL_24 & _EVAL_191;
  assign _EVAL_181 = _EVAL_130 | _EVAL_4;
  assign _EVAL_43 = _EVAL_6 <= 2'h2;
  assign _EVAL_114 = _EVAL_8 == 3'h5;
  assign _EVAL_238 = $signed(_EVAL_183) & -33'sh1000;
  assign _EVAL_170 = {1'b0,$signed(_EVAL_197)};
  assign _EVAL_127 = {1'b0,$signed(_EVAL_36)};
  assign _EVAL_137 = _EVAL_0 == 3'h4;
  assign _EVAL_144 = _EVAL_90[7:0];
  assign _EVAL_267 = ~_EVAL_129;
  assign _EVAL_184 = _EVAL_168 & _EVAL_47;
  assign _EVAL_189 = _EVAL_254 | _EVAL_259;
  assign _EVAL_56 = ~_EVAL_122;
  assign _EVAL_298 = $signed(_EVAL_26) & -33'sh4000;
  assign _EVAL_25 = _EVAL_237 | _EVAL_109;
  assign _EVAL_47 = _EVAL_131 & _EVAL_205;
  assign _EVAL_136 = _EVAL_151 & _EVAL_205;
  assign _EVAL_283 = _EVAL_17 & _EVAL_64;
  assign _EVAL_205 = _EVAL_10[0];
  assign _EVAL_293 = _EVAL_228;
  assign _EVAL_134 = _EVAL_164[5:0];
  assign _EVAL_157 = $signed(_EVAL_252) == 33'sh0;
  assign _EVAL_198 = $signed(_EVAL_209) == 33'sh0;
  assign _EVAL_196 = _EVAL_0 == _EVAL_132;
  assign _EVAL_129 = _EVAL_92 | _EVAL_4;
  assign _EVAL_37 = $signed(_EVAL_127) & -33'sh10000;
  assign _EVAL_156 = ~_EVAL_73;
  assign _EVAL_48 = _EVAL_292 | _EVAL_17;
  assign _EVAL_264 = _EVAL_6 == _EVAL_32;
  assign _EVAL_23 = _EVAL_254 | _EVAL_213;
  assign _EVAL_265 = _EVAL_11 & _EVAL_31;
  assign _EVAL_152 = ~_EVAL_85;
  assign _EVAL_133 = _EVAL_299 | _EVAL_4;
  assign _EVAL_38 = _EVAL_68 | _EVAL_4;
  assign _EVAL_251 = ~_EVAL_140;
  assign _EVAL_301 = _EVAL_25 | _EVAL_276;
  assign _EVAL_252 = _EVAL_37;
  always @(posedge _EVAL_1) begin
    if (_EVAL_283) begin
      _EVAL_32 <= _EVAL_6;
    end
    if (_EVAL_283) begin
      _EVAL_51 <= _EVAL_12;
    end
    if (_EVAL_4) begin
      _EVAL_71 <= 6'h0;
    end else if (_EVAL_292) begin
      if (_EVAL_39) begin
        if (_EVAL_82) begin
          _EVAL_71 <= _EVAL_295;
        end else begin
          _EVAL_71 <= 6'h0;
        end
      end else begin
        _EVAL_71 <= _EVAL_160;
      end
    end
    if (_EVAL_4) begin
      _EVAL_100 <= 1'h0;
    end else begin
      _EVAL_100 <= _EVAL_40;
    end
    if (_EVAL_4) begin
      _EVAL_104 <= 6'h0;
    end else if (_EVAL_292) begin
      if (_EVAL_256) begin
        if (_EVAL_82) begin
          _EVAL_104 <= _EVAL_295;
        end else begin
          _EVAL_104 <= 6'h0;
        end
      end else begin
        _EVAL_104 <= _EVAL_271;
      end
    end
    if (_EVAL_4) begin
      _EVAL_110 <= 32'h0;
    end else if (_EVAL_48) begin
      _EVAL_110 <= 32'h0;
    end else begin
      _EVAL_110 <= _EVAL_210;
    end
    if (_EVAL_283) begin
      _EVAL_125 <= _EVAL_8;
    end
    if (_EVAL_63) begin
      _EVAL_132 <= _EVAL_0;
    end
    if (_EVAL_4) begin
      _EVAL_142 <= 6'h0;
    end else if (_EVAL_17) begin
      if (_EVAL_244) begin
        if (_EVAL_123) begin
          _EVAL_142 <= _EVAL_61;
        end else begin
          _EVAL_142 <= 6'h0;
        end
      end else begin
        _EVAL_142 <= _EVAL_134;
      end
    end
    if (_EVAL_63) begin
      _EVAL_143 <= _EVAL_10;
    end
    if (_EVAL_283) begin
      _EVAL_173 <= _EVAL_3;
    end
    if (_EVAL_63) begin
      _EVAL_219 <= _EVAL_2;
    end
    if (_EVAL_4) begin
      _EVAL_220 <= 6'h0;
    end else if (_EVAL_17) begin
      if (_EVAL_64) begin
        if (_EVAL_123) begin
          _EVAL_220 <= _EVAL_61;
        end else begin
          _EVAL_220 <= 6'h0;
        end
      end else begin
        _EVAL_220 <= _EVAL_53;
      end
    end
    if (_EVAL_283) begin
      _EVAL_255 <= _EVAL_15;
    end
    if (_EVAL_283) begin
      _EVAL_270 <= _EVAL_14;
    end
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fb863f89)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_93) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_27) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7e8fc4b7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(45ff551c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_304) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d5cbdabf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_57) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_58) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7269f02f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc2beeb7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4786552)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(959cdfb8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_112) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc1b563c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5470e69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20e5d3c6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86ee7805)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e9b716c2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5561b88c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_83) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7b975e1b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_98) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3edf9fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_87) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5209d544)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_101) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(48a65634)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(65037290)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_11 & _EVAL_27) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_267) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cfb18c54)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_290) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cc01abd7)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(daa65bf4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9a213a79)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(28bf60e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bcb42a3d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_87) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(515c8c44)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b362f37)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bed45654)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9dad243b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6eeaace6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bd594864)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_234) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e0c8a470)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_263) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(62110a58)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5f763b70)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_98) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(468cdacc)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_251) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(15ef6059)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_262) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5ca9fc19)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_193) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(60452c0d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_33) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b657a8b0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_217 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_204) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2088c703)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_84) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b0fc9a2f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(3c59e8e6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_29) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_33) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a53e48bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(756755aa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_58) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_290) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_119) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e2c3572)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_182 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_93) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(24eba295)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1e10d3f8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_246 & _EVAL_29) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(fd082d6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(70ed1356)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b9e4e60d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(edf4ee28)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f42a5f4b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_83) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(aba38fd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_57) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f02a065f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1988960c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b405ca42)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_126) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(763446f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_156) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8b32ea5)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_113 & _EVAL_304) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e250f357)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_251) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(34ff87b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_126) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd2e1baa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_59) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b088ee76)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_112) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_52 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_101) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d1ff70c0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f3039c18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_156) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(21e33c08)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_193) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ed4ecac8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_258 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_117 & _EVAL_229) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a196fa6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_178 & _EVAL_234) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ac43fcff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9f89cf0c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_240 & _EVAL_78) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9dad243b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_84) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_139 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_277) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7c3d61eb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_265 & _EVAL_119) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_65 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_111) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a1d7925a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_288 & _EVAL_263) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_20 & _EVAL_59) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_194 & _EVAL_78) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_107 & _EVAL_204) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_287 & _EVAL_229) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_32 = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_51 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_71 = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_100 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_104 = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_110 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_125 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_132 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_142 = _RAND_8[5:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_143 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_173 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_219 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_220 = _RAND_12[5:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_255 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_270 = _RAND_14[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
