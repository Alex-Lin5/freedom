//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_138(
  input         _EVAL,
  input  [3:0]  _EVAL_0,
  input         _EVAL_1,
  output [2:0]  _EVAL_2,
  input  [3:0]  _EVAL_3,
  output        _EVAL_4,
  input  [1:0]  _EVAL_5,
  output        _EVAL_6,
  output [3:0]  _EVAL_7,
  input  [1:0]  _EVAL_8,
  output        _EVAL_9,
  input  [31:0] _EVAL_10,
  output        _EVAL_11,
  input  [3:0]  _EVAL_12,
  output        _EVAL_13,
  output        _EVAL_14,
  input  [2:0]  _EVAL_15,
  input  [2:0]  _EVAL_16,
  output        _EVAL_17,
  output        _EVAL_18,
  output [3:0]  _EVAL_19,
  input  [31:0] _EVAL_20,
  output        _EVAL_21,
  output [3:0]  _EVAL_22,
  input         _EVAL_23,
  output [1:0]  _EVAL_24,
  output [31:0] _EVAL_25,
  output        _EVAL_26,
  input         _EVAL_27,
  input  [3:0]  _EVAL_28,
  output [2:0]  _EVAL_29,
  input         _EVAL_30,
  input         _EVAL_31,
  input         _EVAL_32,
  input         _EVAL_33,
  output [3:0]  _EVAL_34,
  input  [3:0]  _EVAL_35,
  output        _EVAL_36,
  input  [31:0] _EVAL_37,
  output        _EVAL_38,
  output [31:0] _EVAL_39,
  input         _EVAL_40,
  input  [2:0]  _EVAL_41,
  input         _EVAL_42,
  output        _EVAL_43,
  output [2:0]  _EVAL_44,
  output [31:0] _EVAL_45,
  input         _EVAL_46,
  input         _EVAL_47,
  output [3:0]  _EVAL_48,
  output        _EVAL_49,
  output [1:0]  _EVAL_50,
  output [31:0] _EVAL_51,
  input         _EVAL_52,
  output [2:0]  _EVAL_53,
  input  [2:0]  _EVAL_54,
  input  [31:0] _EVAL_55,
  output [31:0] _EVAL_56,
  input  [1:0]  _EVAL_57,
  output        _EVAL_58,
  output [1:0]  _EVAL_59,
  output [3:0]  _EVAL_60,
  input         _EVAL_61,
  output [3:0]  _EVAL_62,
  input  [1:0]  _EVAL_63,
  input         _EVAL_64,
  output        _EVAL_65,
  input  [3:0]  _EVAL_66,
  output [3:0]  _EVAL_67,
  input         _EVAL_68,
  output        _EVAL_69,
  input         _EVAL_70,
  output [2:0]  _EVAL_71,
  input  [3:0]  _EVAL_72
);
  wire  bundleIn_0_d_sink__EVAL;
  wire [3:0] bundleIn_0_d_sink__EVAL_0;
  wire  bundleIn_0_d_sink__EVAL_1;
  wire  bundleIn_0_d_sink__EVAL_2;
  wire [31:0] bundleIn_0_d_sink__EVAL_3;
  wire  bundleIn_0_d_sink__EVAL_4;
  wire [1:0] bundleIn_0_d_sink__EVAL_5;
  wire  bundleIn_0_d_sink__EVAL_6;
  wire [31:0] bundleIn_0_d_sink__EVAL_7;
  wire [1:0] bundleIn_0_d_sink__EVAL_8;
  wire [1:0] bundleIn_0_d_sink__EVAL_9;
  wire  bundleIn_0_d_sink__EVAL_10;
  wire  bundleIn_0_d_sink__EVAL_11;
  wire  bundleIn_0_d_sink__EVAL_12;
  wire [1:0] bundleIn_0_d_sink__EVAL_13;
  wire [2:0] bundleIn_0_d_sink__EVAL_14;
  wire  bundleIn_0_d_sink__EVAL_15;
  wire  bundleIn_0_d_sink__EVAL_16;
  wire [1:0] bundleIn_0_d_sink__EVAL_17;
  wire  bundleIn_0_d_sink__EVAL_18;
  wire  bundleIn_0_d_sink__EVAL_19;
  wire [2:0] bundleIn_0_d_sink__EVAL_20;
  wire  bundleIn_0_d_sink__EVAL_21;
  wire [3:0] bundleIn_0_d_sink__EVAL_22;
  wire [3:0] bundleIn_0_d_sink__EVAL_23;
  wire [3:0] bundleIn_0_d_sink__EVAL_24;
  wire [3:0] bundleIn_0_d_sink__EVAL_25;
  wire  bundleIn_0_d_sink__EVAL_26;
  wire [2:0] bundleIn_0_d_sink__EVAL_27;
  wire [3:0] bundleIn_0_d_sink__EVAL_28;
  wire [31:0] bundleIn_0_d_sink__EVAL_29;
  wire  bundleIn_0_d_sink__EVAL_30;
  wire [31:0] bundleOut_0_a_source__EVAL;
  wire  bundleOut_0_a_source__EVAL_0;
  wire [2:0] bundleOut_0_a_source__EVAL_1;
  wire  bundleOut_0_a_source__EVAL_2;
  wire  bundleOut_0_a_source__EVAL_3;
  wire [2:0] bundleOut_0_a_source__EVAL_4;
  wire [2:0] bundleOut_0_a_source__EVAL_5;
  wire  bundleOut_0_a_source__EVAL_6;
  wire [31:0] bundleOut_0_a_source__EVAL_7;
  wire [31:0] bundleOut_0_a_source__EVAL_8;
  wire  bundleOut_0_a_source__EVAL_9;
  wire [3:0] bundleOut_0_a_source__EVAL_10;
  wire  bundleOut_0_a_source__EVAL_11;
  wire  bundleOut_0_a_source__EVAL_12;
  wire  bundleOut_0_a_source__EVAL_13;
  wire [3:0] bundleOut_0_a_source__EVAL_14;
  wire  bundleOut_0_a_source__EVAL_15;
  wire [1:0] bundleOut_0_a_source__EVAL_16;
  wire  bundleOut_0_a_source__EVAL_17;
  wire  bundleOut_0_a_source__EVAL_18;
  wire [3:0] bundleOut_0_a_source__EVAL_19;
  wire  bundleOut_0_a_source__EVAL_20;
  wire [3:0] bundleOut_0_a_source__EVAL_21;
  wire  bundleOut_0_a_source__EVAL_22;
  wire  bundleOut_0_a_source__EVAL_23;
  wire  bundleOut_0_a_source__EVAL_24;
  wire [2:0] bundleOut_0_a_source__EVAL_25;
  wire [31:0] bundleOut_0_a_source__EVAL_26;
  wire  bundleOut_0_a_source__EVAL_27;
  wire  bundleOut_0_a_source__EVAL_28;
  wire [31:0] bundleOut_0_a_source__EVAL_29;
  wire  bundleOut_0_a_source__EVAL_30;
  wire [3:0] bundleOut_0_a_source__EVAL_31;
  wire  bundleOut_0_a_source__EVAL_32;
  wire [31:0] bundleOut_0_a_source__EVAL_33;
  wire [3:0] bundleOut_0_a_source__EVAL_34;
  wire [3:0] bundleOut_0_a_source__EVAL_35;
  wire [2:0] bundleOut_0_a_source__EVAL_36;
  wire  bundleOut_0_a_source__EVAL_37;
  wire  bundleOut_0_a_source__EVAL_38;
  wire [2:0] bundleOut_0_a_source__EVAL_39;
  wire [3:0] bundleOut_0_a_source__EVAL_40;
  wire [3:0] bundleOut_0_a_source__EVAL_41;
  wire [1:0] bundleOut_0_a_source__EVAL_42;
  _EVAL_137 bundleIn_0_d_sink (
    ._EVAL(bundleIn_0_d_sink__EVAL),
    ._EVAL_0(bundleIn_0_d_sink__EVAL_0),
    ._EVAL_1(bundleIn_0_d_sink__EVAL_1),
    ._EVAL_2(bundleIn_0_d_sink__EVAL_2),
    ._EVAL_3(bundleIn_0_d_sink__EVAL_3),
    ._EVAL_4(bundleIn_0_d_sink__EVAL_4),
    ._EVAL_5(bundleIn_0_d_sink__EVAL_5),
    ._EVAL_6(bundleIn_0_d_sink__EVAL_6),
    ._EVAL_7(bundleIn_0_d_sink__EVAL_7),
    ._EVAL_8(bundleIn_0_d_sink__EVAL_8),
    ._EVAL_9(bundleIn_0_d_sink__EVAL_9),
    ._EVAL_10(bundleIn_0_d_sink__EVAL_10),
    ._EVAL_11(bundleIn_0_d_sink__EVAL_11),
    ._EVAL_12(bundleIn_0_d_sink__EVAL_12),
    ._EVAL_13(bundleIn_0_d_sink__EVAL_13),
    ._EVAL_14(bundleIn_0_d_sink__EVAL_14),
    ._EVAL_15(bundleIn_0_d_sink__EVAL_15),
    ._EVAL_16(bundleIn_0_d_sink__EVAL_16),
    ._EVAL_17(bundleIn_0_d_sink__EVAL_17),
    ._EVAL_18(bundleIn_0_d_sink__EVAL_18),
    ._EVAL_19(bundleIn_0_d_sink__EVAL_19),
    ._EVAL_20(bundleIn_0_d_sink__EVAL_20),
    ._EVAL_21(bundleIn_0_d_sink__EVAL_21),
    ._EVAL_22(bundleIn_0_d_sink__EVAL_22),
    ._EVAL_23(bundleIn_0_d_sink__EVAL_23),
    ._EVAL_24(bundleIn_0_d_sink__EVAL_24),
    ._EVAL_25(bundleIn_0_d_sink__EVAL_25),
    ._EVAL_26(bundleIn_0_d_sink__EVAL_26),
    ._EVAL_27(bundleIn_0_d_sink__EVAL_27),
    ._EVAL_28(bundleIn_0_d_sink__EVAL_28),
    ._EVAL_29(bundleIn_0_d_sink__EVAL_29),
    ._EVAL_30(bundleIn_0_d_sink__EVAL_30)
  );
  _EVAL_136 bundleOut_0_a_source (
    ._EVAL(bundleOut_0_a_source__EVAL),
    ._EVAL_0(bundleOut_0_a_source__EVAL_0),
    ._EVAL_1(bundleOut_0_a_source__EVAL_1),
    ._EVAL_2(bundleOut_0_a_source__EVAL_2),
    ._EVAL_3(bundleOut_0_a_source__EVAL_3),
    ._EVAL_4(bundleOut_0_a_source__EVAL_4),
    ._EVAL_5(bundleOut_0_a_source__EVAL_5),
    ._EVAL_6(bundleOut_0_a_source__EVAL_6),
    ._EVAL_7(bundleOut_0_a_source__EVAL_7),
    ._EVAL_8(bundleOut_0_a_source__EVAL_8),
    ._EVAL_9(bundleOut_0_a_source__EVAL_9),
    ._EVAL_10(bundleOut_0_a_source__EVAL_10),
    ._EVAL_11(bundleOut_0_a_source__EVAL_11),
    ._EVAL_12(bundleOut_0_a_source__EVAL_12),
    ._EVAL_13(bundleOut_0_a_source__EVAL_13),
    ._EVAL_14(bundleOut_0_a_source__EVAL_14),
    ._EVAL_15(bundleOut_0_a_source__EVAL_15),
    ._EVAL_16(bundleOut_0_a_source__EVAL_16),
    ._EVAL_17(bundleOut_0_a_source__EVAL_17),
    ._EVAL_18(bundleOut_0_a_source__EVAL_18),
    ._EVAL_19(bundleOut_0_a_source__EVAL_19),
    ._EVAL_20(bundleOut_0_a_source__EVAL_20),
    ._EVAL_21(bundleOut_0_a_source__EVAL_21),
    ._EVAL_22(bundleOut_0_a_source__EVAL_22),
    ._EVAL_23(bundleOut_0_a_source__EVAL_23),
    ._EVAL_24(bundleOut_0_a_source__EVAL_24),
    ._EVAL_25(bundleOut_0_a_source__EVAL_25),
    ._EVAL_26(bundleOut_0_a_source__EVAL_26),
    ._EVAL_27(bundleOut_0_a_source__EVAL_27),
    ._EVAL_28(bundleOut_0_a_source__EVAL_28),
    ._EVAL_29(bundleOut_0_a_source__EVAL_29),
    ._EVAL_30(bundleOut_0_a_source__EVAL_30),
    ._EVAL_31(bundleOut_0_a_source__EVAL_31),
    ._EVAL_32(bundleOut_0_a_source__EVAL_32),
    ._EVAL_33(bundleOut_0_a_source__EVAL_33),
    ._EVAL_34(bundleOut_0_a_source__EVAL_34),
    ._EVAL_35(bundleOut_0_a_source__EVAL_35),
    ._EVAL_36(bundleOut_0_a_source__EVAL_36),
    ._EVAL_37(bundleOut_0_a_source__EVAL_37),
    ._EVAL_38(bundleOut_0_a_source__EVAL_38),
    ._EVAL_39(bundleOut_0_a_source__EVAL_39),
    ._EVAL_40(bundleOut_0_a_source__EVAL_40),
    ._EVAL_41(bundleOut_0_a_source__EVAL_41),
    ._EVAL_42(bundleOut_0_a_source__EVAL_42)
  );
  assign bundleOut_0_a_source__EVAL_24 = _EVAL_61;
  assign bundleOut_0_a_source__EVAL_23 = _EVAL_30;
  assign _EVAL_53 = bundleOut_0_a_source__EVAL_25;
  assign bundleOut_0_a_source__EVAL_40 = _EVAL_0;
  assign bundleIn_0_d_sink__EVAL_20 = _EVAL_16;
  assign _EVAL_21 = bundleOut_0_a_source__EVAL_37;
  assign bundleIn_0_d_sink__EVAL_8 = _EVAL_63;
  assign _EVAL_25 = bundleOut_0_a_source__EVAL_8;
  assign bundleIn_0_d_sink__EVAL_18 = _EVAL_30;
  assign bundleIn_0_d_sink__EVAL_11 = _EVAL_64;
  assign _EVAL_18 = bundleIn_0_d_sink__EVAL_4;
  assign _EVAL_43 = bundleOut_0_a_source__EVAL_11;
  assign _EVAL_48 = bundleOut_0_a_source__EVAL_35;
  assign bundleOut_0_a_source__EVAL_9 = _EVAL_23;
  assign bundleOut_0_a_source__EVAL_15 = _EVAL_1;
  assign bundleOut_0_a_source__EVAL_31 = _EVAL_35;
  assign bundleIn_0_d_sink__EVAL_10 = _EVAL_46;
  assign bundleIn_0_d_sink__EVAL_6 = _EVAL_33;
  assign _EVAL_17 = bundleIn_0_d_sink__EVAL_21;
  assign bundleOut_0_a_source__EVAL_16 = _EVAL_8;
  assign _EVAL_34 = bundleOut_0_a_source__EVAL_10;
  assign bundleOut_0_a_source__EVAL_28 = _EVAL_47;
  assign bundleIn_0_d_sink__EVAL_19 = _EVAL_31;
  assign bundleIn_0_d_sink__EVAL_0 = _EVAL_72;
  assign bundleIn_0_d_sink__EVAL_2 = _EVAL_27;
  assign bundleIn_0_d_sink__EVAL_26 = _EVAL_70;
  assign _EVAL_6 = bundleOut_0_a_source__EVAL_0;
  assign bundleIn_0_d_sink__EVAL_15 = _EVAL_42;
  assign bundleIn_0_d_sink__EVAL_22 = _EVAL_66;
  assign _EVAL_67 = bundleOut_0_a_source__EVAL_19;
  assign bundleOut_0_a_source__EVAL_7 = _EVAL_55;
  assign _EVAL_44 = bundleOut_0_a_source__EVAL_39;
  assign bundleIn_0_d_sink__EVAL = _EVAL_40;
  assign bundleIn_0_d_sink__EVAL_12 = _EVAL_68;
  assign bundleIn_0_d_sink__EVAL_25 = _EVAL_3;
  assign _EVAL_14 = bundleOut_0_a_source__EVAL_18;
  assign _EVAL_38 = bundleOut_0_a_source__EVAL_13;
  assign bundleOut_0_a_source__EVAL_27 = _EVAL_32;
  assign _EVAL_51 = bundleOut_0_a_source__EVAL;
  assign _EVAL_9 = bundleIn_0_d_sink__EVAL_1;
  assign bundleIn_0_d_sink__EVAL_17 = _EVAL_5;
  assign _EVAL_50 = bundleIn_0_d_sink__EVAL_13;
  assign bundleOut_0_a_source__EVAL_14 = _EVAL_12;
  assign _EVAL_69 = bundleOut_0_a_source__EVAL_30;
  assign _EVAL_26 = bundleOut_0_a_source__EVAL_22;
  assign _EVAL_49 = bundleOut_0_a_source__EVAL_6;
  assign bundleIn_0_d_sink__EVAL_5 = _EVAL_57;
  assign _EVAL_7 = bundleIn_0_d_sink__EVAL_24;
  assign bundleOut_0_a_source__EVAL_2 = _EVAL_52;
  assign _EVAL_65 = bundleOut_0_a_source__EVAL_32;
  assign _EVAL_59 = bundleOut_0_a_source__EVAL_42;
  assign _EVAL_2 = bundleOut_0_a_source__EVAL_36;
  assign _EVAL_11 = bundleOut_0_a_source__EVAL_12;
  assign _EVAL_13 = bundleOut_0_a_source__EVAL_3;
  assign _EVAL_60 = bundleOut_0_a_source__EVAL_34;
  assign _EVAL_45 = bundleIn_0_d_sink__EVAL_7;
  assign bundleIn_0_d_sink__EVAL_23 = _EVAL_28;
  assign _EVAL_39 = bundleOut_0_a_source__EVAL_33;
  assign bundleIn_0_d_sink__EVAL_29 = _EVAL_20;
  assign _EVAL_71 = bundleIn_0_d_sink__EVAL_14;
  assign _EVAL_19 = bundleOut_0_a_source__EVAL_41;
  assign _EVAL_22 = bundleIn_0_d_sink__EVAL_28;
  assign bundleIn_0_d_sink__EVAL_3 = _EVAL_37;
  assign _EVAL_62 = bundleOut_0_a_source__EVAL_21;
  assign bundleOut_0_a_source__EVAL_29 = _EVAL_10;
  assign bundleIn_0_d_sink__EVAL_27 = _EVAL_15;
  assign bundleOut_0_a_source__EVAL_38 = _EVAL;
  assign _EVAL_36 = bundleOut_0_a_source__EVAL_20;
  assign bundleOut_0_a_source__EVAL_17 = _EVAL_31;
  assign _EVAL_56 = bundleOut_0_a_source__EVAL_26;
  assign _EVAL_29 = bundleOut_0_a_source__EVAL_5;
  assign _EVAL_24 = bundleIn_0_d_sink__EVAL_9;
  assign bundleOut_0_a_source__EVAL_1 = _EVAL_54;
  assign _EVAL_58 = bundleIn_0_d_sink__EVAL_16;
  assign bundleOut_0_a_source__EVAL_4 = _EVAL_41;
  assign _EVAL_4 = bundleIn_0_d_sink__EVAL_30;
endmodule
