//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_14(
  input  [2:0]  _EVAL,
  output        _EVAL_0,
  input  [2:0]  _EVAL_1,
  output        _EVAL_2,
  input         _EVAL_3,
  input  [31:0] _EVAL_4,
  output [4:0]  _EVAL_5,
  output [31:0] _EVAL_6,
  input         _EVAL_7,
  input  [4:0]  _EVAL_8,
  output        _EVAL_9,
  output        _EVAL_10,
  input         _EVAL_11,
  output [2:0]  _EVAL_12,
  output        _EVAL_13,
  output [1:0]  _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  output [2:0]  _EVAL_17,
  input         _EVAL_18
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_19;
  reg [31:0] _EVAL_20 [0:2];
  wire [31:0] _EVAL_20__EVAL_21_data;
  wire [1:0] _EVAL_20__EVAL_21_addr;
  wire [31:0] _EVAL_20__EVAL_22_data;
  wire [1:0] _EVAL_20__EVAL_22_addr;
  wire  _EVAL_20__EVAL_22_mask;
  wire  _EVAL_20__EVAL_22_en;
  wire [2:0] _EVAL_24;
  wire  _EVAL_26;
  reg  _EVAL_27 [0:2];
  wire  _EVAL_27__EVAL_28_data;
  wire [1:0] _EVAL_27__EVAL_28_addr;
  wire  _EVAL_27__EVAL_29_data;
  wire [1:0] _EVAL_27__EVAL_29_addr;
  wire  _EVAL_27__EVAL_29_mask;
  wire  _EVAL_27__EVAL_29_en;
  reg  _EVAL_31 [0:2];
  wire  _EVAL_31__EVAL_32_data;
  wire [1:0] _EVAL_31__EVAL_32_addr;
  wire  _EVAL_31__EVAL_33_data;
  wire [1:0] _EVAL_31__EVAL_33_addr;
  wire  _EVAL_31__EVAL_33_mask;
  wire  _EVAL_31__EVAL_33_en;
  wire [1:0] _EVAL_34;
  reg  _EVAL_35;
  reg [1:0] _EVAL_36;
  reg [1:0] _EVAL_37;
  wire [1:0] _EVAL_38;
  wire  _EVAL_39;
  wire  _EVAL_40;
  reg [2:0] _EVAL_41 [0:2];
  wire [2:0] _EVAL_41__EVAL_42_data;
  wire [1:0] _EVAL_41__EVAL_42_addr;
  wire [2:0] _EVAL_41__EVAL_43_data;
  wire [1:0] _EVAL_41__EVAL_43_addr;
  wire  _EVAL_41__EVAL_43_mask;
  wire  _EVAL_41__EVAL_43_en;
  wire  _EVAL_44;
  reg [4:0] _EVAL_45 [0:2];
  wire [4:0] _EVAL_45__EVAL_46_data;
  wire [1:0] _EVAL_45__EVAL_46_addr;
  wire [4:0] _EVAL_45__EVAL_47_data;
  wire [1:0] _EVAL_45__EVAL_47_addr;
  wire  _EVAL_45__EVAL_47_mask;
  wire  _EVAL_45__EVAL_47_en;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire  _EVAL_51;
  reg [1:0] _EVAL_53 [0:2];
  wire [1:0] _EVAL_53__EVAL_54_data;
  wire [1:0] _EVAL_53__EVAL_54_addr;
  wire [1:0] _EVAL_53__EVAL_55_data;
  wire [1:0] _EVAL_53__EVAL_55_addr;
  wire  _EVAL_53__EVAL_55_mask;
  wire  _EVAL_53__EVAL_55_en;
  wire  _EVAL_56;
  wire [2:0] _EVAL_57;
  wire  _EVAL_58;
  reg  _EVAL_59 [0:2];
  wire  _EVAL_59__EVAL_60_data;
  wire [1:0] _EVAL_59__EVAL_60_addr;
  wire  _EVAL_59__EVAL_61_data;
  wire [1:0] _EVAL_59__EVAL_61_addr;
  wire  _EVAL_59__EVAL_61_mask;
  wire  _EVAL_59__EVAL_61_en;
  wire  _EVAL_63;
  wire  _EVAL_64;
  reg [2:0] _EVAL_65 [0:2];
  wire [2:0] _EVAL_65__EVAL_66_data;
  wire [1:0] _EVAL_65__EVAL_66_addr;
  wire [2:0] _EVAL_65__EVAL_67_data;
  wire [1:0] _EVAL_65__EVAL_67_addr;
  wire  _EVAL_65__EVAL_67_mask;
  wire  _EVAL_65__EVAL_67_en;
  assign _EVAL_20__EVAL_21_addr = _EVAL_37;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _EVAL_20__EVAL_21_data = _EVAL_20[_EVAL_20__EVAL_21_addr];
  `else
  assign _EVAL_20__EVAL_21_data = _EVAL_20__EVAL_21_addr >= 2'h3 ? _RAND_1[31:0] : _EVAL_20[_EVAL_20__EVAL_21_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _EVAL_20__EVAL_22_data = _EVAL_4;
  assign _EVAL_20__EVAL_22_addr = _EVAL_36;
  assign _EVAL_20__EVAL_22_mask = 1'h1;
  assign _EVAL_20__EVAL_22_en = _EVAL_58 ? _EVAL_64 : _EVAL_19;
  assign _EVAL_27__EVAL_28_addr = _EVAL_37;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _EVAL_27__EVAL_28_data = _EVAL_27[_EVAL_27__EVAL_28_addr];
  `else
  assign _EVAL_27__EVAL_28_data = _EVAL_27__EVAL_28_addr >= 2'h3 ? _RAND_3[0:0] : _EVAL_27[_EVAL_27__EVAL_28_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _EVAL_27__EVAL_29_data = _EVAL_7;
  assign _EVAL_27__EVAL_29_addr = _EVAL_36;
  assign _EVAL_27__EVAL_29_mask = 1'h1;
  assign _EVAL_27__EVAL_29_en = _EVAL_58 ? _EVAL_64 : _EVAL_19;
  assign _EVAL_31__EVAL_32_addr = _EVAL_37;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _EVAL_31__EVAL_32_data = _EVAL_31[_EVAL_31__EVAL_32_addr];
  `else
  assign _EVAL_31__EVAL_32_data = _EVAL_31__EVAL_32_addr >= 2'h3 ? _RAND_5[0:0] : _EVAL_31[_EVAL_31__EVAL_32_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _EVAL_31__EVAL_33_data = _EVAL_3;
  assign _EVAL_31__EVAL_33_addr = _EVAL_36;
  assign _EVAL_31__EVAL_33_mask = 1'h1;
  assign _EVAL_31__EVAL_33_en = _EVAL_58 ? _EVAL_64 : _EVAL_19;
  assign _EVAL_41__EVAL_42_addr = _EVAL_37;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _EVAL_41__EVAL_42_data = _EVAL_41[_EVAL_41__EVAL_42_addr];
  `else
  assign _EVAL_41__EVAL_42_data = _EVAL_41__EVAL_42_addr >= 2'h3 ? _RAND_10[2:0] : _EVAL_41[_EVAL_41__EVAL_42_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _EVAL_41__EVAL_43_data = _EVAL;
  assign _EVAL_41__EVAL_43_addr = _EVAL_36;
  assign _EVAL_41__EVAL_43_mask = 1'h1;
  assign _EVAL_41__EVAL_43_en = _EVAL_58 ? _EVAL_64 : _EVAL_19;
  assign _EVAL_45__EVAL_46_addr = _EVAL_37;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _EVAL_45__EVAL_46_data = _EVAL_45[_EVAL_45__EVAL_46_addr];
  `else
  assign _EVAL_45__EVAL_46_data = _EVAL_45__EVAL_46_addr >= 2'h3 ? _RAND_12[4:0] : _EVAL_45[_EVAL_45__EVAL_46_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _EVAL_45__EVAL_47_data = _EVAL_8;
  assign _EVAL_45__EVAL_47_addr = _EVAL_36;
  assign _EVAL_45__EVAL_47_mask = 1'h1;
  assign _EVAL_45__EVAL_47_en = _EVAL_58 ? _EVAL_64 : _EVAL_19;
  assign _EVAL_53__EVAL_54_addr = _EVAL_37;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _EVAL_53__EVAL_54_data = _EVAL_53[_EVAL_53__EVAL_54_addr];
  `else
  assign _EVAL_53__EVAL_54_data = _EVAL_53__EVAL_54_addr >= 2'h3 ? _RAND_14[1:0] : _EVAL_53[_EVAL_53__EVAL_54_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _EVAL_53__EVAL_55_data = 2'h0;
  assign _EVAL_53__EVAL_55_addr = _EVAL_36;
  assign _EVAL_53__EVAL_55_mask = 1'h1;
  assign _EVAL_53__EVAL_55_en = _EVAL_58 ? _EVAL_64 : _EVAL_19;
  assign _EVAL_59__EVAL_60_addr = _EVAL_37;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _EVAL_59__EVAL_60_data = _EVAL_59[_EVAL_59__EVAL_60_addr];
  `else
  assign _EVAL_59__EVAL_60_data = _EVAL_59__EVAL_60_addr >= 2'h3 ? _RAND_16[0:0] : _EVAL_59[_EVAL_59__EVAL_60_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _EVAL_59__EVAL_61_data = 1'h0;
  assign _EVAL_59__EVAL_61_addr = _EVAL_36;
  assign _EVAL_59__EVAL_61_mask = 1'h1;
  assign _EVAL_59__EVAL_61_en = _EVAL_58 ? _EVAL_64 : _EVAL_19;
  assign _EVAL_65__EVAL_66_addr = _EVAL_37;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _EVAL_65__EVAL_66_data = _EVAL_65[_EVAL_65__EVAL_66_addr];
  `else
  assign _EVAL_65__EVAL_66_data = _EVAL_65__EVAL_66_addr >= 2'h3 ? _RAND_18[2:0] : _EVAL_65[_EVAL_65__EVAL_66_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _EVAL_65__EVAL_67_data = _EVAL_1;
  assign _EVAL_65__EVAL_67_addr = _EVAL_36;
  assign _EVAL_65__EVAL_67_mask = 1'h1;
  assign _EVAL_65__EVAL_67_en = _EVAL_58 ? _EVAL_64 : _EVAL_19;
  assign _EVAL_12 = _EVAL_58 ? _EVAL_1 : _EVAL_65__EVAL_66_data;
  assign _EVAL_64 = _EVAL_11 ? 1'h0 : _EVAL_19;
  assign _EVAL_63 = _EVAL_58 ? _EVAL_64 : _EVAL_19;
  assign _EVAL_48 = _EVAL_11 & _EVAL_10;
  assign _EVAL_24 = _EVAL_37 + 2'h1;
  assign _EVAL_50 = _EVAL_36 == _EVAL_37;
  assign _EVAL_9 = _EVAL_58 ? _EVAL_7 : _EVAL_27__EVAL_28_data;
  assign _EVAL_6 = _EVAL_58 ? _EVAL_4 : _EVAL_20__EVAL_21_data;
  assign _EVAL_58 = _EVAL_50 & _EVAL_44;
  assign _EVAL_56 = _EVAL_50 & _EVAL_35;
  assign _EVAL_19 = _EVAL_13 & _EVAL_15;
  assign _EVAL_26 = _EVAL_36 == 2'h2;
  assign _EVAL_10 = _EVAL_15 | _EVAL_51;
  assign _EVAL_57 = _EVAL_36 + 2'h1;
  assign _EVAL_17 = _EVAL_58 ? _EVAL : _EVAL_41__EVAL_42_data;
  assign _EVAL_39 = _EVAL_63 != _EVAL_40;
  assign _EVAL_34 = _EVAL_24[1:0];
  assign _EVAL_5 = _EVAL_58 ? _EVAL_8 : _EVAL_45__EVAL_46_data;
  assign _EVAL_51 = ~_EVAL_58;
  assign _EVAL_13 = ~_EVAL_56;
  assign _EVAL_14 = _EVAL_58 ? 2'h0 : _EVAL_53__EVAL_54_data;
  assign _EVAL_40 = _EVAL_58 ? 1'h0 : _EVAL_48;
  assign _EVAL_0 = _EVAL_58 ? _EVAL_3 : _EVAL_31__EVAL_32_data;
  assign _EVAL_49 = _EVAL_37 == 2'h2;
  assign _EVAL_2 = _EVAL_58 ? 1'h0 : _EVAL_59__EVAL_60_data;
  assign _EVAL_44 = ~_EVAL_35;
  assign _EVAL_38 = _EVAL_57[1:0];
  always @(posedge _EVAL_16) begin
    if(_EVAL_20__EVAL_22_en & _EVAL_20__EVAL_22_mask) begin
      _EVAL_20[_EVAL_20__EVAL_22_addr] <= _EVAL_20__EVAL_22_data;
    end
    if(_EVAL_27__EVAL_29_en & _EVAL_27__EVAL_29_mask) begin
      _EVAL_27[_EVAL_27__EVAL_29_addr] <= _EVAL_27__EVAL_29_data;
    end
    if(_EVAL_31__EVAL_33_en & _EVAL_31__EVAL_33_mask) begin
      _EVAL_31[_EVAL_31__EVAL_33_addr] <= _EVAL_31__EVAL_33_data;
    end
    if (_EVAL_18) begin
      _EVAL_35 <= 1'h0;
    end else if (_EVAL_39) begin
      if (_EVAL_58) begin
        if (_EVAL_11) begin
          _EVAL_35 <= 1'h0;
        end else begin
          _EVAL_35 <= _EVAL_19;
        end
      end else begin
        _EVAL_35 <= _EVAL_19;
      end
    end
    if (_EVAL_18) begin
      _EVAL_36 <= 2'h0;
    end else if (_EVAL_63) begin
      if (_EVAL_26) begin
        _EVAL_36 <= 2'h0;
      end else begin
        _EVAL_36 <= _EVAL_38;
      end
    end
    if (_EVAL_18) begin
      _EVAL_37 <= 2'h0;
    end else if (_EVAL_40) begin
      if (_EVAL_49) begin
        _EVAL_37 <= 2'h0;
      end else begin
        _EVAL_37 <= _EVAL_34;
      end
    end
    if(_EVAL_41__EVAL_43_en & _EVAL_41__EVAL_43_mask) begin
      _EVAL_41[_EVAL_41__EVAL_43_addr] <= _EVAL_41__EVAL_43_data;
    end
    if(_EVAL_45__EVAL_47_en & _EVAL_45__EVAL_47_mask) begin
      _EVAL_45[_EVAL_45__EVAL_47_addr] <= _EVAL_45__EVAL_47_data;
    end
    if(_EVAL_53__EVAL_55_en & _EVAL_53__EVAL_55_mask) begin
      _EVAL_53[_EVAL_53__EVAL_55_addr] <= _EVAL_53__EVAL_55_data;
    end
    if(_EVAL_59__EVAL_61_en & _EVAL_59__EVAL_61_mask) begin
      _EVAL_59[_EVAL_59__EVAL_61_addr] <= _EVAL_59__EVAL_61_data;
    end
    if(_EVAL_65__EVAL_67_en & _EVAL_65__EVAL_67_mask) begin
      _EVAL_65[_EVAL_65__EVAL_67_addr] <= _EVAL_65__EVAL_67_data;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_5 = {1{`RANDOM}};
  _RAND_10 = {1{`RANDOM}};
  _RAND_12 = {1{`RANDOM}};
  _RAND_14 = {1{`RANDOM}};
  _RAND_16 = {1{`RANDOM}};
  _RAND_18 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _EVAL_20[initvar] = _RAND_0[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _EVAL_27[initvar] = _RAND_2[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _EVAL_31[initvar] = _RAND_4[0:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _EVAL_41[initvar] = _RAND_9[2:0];
  _RAND_11 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _EVAL_45[initvar] = _RAND_11[4:0];
  _RAND_13 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _EVAL_53[initvar] = _RAND_13[1:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _EVAL_59[initvar] = _RAND_15[0:0];
  _RAND_17 = {1{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _EVAL_65[initvar] = _RAND_17[2:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _EVAL_35 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_36 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_37 = _RAND_8[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
