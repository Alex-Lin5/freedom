//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_92_assert(
  input  [2:0]  _EVAL_0,
  input         _EVAL_2,
  input  [9:0]  _EVAL_6,
  input  [2:0]  _EVAL_9,
  input         _EVAL_11,
  input  [4:0]  _EVAL_12,
  input  [3:0]  _EVAL_14,
  input  [2:0]  _EVAL_15,
  input         _EVAL_16,
  input  [14:0] _EVAL_21,
  input         _EVAL_26,
  input         _EVAL_27,
  input  [2:0]  _EVAL_28,
  input         _EVAL_30,
  input         _EVAL_41,
  input  [2:0]  _EVAL_45,
  input         _EVAL_89,
  input         _EVAL_98,
  input  [2:0]  _EVAL_115,
  input         repeater__EVAL_10,
  input         repeater__EVAL_15,
  input  [3:0]  repeater__EVAL_20
);
  wire  _EVAL_40;
  wire  _EVAL_55;
  wire  _EVAL_58;
  wire [2:0] monitor__EVAL;
  wire [2:0] monitor__EVAL_0;
  wire  monitor__EVAL_1;
  wire [4:0] monitor__EVAL_2;
  wire  monitor__EVAL_3;
  wire  monitor__EVAL_4;
  wire [2:0] monitor__EVAL_5;
  wire  monitor__EVAL_6;
  wire  monitor__EVAL_7;
  wire  monitor__EVAL_8;
  wire [3:0] monitor__EVAL_9;
  wire [4:0] monitor__EVAL_10;
  wire [2:0] monitor__EVAL_11;
  wire  monitor__EVAL_12;
  wire [14:0] monitor__EVAL_13;
  wire [2:0] monitor__EVAL_14;
  wire  _EVAL_70;
  wire  _EVAL_80;
  wire  _EVAL_100;
  wire  _EVAL_114;
  wire  _EVAL_123;
  _EVAL_90_assert monitor (
    ._EVAL(monitor__EVAL),
    ._EVAL_0(monitor__EVAL_0),
    ._EVAL_1(monitor__EVAL_1),
    ._EVAL_2(monitor__EVAL_2),
    ._EVAL_3(monitor__EVAL_3),
    ._EVAL_4(monitor__EVAL_4),
    ._EVAL_5(monitor__EVAL_5),
    ._EVAL_6(monitor__EVAL_6),
    ._EVAL_7(monitor__EVAL_7),
    ._EVAL_8(monitor__EVAL_8),
    ._EVAL_9(monitor__EVAL_9),
    ._EVAL_10(monitor__EVAL_10),
    ._EVAL_11(monitor__EVAL_11),
    ._EVAL_12(monitor__EVAL_12),
    ._EVAL_13(monitor__EVAL_13),
    ._EVAL_14(monitor__EVAL_14)
  );
  assign monitor__EVAL_13 = _EVAL_21;
  assign _EVAL_70 = _EVAL_100 | _EVAL_58;
  assign _EVAL_40 = _EVAL_100 | _EVAL_98;
  assign _EVAL_55 = ~_EVAL_80;
  assign monitor__EVAL_12 = repeater__EVAL_10;
  assign monitor__EVAL_7 = _EVAL_30;
  assign _EVAL_123 = ~_EVAL_114;
  assign monitor__EVAL_11 = _EVAL_9;
  assign monitor__EVAL_6 = _EVAL_2;
  assign monitor__EVAL_9 = _EVAL_14;
  assign monitor__EVAL_14 = _EVAL_28;
  assign monitor__EVAL_3 = _EVAL_26 & _EVAL_89;
  assign _EVAL_100 = ~repeater__EVAL_15;
  assign monitor__EVAL_2 = _EVAL_12;
  assign monitor__EVAL_5 = _EVAL_15;
  assign monitor__EVAL_8 = _EVAL_27;
  assign monitor__EVAL_0 = _EVAL_41 ? _EVAL_45 : _EVAL_115;
  assign monitor__EVAL_10 = _EVAL_6[9:5];
  assign monitor__EVAL_1 = _EVAL_16;
  assign monitor__EVAL = _EVAL_0;
  assign _EVAL_58 = repeater__EVAL_20 == 4'hf;
  assign _EVAL_114 = _EVAL_40 | _EVAL_27;
  assign monitor__EVAL_4 = _EVAL_11;
  assign _EVAL_80 = _EVAL_70 | _EVAL_27;
  always @(posedge _EVAL_16) begin
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_123) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b22d1eaf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7986d96b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_123) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end

endmodule
