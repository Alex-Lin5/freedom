//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_128(
  input  [31:0] _EVAL,
  input         _EVAL_0,
  input         _EVAL_1,
  output        _EVAL_2,
  output        _EVAL_3,
  input         _EVAL_4,
  input         _EVAL_5,
  output        _EVAL_6,
  input  [1:0]  _EVAL_7,
  input  [31:0] _EVAL_8,
  output        _EVAL_9,
  input         _EVAL_10,
  input         _EVAL_11,
  input         _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input         _EVAL_17,
  input  [1:0]  _EVAL_18,
  input  [1:0]  _EVAL_19,
  input         _EVAL_20,
  input  [31:0] _EVAL_21,
  input         _EVAL_22,
  input  [31:0] _EVAL_23,
  input         _EVAL_24,
  output        _EVAL_25,
  input         _EVAL_26,
  input         _EVAL_27,
  output        _EVAL_28,
  input  [31:0] _EVAL_29,
  input         _EVAL_30,
  input  [31:0] _EVAL_31,
  input         _EVAL_32,
  input         _EVAL_33,
  input  [1:0]  _EVAL_34,
  input         _EVAL_35,
  input         _EVAL_36,
  input         _EVAL_37,
  input         _EVAL_38,
  input         _EVAL_39,
  input         _EVAL_40,
  input         _EVAL_41,
  input  [1:0]  _EVAL_42,
  input         _EVAL_43
);
  wire  _EVAL_44;
  wire  _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire  _EVAL_49;
  wire  _EVAL_50;
  wire [31:0] _EVAL_51;
  wire  _EVAL_52;
  wire  _EVAL_53;
  wire  _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_60;
  wire  _EVAL_61;
  wire  _EVAL_62;
  wire [3:0] _EVAL_63;
  wire  _EVAL_64;
  wire [3:0] _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire [31:0] _EVAL_69;
  wire  _EVAL_70;
  wire [31:0] _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire  _EVAL_77;
  wire  _EVAL_78;
  wire [3:0] _EVAL_79;
  wire  _EVAL_80;
  wire  _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire  _EVAL_84;
  wire [31:0] _EVAL_85;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire [31:0] _EVAL_88;
  wire  _EVAL_89;
  wire [31:0] _EVAL_90;
  wire  _EVAL_91;
  wire  _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_97;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire [31:0] _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire  _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_109;
  wire  _EVAL_110;
  wire  _EVAL_111;
  wire  _EVAL_112;
  wire [31:0] _EVAL_113;
  wire  _EVAL_114;
  wire  _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire [3:0] _EVAL_118;
  wire  _EVAL_119;
  wire  _EVAL_120;
  wire  _EVAL_121;
  wire  _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire [31:0] _EVAL_126;
  wire  _EVAL_127;
  wire [3:0] _EVAL_128;
  wire  _EVAL_129;
  wire  _EVAL_130;
  wire  _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire [3:0] _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_136;
  wire  _EVAL_137;
  wire [31:0] _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_141;
  wire  _EVAL_142;
  wire  _EVAL_143;
  wire [31:0] _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire  _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire  _EVAL_155;
  wire  _EVAL_156;
  wire [3:0] _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire  _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire [31:0] _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire  _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire [31:0] _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire  _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire [3:0] _EVAL_180;
  wire  _EVAL_181;
  wire  _EVAL_182;
  wire [3:0] _EVAL_183;
  wire [31:0] _EVAL_184;
  wire  _EVAL_185;
  wire [3:0] _EVAL_186;
  wire [31:0] _EVAL_187;
  wire  _EVAL_188;
  wire  _EVAL_189;
  wire  _EVAL_190;
  wire [31:0] _EVAL_191;
  wire [31:0] _EVAL_192;
  wire  _EVAL_193;
  wire [31:0] _EVAL_194;
  wire [31:0] _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire  _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire [3:0] _EVAL_203;
  wire  _EVAL_204;
  wire  _EVAL_205;
  wire  _EVAL_206;
  wire [31:0] _EVAL_207;
  wire  _EVAL_208;
  wire  _EVAL_209;
  wire  _EVAL_210;
  wire  _EVAL_211;
  wire [31:0] _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire  _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire [3:0] _EVAL_221;
  wire  _EVAL_222;
  wire [31:0] _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  assign _EVAL_113 = _EVAL_126 | _EVAL_69;
  assign _EVAL_209 = _EVAL_64 & _EVAL_37;
  assign _EVAL_98 = _EVAL_82 & _EVAL_77;
  assign _EVAL_169 = _EVAL_156 ? _EVAL_114 : _EVAL_222;
  assign _EVAL_179 = _EVAL_34[0];
  assign _EVAL_90 = _EVAL_207 | _EVAL_138;
  assign _EVAL_198 = _EVAL_140 & _EVAL_33;
  assign _EVAL_163 = _EVAL_188 & _EVAL_80;
  assign _EVAL_158 = _EVAL_21[0];
  assign _EVAL_115 = _EVAL_29 >= _EVAL_8;
  assign _EVAL_54 = _EVAL_170 ? _EVAL_149 : _EVAL_200;
  assign _EVAL_72 = _EVAL_127 & _EVAL_67;
  assign _EVAL_3 = _EVAL_116 ? _EVAL_45 : _EVAL_181;
  assign _EVAL_196 = _EVAL_217 & _EVAL_225;
  assign _EVAL_118 = {_EVAL_14,1'h0,1'h0,_EVAL_15};
  assign _EVAL_141 = _EVAL_199 & _EVAL_169;
  assign _EVAL_116 = _EVAL_91 & _EVAL_84;
  assign _EVAL_105 = _EVAL_68 & _EVAL_78;
  assign _EVAL_123 = _EVAL_204 & _EVAL_141;
  assign _EVAL_107 = _EVAL_204 | _EVAL_145;
  assign _EVAL_138 = {{28'd0}, _EVAL_65};
  assign _EVAL_67 = _EVAL_8[1];
  assign _EVAL_63 = {_EVAL_94,_EVAL_100,_EVAL_185,_EVAL_179};
  assign _EVAL_214 = _EVAL_19[0];
  assign _EVAL_117 = _EVAL_7[1];
  assign _EVAL_165 = _EVAL_51 == _EVAL_144;
  assign _EVAL_25 = _EVAL_125 ? _EVAL_45 : _EVAL_215;
  assign _EVAL_66 = _EVAL_88 == _EVAL_85;
  assign _EVAL_187 = _EVAL_126 | _EVAL_192;
  assign _EVAL_121 = _EVAL_210 ? _EVAL_5 : _EVAL_104;
  assign _EVAL_172 = _EVAL_29 >= _EVAL_21;
  assign _EVAL_99 = _EVAL_156 ? _EVAL_60 : _EVAL_66;
  assign _EVAL_140 = _EVAL_188 & _EVAL_190;
  assign _EVAL_60 = _EVAL_47 ^ _EVAL_130;
  assign _EVAL_152 = _EVAL_105 ? _EVAL_174 : _EVAL_44;
  assign _EVAL_120 = _EVAL_220 ? _EVAL_32 : _EVAL_119;
  assign _EVAL_89 = _EVAL_31[1];
  assign _EVAL_128 = _EVAL_180 >> _EVAL_42;
  assign _EVAL_211 = _EVAL_163 & _EVAL_38;
  assign _EVAL_61 = _EVAL_19[1];
  assign _EVAL_114 = _EVAL_101 ^ _EVAL_130;
  assign _EVAL_203 = _EVAL_118 >> _EVAL_42;
  assign _EVAL_174 = ~_EVAL_5;
  assign _EVAL_147 = _EVAL_76 & _EVAL_59;
  assign _EVAL_218 = _EVAL_81 & _EVAL_13;
  assign _EVAL_171 = _EVAL_210 ? _EVAL_174 : _EVAL_139;
  assign _EVAL_220 = _EVAL_123 & _EVAL_108;
  assign _EVAL_219 = _EVAL_105 ? _EVAL_5 : _EVAL_131;
  assign _EVAL_97 = _EVAL_56 | _EVAL_135;
  assign _EVAL_46 = _EVAL_75 & _EVAL_89;
  assign _EVAL_95 = _EVAL[2];
  assign _EVAL_47 = _EVAL_23 >= _EVAL_31;
  assign _EVAL_112 = _EVAL_7[0];
  assign _EVAL_201 = _EVAL_79[0];
  assign _EVAL_212 = _EVAL_71 | _EVAL_138;
  assign _EVAL_144 = _EVAL_166 | _EVAL_194;
  assign _EVAL_85 = _EVAL_173 | _EVAL_192;
  assign _EVAL_186 = {_EVAL_111,_EVAL_49,_EVAL_132,_EVAL_112};
  assign _EVAL_178 = _EVAL_74 | _EVAL_197;
  assign _EVAL_131 = _EVAL_202 & _EVAL_13;
  assign _EVAL_75 = _EVAL_130 & _EVAL_150;
  assign _EVAL_157 = {_EVAL_36,1'h0,1'h0,_EVAL_27};
  assign _EVAL_68 = _EVAL_74 & _EVAL_175;
  assign _EVAL_100 = _EVAL_185 & _EVAL_124;
  assign _EVAL_184 = ~_EVAL_21;
  assign _EVAL_2 = _EVAL_147 ? _EVAL_45 : _EVAL_133;
  assign _EVAL_130 = _EVAL_18[0];
  assign _EVAL_111 = _EVAL_49 & _EVAL_52;
  assign _EVAL_62 = _EVAL_211 & _EVAL_99;
  assign _EVAL_91 = _EVAL_198 & _EVAL_77;
  assign _EVAL_180 = {_EVAL_0,1'h0,1'h0,_EVAL_16};
  assign _EVAL_59 = _EVAL_204 | _EVAL_62;
  assign _EVAL_52 = _EVAL_21[2];
  assign _EVAL_69 = {{28'd0}, _EVAL_186};
  assign _EVAL_192 = {{28'd0}, _EVAL_183};
  assign _EVAL_119 = _EVAL_196 ? _EVAL_5 : _EVAL_218;
  assign _EVAL_143 = ~_EVAL_32;
  assign _EVAL_175 = _EVAL_209 & _EVAL_155;
  assign _EVAL_78 = _EVAL_56 | _EVAL_164;
  assign _EVAL_193 = _EVAL_204 & _EVAL_145;
  assign _EVAL_125 = _EVAL_98 & _EVAL_107;
  assign _EVAL_55 = _EVAL_81 & _EVAL_70;
  assign _EVAL_92 = _EVAL_72 & _EVAL_48;
  assign _EVAL_161 = _EVAL_191 == _EVAL_103;
  assign _EVAL_206 = _EVAL_113 == _EVAL_103;
  assign _EVAL_73 = _EVAL_163 & _EVAL_1;
  assign _EVAL_223 = _EVAL_207 | _EVAL_194;
  assign _EVAL_81 = _EVAL_56 & _EVAL_57;
  assign _EVAL_83 = _EVAL_140 & _EVAL_26;
  assign _EVAL_136 = _EVAL_61 ? _EVAL_216 : _EVAL_208;
  assign _EVAL_189 = _EVAL_90 == _EVAL_212;
  assign _EVAL_154 = _EVAL_53 ^ _EVAL_179;
  assign _EVAL_133 = _EVAL_205 ? _EVAL_143 : _EVAL_171;
  assign _EVAL_188 = ~_EVAL_11;
  assign _EVAL_53 = _EVAL_29 >= _EVAL;
  assign _EVAL_149 = _EVAL_160 ^ _EVAL_179;
  assign _EVAL_151 = _EVAL_23 >= _EVAL_21;
  assign _EVAL_202 = _EVAL_56 & _EVAL_164;
  assign _EVAL_82 = _EVAL_140 & _EVAL_41;
  assign _EVAL_109 = _EVAL_23 >= _EVAL_8;
  assign _EVAL_49 = _EVAL_132 & _EVAL_226;
  assign _EVAL_84 = _EVAL_204 | _EVAL_141;
  assign _EVAL_164 = _EVAL_93 & _EVAL_136;
  assign _EVAL_94 = _EVAL_100 & _EVAL_95;
  assign _EVAL_56 = ~_EVAL_20;
  assign _EVAL_226 = _EVAL_21[1];
  assign _EVAL_145 = _EVAL_73 & _EVAL_169;
  assign _EVAL_176 = _EVAL_74 | _EVAL_175;
  assign _EVAL_44 = _EVAL_202 & _EVAL_70;
  assign _EVAL_173 = ~_EVAL_31;
  assign _EVAL_153 = _EVAL[0];
  assign _EVAL_122 = _EVAL_64 & _EVAL_10;
  assign _EVAL_71 = ~_EVAL_8;
  assign _EVAL_65 = {_EVAL_92,_EVAL_72,_EVAL_127,_EVAL_214};
  assign _EVAL_181 = _EVAL_220 ? _EVAL_143 : _EVAL_148;
  assign _EVAL_58 = _EVAL_204 & _EVAL_62;
  assign _EVAL_159 = _EVAL_117 ? _EVAL_213 : _EVAL_161;
  assign _EVAL_104 = _EVAL_102 & _EVAL_13;
  assign _EVAL_64 = _EVAL_188 & _EVAL_201;
  assign _EVAL_88 = _EVAL_207 | _EVAL_192;
  assign _EVAL_127 = _EVAL_214 & _EVAL_96;
  assign _EVAL_194 = {{28'd0}, _EVAL_63};
  assign _EVAL_87 = _EVAL_128[0];
  assign _EVAL_9 = _EVAL_147 ? _EVAL_40 : _EVAL_137;
  assign _EVAL_207 = ~_EVAL_23;
  assign _EVAL_6 = _EVAL_125 ? _EVAL_40 : _EVAL_146;
  assign _EVAL_204 = ~_EVAL_17;
  assign _EVAL_93 = _EVAL_50 & _EVAL_12;
  assign _EVAL_156 = _EVAL_18[1];
  assign _EVAL_135 = _EVAL_106 & _EVAL_182;
  assign _EVAL_215 = _EVAL_129 ? _EVAL_143 : _EVAL_152;
  assign _EVAL_150 = _EVAL_31[0];
  assign _EVAL_167 = _EVAL_172 ^ _EVAL_112;
  assign _EVAL_217 = _EVAL_74 & _EVAL_142;
  assign _EVAL_126 = ~_EVAL_29;
  assign _EVAL_160 = _EVAL_23 >= _EVAL;
  assign _EVAL_166 = ~_EVAL;
  assign _EVAL_185 = _EVAL_179 & _EVAL_153;
  assign _EVAL_106 = _EVAL_50 & _EVAL_22;
  assign _EVAL_108 = _EVAL_74 | _EVAL_142;
  assign _EVAL_48 = _EVAL_8[2];
  assign _EVAL_183 = {_EVAL_110,_EVAL_46,_EVAL_75,_EVAL_130};
  assign _EVAL_103 = _EVAL_184 | _EVAL_69;
  assign _EVAL_170 = _EVAL_34[1];
  assign _EVAL_146 = _EVAL_129 ? _EVAL_32 : _EVAL_219;
  assign _EVAL_208 = _EVAL_195 == _EVAL_212;
  assign _EVAL_86 = _EVAL_109 ^ _EVAL_214;
  assign _EVAL_51 = _EVAL_126 | _EVAL_194;
  assign _EVAL_28 = _EVAL_116 ? _EVAL_40 : _EVAL_120;
  assign _EVAL_195 = _EVAL_126 | _EVAL_138;
  assign _EVAL_57 = _EVAL_162 & _EVAL_136;
  assign _EVAL_222 = _EVAL_187 == _EVAL_85;
  assign _EVAL_221 = {_EVAL_24,1'h0,1'h0,_EVAL_4};
  assign _EVAL_129 = _EVAL_193 & _EVAL_176;
  assign _EVAL_200 = _EVAL_223 == _EVAL_144;
  assign _EVAL_45 = ~_EVAL_40;
  assign _EVAL_213 = _EVAL_151 ^ _EVAL_112;
  assign _EVAL_139 = _EVAL_102 & _EVAL_70;
  assign _EVAL_134 = _EVAL_157 >> _EVAL_42;
  assign _EVAL_205 = _EVAL_58 & _EVAL_178;
  assign _EVAL_137 = _EVAL_205 ? _EVAL_32 : _EVAL_121;
  assign _EVAL_177 = _EVAL_74 & _EVAL_197;
  assign _EVAL_182 = _EVAL_61 ? _EVAL_86 : _EVAL_189;
  assign _EVAL_50 = _EVAL_188 & _EVAL_87;
  assign _EVAL_225 = _EVAL_56 | _EVAL_57;
  assign _EVAL_74 = ~_EVAL_30;
  assign _EVAL_102 = _EVAL_56 & _EVAL_135;
  assign _EVAL_190 = _EVAL_134[0];
  assign _EVAL_155 = _EVAL_117 ? _EVAL_167 : _EVAL_206;
  assign _EVAL_168 = _EVAL_31[2];
  assign _EVAL_224 = _EVAL_64 & _EVAL_43;
  assign _EVAL_199 = _EVAL_163 & _EVAL_35;
  assign _EVAL_79 = _EVAL_221 >> _EVAL_42;
  assign _EVAL_210 = _EVAL_177 & _EVAL_97;
  assign _EVAL_197 = _EVAL_224 & _EVAL_159;
  assign _EVAL_70 = ~_EVAL_13;
  assign _EVAL_77 = _EVAL_170 ? _EVAL_154 : _EVAL_165;
  assign _EVAL_96 = _EVAL_8[0];
  assign _EVAL_101 = _EVAL_29 >= _EVAL_31;
  assign _EVAL_80 = _EVAL_203[0];
  assign _EVAL_148 = _EVAL_196 ? _EVAL_174 : _EVAL_55;
  assign _EVAL_142 = _EVAL_122 & _EVAL_155;
  assign _EVAL_216 = _EVAL_115 ^ _EVAL_214;
  assign _EVAL_124 = _EVAL[1];
  assign _EVAL_162 = _EVAL_50 & _EVAL_39;
  assign _EVAL_76 = _EVAL_83 & _EVAL_54;
  assign _EVAL_191 = _EVAL_207 | _EVAL_69;
  assign _EVAL_132 = _EVAL_112 & _EVAL_158;
  assign _EVAL_110 = _EVAL_46 & _EVAL_168;
endmodule
