//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
module _EVAL_33(
  output [7:0]  _EVAL,
  output        _EVAL_0,
  output [2:0]  _EVAL_1,
  input         _EVAL_2,
  input  [3:0]  _EVAL_3,
  output [3:0]  _EVAL_4,
  input         _EVAL_5,
  input         _EVAL_6,
  output        _EVAL_7,
  output        _EVAL_8,
  input  [31:0] _EVAL_9,
  output        _EVAL_10,
  input  [3:0]  _EVAL_11,
  input  [2:0]  _EVAL_12,
  output        _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  output [31:0] _EVAL_16,
  input         _EVAL_17,
  output        _EVAL_18,
  input         _EVAL_19,
  input  [7:0]  _EVAL_20,
  input         _EVAL_21,
  output [3:0]  _EVAL_22,
  input  [2:0]  _EVAL_23,
  output [31:0] _EVAL_24,
  input  [31:0] _EVAL_25,
  input         _EVAL_26,
  input  [1:0]  _EVAL_27
);
  wire  widget__EVAL;
  wire [1:0] widget__EVAL_0;
  wire  widget__EVAL_1;
  wire [7:0] widget__EVAL_2;
  wire [7:0] widget__EVAL_3;
  wire [3:0] widget__EVAL_4;
  wire  widget__EVAL_5;
  wire [2:0] widget__EVAL_6;
  wire [3:0] widget__EVAL_7;
  wire [2:0] widget__EVAL_8;
  wire  widget__EVAL_9;
  wire  widget__EVAL_10;
  wire  widget__EVAL_11;
  wire  widget__EVAL_12;
  wire  widget__EVAL_13;
  wire  widget__EVAL_14;
  wire  widget__EVAL_15;
  wire  widget__EVAL_16;
  wire [31:0] widget__EVAL_17;
  wire [31:0] widget__EVAL_18;
  wire  widget__EVAL_19;
  wire  widget__EVAL_20;
  wire  widget__EVAL_21;
  wire  widget__EVAL_22;
  wire [3:0] widget__EVAL_23;
  wire [31:0] widget__EVAL_24;
  wire [3:0] widget__EVAL_25;
  wire [2:0] widget__EVAL_26;
  wire [31:0] widget__EVAL_27;
  _EVAL_32 widget (
    ._EVAL(widget__EVAL),
    ._EVAL_0(widget__EVAL_0),
    ._EVAL_1(widget__EVAL_1),
    ._EVAL_2(widget__EVAL_2),
    ._EVAL_3(widget__EVAL_3),
    ._EVAL_4(widget__EVAL_4),
    ._EVAL_5(widget__EVAL_5),
    ._EVAL_6(widget__EVAL_6),
    ._EVAL_7(widget__EVAL_7),
    ._EVAL_8(widget__EVAL_8),
    ._EVAL_9(widget__EVAL_9),
    ._EVAL_10(widget__EVAL_10),
    ._EVAL_11(widget__EVAL_11),
    ._EVAL_12(widget__EVAL_12),
    ._EVAL_13(widget__EVAL_13),
    ._EVAL_14(widget__EVAL_14),
    ._EVAL_15(widget__EVAL_15),
    ._EVAL_16(widget__EVAL_16),
    ._EVAL_17(widget__EVAL_17),
    ._EVAL_18(widget__EVAL_18),
    ._EVAL_19(widget__EVAL_19),
    ._EVAL_20(widget__EVAL_20),
    ._EVAL_21(widget__EVAL_21),
    ._EVAL_22(widget__EVAL_22),
    ._EVAL_23(widget__EVAL_23),
    ._EVAL_24(widget__EVAL_24),
    ._EVAL_25(widget__EVAL_25),
    ._EVAL_26(widget__EVAL_26),
    ._EVAL_27(widget__EVAL_27)
  );
  assign _EVAL_8 = widget__EVAL_11;
  assign widget__EVAL_22 = _EVAL_14;
  assign _EVAL_7 = widget__EVAL_15;
  assign widget__EVAL_3 = _EVAL_20;
  assign widget__EVAL_19 = _EVAL_17;
  assign widget__EVAL_26 = _EVAL_12;
  assign widget__EVAL_12 = _EVAL_6;
  assign _EVAL = widget__EVAL_2;
  assign widget__EVAL_5 = _EVAL_5;
  assign widget__EVAL_14 = _EVAL_26;
  assign _EVAL_1 = widget__EVAL_6;
  assign _EVAL_0 = widget__EVAL_9;
  assign _EVAL_4 = widget__EVAL_25;
  assign _EVAL_10 = widget__EVAL_10;
  assign _EVAL_18 = widget__EVAL_21;
  assign widget__EVAL = _EVAL_21;
  assign widget__EVAL_20 = _EVAL_15;
  assign _EVAL_16 = widget__EVAL_17;
  assign widget__EVAL_1 = _EVAL_2;
  assign widget__EVAL_8 = _EVAL_23;
  assign _EVAL_13 = widget__EVAL_13;
  assign widget__EVAL_27 = _EVAL_25;
  assign widget__EVAL_23 = _EVAL_11;
  assign widget__EVAL_16 = _EVAL_19;
  assign _EVAL_22 = widget__EVAL_7;
  assign widget__EVAL_24 = _EVAL_9;
  assign widget__EVAL_4 = _EVAL_3;
  assign _EVAL_24 = widget__EVAL_18;
  assign widget__EVAL_0 = _EVAL_27;
endmodule
