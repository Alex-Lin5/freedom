//
// Copyright (c) 2016-2020 SiFive, Inc. -- Proprietary and Confidential
// All Rights Reserved.
//
// NOTICE: All information contained herein is, and remains the
// property of SiFive, Inc. The intellectual and technical concepts
// contained herein are proprietary to SiFive, Inc. and may be covered
// by U.S. and Foreign Patents, patents in process, and are protected by
// trade secret or copyright law.
//
// This work may not be copied, modified, re-published, uploaded,
// executed, or distributed in any way, in any medium, whether in whole
// or in part, without prior written permission from SiFive, Inc.
//
// The copyright notice above does not evidence any actual or intended
// publication or disclosure of this source code, which includes
// information that is confidential and/or proprietary, and is a trade
// secret, of SiFive, Inc.
//
// Instance ID: 3182346c-d10e-418d-aa89-6f3d35a9b6fb, 00000000-0000-0000-0000-000000000000, 00000000-0000-0000-0000-000000000000
//VCS coverage exclude_file
module _EVAL_1_assert(
  input         _EVAL,
  input         _EVAL_0,
  input  [1:0]  _EVAL_1,
  input  [2:0]  _EVAL_2,
  input         _EVAL_3,
  input         _EVAL_4,
  input  [3:0]  _EVAL_5,
  input  [31:0] _EVAL_6,
  input  [2:0]  _EVAL_7,
  input         _EVAL_8,
  input         _EVAL_9,
  input  [3:0]  _EVAL_10,
  input         _EVAL_11,
  input  [2:0]  _EVAL_12,
  input         _EVAL_13,
  input         _EVAL_14,
  input         _EVAL_15,
  input         _EVAL_16,
  input  [3:0]  _EVAL_17,
  input         _EVAL_18
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  _EVAL_19;
  reg [2:0] _EVAL_20;
  wire [1:0] _EVAL_21;
  wire [6:0] _EVAL_22;
  wire  _EVAL_23;
  wire  _EVAL_24;
  wire [5:0] _EVAL_25;
  reg [3:0] _EVAL_26;
  wire [7:0] _EVAL_27;
  wire  _EVAL_28;
  wire  _EVAL_29;
  wire  _EVAL_30;
  wire [32:0] _EVAL_31;
  wire  _EVAL_32;
  wire  _EVAL_33;
  wire  _EVAL_34;
  reg  _EVAL_35;
  wire  _EVAL_36;
  wire  _EVAL_37;
  wire  _EVAL_38;
  wire [32:0] _EVAL_39;
  wire  _EVAL_40;
  wire  _EVAL_41;
  wire  _EVAL_42;
  wire [6:0] _EVAL_43;
  wire  _EVAL_44;
  wire [32:0] _EVAL_45;
  wire  _EVAL_46;
  wire  _EVAL_47;
  wire  _EVAL_48;
  wire [31:0] _EVAL_49;
  wire  _EVAL_50;
  wire [6:0] _EVAL_51;
  wire  _EVAL_52;
  wire [32:0] _EVAL_53;
  wire [32:0] _EVAL_54;
  wire  _EVAL_55;
  wire  _EVAL_56;
  wire  _EVAL_57;
  wire  _EVAL_58;
  wire  _EVAL_59;
  wire  _EVAL_61;
  wire [5:0] _EVAL_62;
  wire  _EVAL_63;
  wire [32:0] _EVAL_64;
  wire  _EVAL_65;
  wire  _EVAL_66;
  wire  _EVAL_67;
  wire  _EVAL_68;
  wire  _EVAL_69;
  wire  _EVAL_70;
  wire [1:0] _EVAL_71;
  wire  _EVAL_72;
  wire  _EVAL_73;
  wire  _EVAL_74;
  wire  _EVAL_75;
  wire  _EVAL_76;
  wire [32:0] _EVAL_77;
  wire  _EVAL_78;
  wire  _EVAL_79;
  wire  _EVAL_80;
  wire [32:0] _EVAL_81;
  wire  _EVAL_82;
  wire  _EVAL_83;
  wire [22:0] _EVAL_84;
  wire  _EVAL_86;
  wire  _EVAL_87;
  wire  _EVAL_88;
  wire  _EVAL_89;
  wire  _EVAL_90;
  wire  _EVAL_91;
  wire [1:0] _EVAL_92;
  wire  _EVAL_93;
  wire  _EVAL_94;
  wire  _EVAL_95;
  wire  _EVAL_96;
  wire  _EVAL_98;
  wire  _EVAL_99;
  wire  _EVAL_100;
  wire  _EVAL_101;
  wire  _EVAL_102;
  wire [1:0] _EVAL_103;
  wire  _EVAL_104;
  wire  _EVAL_105;
  wire [32:0] _EVAL_106;
  wire  _EVAL_107;
  wire  _EVAL_108;
  wire  _EVAL_110;
  wire [1:0] _EVAL_111;
  wire  _EVAL_112;
  wire  _EVAL_113;
  wire [31:0] _EVAL_114;
  wire [1:0] _EVAL_115;
  wire  _EVAL_116;
  wire  _EVAL_117;
  wire [32:0] _EVAL_118;
  wire  _EVAL_119;
  wire [32:0] _EVAL_120;
  wire [32:0] _EVAL_121;
  reg [2:0] _EVAL_122;
  wire  _EVAL_123;
  wire  _EVAL_124;
  wire  _EVAL_125;
  wire [31:0] _EVAL_126;
  wire  _EVAL_127;
  wire  _EVAL_128;
  wire  _EVAL_129;
  wire [5:0] _EVAL_130;
  wire [32:0] _EVAL_131;
  wire  _EVAL_132;
  wire  _EVAL_133;
  wire [7:0] _EVAL_134;
  wire  _EVAL_135;
  wire  _EVAL_137;
  wire [1:0] _EVAL_138;
  wire  _EVAL_139;
  wire  _EVAL_140;
  wire  _EVAL_142;
  wire [1:0] _EVAL_143;
  wire  _EVAL_144;
  wire  _EVAL_145;
  wire  _EVAL_146;
  wire  _EVAL_147;
  wire  _EVAL_148;
  wire  _EVAL_149;
  wire  _EVAL_150;
  wire [31:0] _EVAL_151;
  wire  _EVAL_152;
  wire  _EVAL_153;
  wire  _EVAL_154;
  wire [32:0] _EVAL_155;
  wire [1:0] _EVAL_156;
  wire  _EVAL_157;
  wire  _EVAL_158;
  wire  _EVAL_159;
  wire  _EVAL_160;
  wire  _EVAL_161;
  wire [32:0] _EVAL_162;
  wire  _EVAL_163;
  wire  _EVAL_164;
  wire  _EVAL_165;
  wire  _EVAL_166;
  wire  _EVAL_167;
  wire  _EVAL_168;
  wire  _EVAL_169;
  wire [6:0] _EVAL_170;
  wire  _EVAL_171;
  wire  _EVAL_172;
  wire  _EVAL_173;
  wire  _EVAL_174;
  wire  _EVAL_175;
  wire  _EVAL_176;
  wire [31:0] _EVAL_177;
  wire  _EVAL_178;
  wire  _EVAL_179;
  wire  _EVAL_180;
  wire [31:0] _EVAL_181;
  wire [32:0] _EVAL_182;
  wire  _EVAL_183;
  wire  _EVAL_184;
  wire  _EVAL_185;
  wire  _EVAL_186;
  reg [2:0] _EVAL_187;
  wire [31:0] _EVAL_189;
  wire  _EVAL_190;
  wire  _EVAL_191;
  wire [31:0] _EVAL_192;
  wire  _EVAL_193;
  wire [32:0] _EVAL_194;
  wire [32:0] _EVAL_195;
  wire  _EVAL_196;
  wire  _EVAL_197;
  wire  _EVAL_198;
  wire  _EVAL_199;
  wire [32:0] _EVAL_200;
  wire  _EVAL_201;
  wire  _EVAL_202;
  wire  _EVAL_203;
  reg [5:0] _EVAL_204;
  reg [5:0] _EVAL_205;
  wire  _EVAL_206;
  wire  _EVAL_207;
  wire  _EVAL_208;
  wire [22:0] _EVAL_210;
  wire  _EVAL_211;
  reg [31:0] _EVAL_212;
  wire  _EVAL_213;
  wire  _EVAL_214;
  wire  _EVAL_215;
  wire  _EVAL_216;
  wire  _EVAL_217;
  wire [32:0] _EVAL_218;
  wire  _EVAL_219;
  wire  _EVAL_220;
  wire  _EVAL_222;
  wire  _EVAL_223;
  wire  _EVAL_224;
  wire  _EVAL_225;
  wire  _EVAL_226;
  wire  _EVAL_227;
  wire  _EVAL_228;
  wire  _EVAL_229;
  wire [32:0] _EVAL_230;
  wire  _EVAL_231;
  wire [7:0] _EVAL_232;
  wire  _EVAL_233;
  wire  _EVAL_234;
  wire  _EVAL_235;
  wire [32:0] _EVAL_236;
  wire [5:0] _EVAL_237;
  wire  _EVAL_238;
  wire  _EVAL_239;
  reg [5:0] _EVAL_240;
  wire  _EVAL_241;
  wire  _EVAL_242;
  wire  _EVAL_244;
  wire  _EVAL_245;
  wire  _EVAL_246;
  wire  _EVAL_247;
  wire  _EVAL_248;
  wire [1:0] _EVAL_249;
  wire  _EVAL_250;
  wire  _EVAL_251;
  wire  _EVAL_252;
  wire  _EVAL_253;
  wire  _EVAL_254;
  wire  _EVAL_255;
  wire  _EVAL_257;
  wire [5:0] _EVAL_258;
  wire  _EVAL_259;
  wire  _EVAL_260;
  wire [7:0] _EVAL_261;
  wire  _EVAL_262;
  reg [1:0] _EVAL_263;
  wire  _EVAL_264;
  wire  _EVAL_265;
  wire  _EVAL_266;
  wire  _EVAL_267;
  wire  _EVAL_268;
  wire  _EVAL_269;
  wire  _EVAL_270;
  wire  _EVAL_271;
  wire  _EVAL_272;
  wire  _EVAL_273;
  wire  _EVAL_274;
  wire  _EVAL_275;
  wire  _EVAL_276;
  wire [1:0] _EVAL_277;
  wire  _EVAL_278;
  wire [32:0] _EVAL_279;
  wire  _EVAL_280;
  wire  _EVAL_281;
  wire  _EVAL_282;
  wire  _EVAL_283;
  wire  _EVAL_284;
  reg  _EVAL_285;
  wire  _EVAL_286;
  reg [31:0] _EVAL_287;
  wire  _EVAL_288;
  wire  _EVAL_289;
  reg [1:0] _EVAL_290;
  wire  _EVAL_291;
  wire  _EVAL_292;
  wire  _EVAL_293;
  wire [32:0] _EVAL_294;
  wire [3:0] _EVAL_295;
  wire  _EVAL_296;
  wire  _EVAL_297;
  wire  _EVAL_298;
  wire  _EVAL_299;
  wire  _EVAL_300;
  wire  _EVAL_301;
  reg [5:0] _EVAL_302;
  wire  _EVAL_303;
  wire  _EVAL_304;
  wire  _EVAL_305;
  wire  _EVAL_306;
  wire  _EVAL_307;
  wire  _EVAL_308;
  wire  _EVAL_309;
  wire  _EVAL_310;
  reg  _EVAL_311;
  wire  _EVAL_312;
  wire  _EVAL_313;
  wire [5:0] _EVAL_314;
  wire  _EVAL_315;
  wire  _EVAL_316;
  wire [31:0] _EVAL_317;
  wire  _EVAL_318;
  wire  _EVAL_319;
  wire  _EVAL_320;
  wire  _EVAL_321;
  wire  _EVAL_322;
  wire  _EVAL_323;
  wire  _EVAL_324;
  wire [31:0] _EVAL_325;
  reg [3:0] _EVAL_326;
  wire  _EVAL_327;
  wire  _EVAL_328;
  wire [1:0] _EVAL_329;
  wire  _EVAL_330;
  wire  _EVAL_331;
  wire  _EVAL_332;
  wire  _EVAL_333;
  wire  _EVAL_334;
  wire [32:0] _EVAL_335;
  wire [3:0] _EVAL_336;
  wire [31:0] plusarg_reader_out;
  wire  _EVAL_337;
  wire [3:0] _EVAL_338;
  wire  _EVAL_339;
  wire  _EVAL_340;
  wire  _EVAL_341;
  wire  _EVAL_342;
  wire  _EVAL_343;
  wire  _EVAL_344;
  wire  _EVAL_345;
  wire [3:0] _EVAL_346;
  reg  _EVAL_347;
  wire  _EVAL_348;
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0), .WIDTH(32)) plusarg_reader (
    .out(plusarg_reader_out)
  );
  assign _EVAL_30 = _EVAL_298 | _EVAL_305;
  assign _EVAL_180 = ~_EVAL_163;
  assign _EVAL_283 = _EVAL_17 <= 4'h2;
  assign _EVAL_74 = _EVAL_317 == 32'h0;
  assign _EVAL_40 = _EVAL_58 | _EVAL_29;
  assign _EVAL_83 = _EVAL & _EVAL_110;
  assign _EVAL_245 = ~_EVAL_251;
  assign _EVAL_69 = _EVAL_12 <= 3'h1;
  assign _EVAL_329 = 2'h1 << _EVAL_0;
  assign _EVAL_81 = $signed(_EVAL_279) & -33'sh10000;
  assign _EVAL_291 = _EVAL_71[1];
  assign _EVAL_50 = ~_EVAL_75;
  assign _EVAL_265 = _EVAL_268 & _EVAL_334;
  assign _EVAL_157 = _EVAL_3 & _EVAL_316;
  assign _EVAL_98 = ~_EVAL_273;
  assign _EVAL_19 = _EVAL_332 | _EVAL_8;
  assign _EVAL_36 = _EVAL_331 | _EVAL_8;
  assign _EVAL_127 = plusarg_reader_out == 32'h0;
  assign _EVAL_52 = _EVAL_7[0];
  assign _EVAL_34 = _EVAL_238 | _EVAL_8;
  assign _EVAL_348 = ~_EVAL_250;
  assign _EVAL_76 = _EVAL_108 & _EVAL_57;
  assign _EVAL_270 = ~_EVAL_44;
  assign _EVAL_140 = _EVAL_191 | _EVAL_127;
  assign _EVAL_120 = _EVAL_53;
  assign _EVAL_210 = 23'hff << _EVAL_10;
  assign _EVAL_296 = ~_EVAL_312;
  assign _EVAL_328 = _EVAL_47 | _EVAL_8;
  assign _EVAL_42 = _EVAL_7 <= 3'h6;
  assign _EVAL_321 = ~_EVAL_73;
  assign _EVAL_27 = _EVAL_210[7:0];
  assign _EVAL_336 = _EVAL_5 & _EVAL_346;
  assign _EVAL_153 = _EVAL_10 == _EVAL_26;
  assign _EVAL_340 = _EVAL_17 == _EVAL_326;
  assign _EVAL_183 = _EVAL_12 <= 3'h3;
  assign _EVAL_189 = _EVAL_6 ^ 32'hc000000;
  assign _EVAL_310 = _EVAL_295 == 4'h0;
  assign _EVAL_190 = ~_EVAL_199;
  assign _EVAL_119 = _EVAL_42 | _EVAL_8;
  assign _EVAL_235 = _EVAL_3 & _EVAL_61;
  assign _EVAL_114 = _EVAL_6 ^ 32'h2000000;
  assign _EVAL_67 = _EVAL_70 | _EVAL_165;
  assign _EVAL_123 = _EVAL_233 & _EVAL_265;
  assign _EVAL_156 = _EVAL_290 | _EVAL_143;
  assign _EVAL_113 = ~_EVAL_82;
  assign _EVAL_169 = _EVAL_3 & _EVAL_135;
  assign _EVAL_305 = $signed(_EVAL_31) == 33'sh0;
  assign _EVAL_171 = _EVAL_183 | _EVAL_8;
  assign _EVAL_308 = _EVAL_300 | _EVAL_108;
  assign _EVAL_80 = _EVAL_300 & _EVAL_91;
  assign _EVAL_56 = ~_EVAL_46;
  assign _EVAL_53 = $signed(_EVAL_194) & -33'sh4000;
  assign _EVAL_148 = _EVAL_96 | _EVAL_29;
  assign _EVAL_184 = _EVAL_340 | _EVAL_8;
  assign _EVAL_59 = _EVAL_167 | _EVAL_8;
  assign _EVAL_128 = _EVAL_3 & _EVAL_95;
  assign _EVAL_31 = _EVAL_54;
  assign _EVAL_100 = _EVAL_300 & _EVAL_276;
  assign _EVAL_99 = ~_EVAL_186;
  assign _EVAL_343 = _EVAL_1 == 2'h0;
  assign _EVAL_227 = _EVAL_173 | _EVAL_8;
  assign _EVAL_314 = _EVAL_170[5:0];
  assign _EVAL_242 = _EVAL_309 & _EVAL_334;
  assign _EVAL_272 = ~_EVAL_125;
  assign _EVAL_106 = $signed(_EVAL_195) & -33'sh2000;
  assign _EVAL_139 = _EVAL_17 <= 4'h8;
  assign _EVAL_58 = $signed(_EVAL_39) == 33'sh0;
  assign _EVAL_47 = _EVAL_262 | _EVAL_254;
  assign _EVAL_333 = _EVAL_291 & _EVAL_309;
  assign _EVAL_249 = _EVAL_257 ? _EVAL_138 : 2'h0;
  assign _EVAL_191 = ~_EVAL_318;
  assign _EVAL_216 = $signed(_EVAL_120) == 33'sh0;
  assign _EVAL_294 = _EVAL_81;
  assign _EVAL_160 = ~_EVAL_253;
  assign _EVAL_254 = _EVAL_267 & _EVAL_159;
  assign _EVAL_88 = _EVAL_2[2];
  assign _EVAL_248 = ~_EVAL_158;
  assign _EVAL_43 = _EVAL_302 - 6'h1;
  assign _EVAL_29 = $signed(_EVAL_45) == 33'sh0;
  assign _EVAL_234 = _EVAL_2 == 3'h3;
  assign _EVAL_182 = $signed(_EVAL_230) & -33'sh2000;
  assign _EVAL_318 = |_EVAL_290;
  assign _EVAL_281 = _EVAL & _EVAL_255;
  assign _EVAL_87 = _EVAL_149 | _EVAL_8;
  assign _EVAL_90 = _EVAL_17 <= 4'hb;
  assign _EVAL_344 = ~_EVAL_129;
  assign _EVAL_86 = _EVAL_309 & _EVAL_260;
  assign _EVAL_105 = _EVAL_72 | _EVAL_8;
  assign _EVAL_288 = ~_EVAL_0;
  assign _EVAL_293 = _EVAL_267 & _EVAL_40;
  assign _EVAL_91 = _EVAL_240 == 6'h0;
  assign _EVAL_306 = _EVAL_0 == _EVAL_311;
  assign _EVAL_101 = _EVAL_2 == 3'h0;
  assign _EVAL_107 = _EVAL_70 | _EVAL_286;
  assign _EVAL_125 = |_EVAL_143;
  assign _EVAL_259 = ~_EVAL_184;
  assign _EVAL_23 = _EVAL_93 | _EVAL_8;
  assign _EVAL_181 = _EVAL_6 ^ 32'h40000000;
  assign _EVAL_161 = ~_EVAL_207;
  assign _EVAL_250 = _EVAL_175 | _EVAL_8;
  assign _EVAL_228 = _EVAL_268 & _EVAL_260;
  assign _EVAL_108 = _EVAL_13 & _EVAL;
  assign _EVAL_186 = _EVAL_153 | _EVAL_8;
  assign _EVAL_178 = _EVAL_90 & _EVAL_288;
  assign _EVAL_271 = ~_EVAL_8;
  assign _EVAL_48 = ~_EVAL_65;
  assign _EVAL_45 = _EVAL_106;
  assign _EVAL_64 = $signed(_EVAL_218) & -33'sh4000;
  assign _EVAL_159 = _EVAL_148 | _EVAL_216;
  assign _EVAL_252 = ~_EVAL_164;
  assign _EVAL_196 = ~_EVAL_264;
  assign _EVAL_327 = _EVAL_1 != 2'h2;
  assign _EVAL_147 = ~_EVAL_34;
  assign _EVAL_309 = ~_EVAL_268;
  assign _EVAL_146 = ~_EVAL_303;
  assign _EVAL_68 = $signed(_EVAL_294) == 33'sh0;
  assign _EVAL_126 = {{24'd0}, _EVAL_134};
  assign _EVAL_151 = _EVAL_118[31:0];
  assign _EVAL_129 = _EVAL_63 | _EVAL_8;
  assign _EVAL_32 = ~_EVAL_59;
  assign _EVAL_94 = _EVAL_3 & _EVAL_78;
  assign _EVAL_155 = _EVAL_64;
  assign _EVAL_282 = _EVAL_3 & _EVAL_297;
  assign _EVAL_104 = ~_EVAL_23;
  assign _EVAL_110 = _EVAL_7 == 3'h5;
  assign _EVAL_335 = _EVAL_131;
  assign _EVAL_276 = _EVAL_204 == 6'h0;
  assign _EVAL_231 = ~_EVAL_133;
  assign _EVAL_202 = ~_EVAL_11;
  assign _EVAL_214 = ~_EVAL_171;
  assign _EVAL_133 = _EVAL_322 | _EVAL_8;
  assign _EVAL_236 = $signed(_EVAL_121) & -33'sh1000;
  assign _EVAL_163 = _EVAL_24 | _EVAL_8;
  assign _EVAL_211 = ~_EVAL_15;
  assign _EVAL_266 = _EVAL_267 & _EVAL_320;
  assign _EVAL_39 = _EVAL_182;
  assign _EVAL_320 = _EVAL_30 | _EVAL_216;
  assign _EVAL_185 = ~_EVAL_36;
  assign _EVAL_262 = _EVAL_139 & _EVAL_152;
  assign _EVAL_275 = ~_EVAL_18;
  assign _EVAL_164 = _EVAL_327 | _EVAL_8;
  assign _EVAL_264 = _EVAL_176 | _EVAL_8;
  assign _EVAL_289 = _EVAL_3 & _EVAL_101;
  assign _EVAL_339 = ~_EVAL_203;
  assign _EVAL_207 = _EVAL_306 | _EVAL_8;
  assign _EVAL_65 = _EVAL_307 | _EVAL_8;
  assign _EVAL_66 = ~_EVAL_328;
  assign _EVAL_24 = _EVAL_12 != 3'h0;
  assign _EVAL_28 = ~_EVAL_88;
  assign _EVAL_278 = _EVAL_17[0];
  assign _EVAL_206 = _EVAL_1 == _EVAL_263;
  assign _EVAL_307 = _EVAL_15 == _EVAL_285;
  assign _EVAL_319 = _EVAL_6 == _EVAL_287;
  assign _EVAL_112 = _EVAL_277[0];
  assign _EVAL_199 = _EVAL_174 | _EVAL_8;
  assign _EVAL_292 = ~_EVAL_315;
  assign _EVAL_315 = _EVAL_198 | _EVAL_8;
  assign _EVAL_238 = _EVAL_5 == _EVAL_338;
  assign _EVAL_332 = ~_EVAL_102;
  assign _EVAL_170 = _EVAL_205 - 6'h1;
  assign _EVAL_173 = _EVAL_202 | _EVAL_18;
  assign _EVAL_301 = ~_EVAL_224;
  assign _EVAL_255 = _EVAL_7 == 3'h2;
  assign _EVAL_176 = _EVAL_93 & _EVAL_47;
  assign _EVAL_273 = _EVAL_205 == 6'h0;
  assign _EVAL_341 = ~_EVAL_79;
  assign _EVAL_277 = _EVAL_115 >> _EVAL_15;
  assign _EVAL_251 = _EVAL_179 | _EVAL_8;
  assign _EVAL_237 = _EVAL_232[7:2];
  assign _EVAL_61 = _EVAL_2 == 3'h2;
  assign _EVAL_346 = ~_EVAL_338;
  assign _EVAL_72 = ~_EVAL_16;
  assign _EVAL_22 = _EVAL_240 - 6'h1;
  assign _EVAL_241 = ~_EVAL_119;
  assign _EVAL_215 = _EVAL_112 | _EVAL_8;
  assign _EVAL_62 = _EVAL_51[5:0];
  assign _EVAL_154 = _EVAL & _EVAL_168;
  assign _EVAL_57 = _EVAL_302 == 6'h0;
  assign _EVAL_280 = _EVAL_319 | _EVAL_8;
  assign _EVAL_194 = {1'b0,$signed(_EVAL_49)};
  assign _EVAL_54 = $signed(_EVAL_77) & -33'sh400000;
  assign _EVAL_230 = {1'b0,$signed(_EVAL_177)};
  assign _EVAL_274 = _EVAL_108 & _EVAL_273;
  assign _EVAL_193 = _EVAL_202 | _EVAL_8;
  assign _EVAL_111 = _EVAL_290 >> _EVAL_0;
  assign _EVAL_145 = _EVAL_144 | _EVAL_217;
  assign _EVAL_313 = _EVAL_17 >= 4'h2;
  assign _EVAL_198 = _EVAL_15 | _EVAL_211;
  assign _EVAL_257 = _EVAL_76 & _EVAL_339;
  assign _EVAL_223 = _EVAL_12 == _EVAL_122;
  assign _EVAL_330 = ~_EVAL_19;
  assign _EVAL_201 = ~_EVAL_105;
  assign _EVAL_131 = $signed(_EVAL_162) & -33'sh5000;
  assign _EVAL_132 = $signed(_EVAL_155) == 33'sh0;
  assign _EVAL_124 = ~_EVAL_213;
  assign _EVAL_298 = _EVAL_345 | _EVAL_68;
  assign _EVAL_192 = _EVAL_6 ^ 32'h3000;
  assign _EVAL_84 = 23'hff << _EVAL_17;
  assign _EVAL_233 = _EVAL_71[0];
  assign _EVAL_268 = _EVAL_6[1];
  assign _EVAL_55 = ~_EVAL_193;
  assign _EVAL_303 = _EVAL_150 | _EVAL_8;
  assign _EVAL_130 = _EVAL_43[5:0];
  assign _EVAL_102 = _EVAL_111[0];
  assign _EVAL_279 = {1'b0,$signed(_EVAL_114)};
  assign _EVAL_325 = _EVAL_6 ^ 32'h1800000;
  assign _EVAL_220 = _EVAL_2 == 3'h7;
  assign _EVAL_41 = ~_EVAL_116;
  assign _EVAL_63 = _EVAL_10 >= 4'h2;
  assign _EVAL_46 = _EVAL_172 | _EVAL_8;
  assign _EVAL_317 = _EVAL_6 & _EVAL_126;
  assign _EVAL_144 = _EVAL_313 | _EVAL_219;
  assign _EVAL_232 = ~_EVAL_27;
  assign _EVAL_70 = _EVAL_313 | _EVAL_333;
  assign _EVAL_342 = ~_EVAL_269;
  assign _EVAL_143 = _EVAL_80 ? _EVAL_329 : 2'h0;
  assign _EVAL_226 = _EVAL_283 & _EVAL_0;
  assign _EVAL_269 = _EVAL_223 | _EVAL_8;
  assign _EVAL_219 = _EVAL_291 & _EVAL_268;
  assign _EVAL_225 = _EVAL_262 | _EVAL_293;
  assign _EVAL_267 = _EVAL_17 <= 4'h6;
  assign _EVAL_337 = _EVAL_33 | _EVAL_272;
  assign _EVAL_316 = _EVAL_2 == 3'h1;
  assign _EVAL_217 = _EVAL_233 & _EVAL_228;
  assign _EVAL_247 = _EVAL_144 | _EVAL_123;
  assign _EVAL_73 = _EVAL_206 | _EVAL_8;
  assign _EVAL_304 = ~_EVAL_324;
  assign _EVAL_165 = _EVAL_233 & _EVAL_242;
  assign _EVAL_179 = _EVAL_336 == 4'h0;
  assign _EVAL_95 = ~_EVAL_276;
  assign _EVAL_175 = _EVAL_7 == _EVAL_20;
  assign _EVAL_224 = _EVAL_313 | _EVAL_8;
  assign _EVAL_239 = _EVAL_12 <= 3'h4;
  assign _EVAL_103 = ~_EVAL_249;
  assign _EVAL_261 = _EVAL_84[7:0];
  assign _EVAL_77 = {1'b0,$signed(_EVAL_189)};
  assign _EVAL_49 = _EVAL_6 ^ 32'h80000000;
  assign _EVAL_222 = _EVAL_3 & _EVAL_220;
  assign _EVAL_71 = _EVAL_21 | 2'h1;
  assign _EVAL_75 = _EVAL_74 | _EVAL_8;
  assign _EVAL_174 = _EVAL_12 == 3'h0;
  assign _EVAL_284 = _EVAL & _EVAL_89;
  assign _EVAL_162 = {1'b0,$signed(_EVAL_6)};
  assign _EVAL_244 = ~_EVAL_280;
  assign _EVAL_300 = _EVAL_14 & _EVAL_3;
  assign _EVAL_195 = {1'b0,$signed(_EVAL_181)};
  assign _EVAL_168 = _EVAL_7 == 3'h1;
  assign _EVAL_38 = _EVAL_262 | _EVAL_266;
  assign _EVAL_121 = {1'b0,$signed(_EVAL_192)};
  assign _EVAL_117 = $signed(_EVAL_335) == 33'sh0;
  assign _EVAL_213 = _EVAL_275 | _EVAL_8;
  assign _EVAL_177 = _EVAL_6 ^ 32'h20000000;
  assign _EVAL_345 = _EVAL_117 | _EVAL_132;
  assign _EVAL_25 = _EVAL_22[5:0];
  assign _EVAL_260 = _EVAL_6[0];
  assign _EVAL_323 = _EVAL & _EVAL_203;
  assign _EVAL_92 = _EVAL_156 & _EVAL_103;
  assign _EVAL_134 = ~_EVAL_261;
  assign _EVAL_197 = _EVAL_3 & _EVAL_234;
  assign _EVAL_118 = _EVAL_212 + 32'h1;
  assign _EVAL_299 = _EVAL_1 <= 2'h2;
  assign _EVAL_78 = _EVAL_2 == 3'h6;
  assign _EVAL_331 = _EVAL_0 | _EVAL_288;
  assign _EVAL_338 = {_EVAL_145,_EVAL_247,_EVAL_107,_EVAL_67};
  assign _EVAL_152 = $signed(_EVAL_200) == 33'sh0;
  assign _EVAL_37 = _EVAL & _EVAL_98;
  assign _EVAL_158 = _EVAL_225 | _EVAL_8;
  assign _EVAL_135 = _EVAL_2 == 3'h5;
  assign _EVAL_208 = _EVAL & _EVAL_229;
  assign _EVAL_200 = _EVAL_236;
  assign _EVAL_79 = _EVAL_239 | _EVAL_8;
  assign _EVAL_33 = _EVAL_143 != _EVAL_249;
  assign _EVAL_21 = 2'h1 << _EVAL_278;
  assign _EVAL_229 = _EVAL_7 == 3'h4;
  assign _EVAL_82 = _EVAL_69 | _EVAL_8;
  assign _EVAL_203 = _EVAL_7 == 3'h6;
  assign _EVAL_93 = _EVAL_226 | _EVAL_178;
  assign _EVAL_96 = _EVAL_30 | _EVAL_58;
  assign _EVAL_246 = ~_EVAL_227;
  assign _EVAL_149 = _EVAL_140 | _EVAL_137;
  assign _EVAL_324 = _EVAL_299 | _EVAL_8;
  assign _EVAL_89 = _EVAL_7 == 3'h0;
  assign _EVAL_172 = _EVAL_4 == _EVAL_347;
  assign _EVAL_115 = _EVAL_143 | _EVAL_290;
  assign _EVAL_44 = _EVAL_337 | _EVAL_8;
  assign _EVAL_258 = _EVAL_134[7:2];
  assign _EVAL_166 = ~_EVAL_215;
  assign _EVAL_218 = {1'b0,$signed(_EVAL_325)};
  assign _EVAL_312 = _EVAL_38 | _EVAL_8;
  assign _EVAL_297 = _EVAL_2 == 3'h4;
  assign _EVAL_51 = _EVAL_204 - 6'h1;
  assign _EVAL_137 = _EVAL_212 < plusarg_reader_out;
  assign _EVAL_295 = ~_EVAL_5;
  assign _EVAL_286 = _EVAL_233 & _EVAL_86;
  assign _EVAL_253 = _EVAL_310 | _EVAL_8;
  assign _EVAL_334 = ~_EVAL_260;
  assign _EVAL_138 = 2'h1 << _EVAL_15;
  assign _EVAL_116 = _EVAL_343 | _EVAL_8;
  assign _EVAL_322 = _EVAL_12 <= 3'h2;
  assign _EVAL_150 = _EVAL_2 == _EVAL_187;
  assign _EVAL_142 = ~_EVAL_87;
  assign _EVAL_167 = _EVAL_11 == _EVAL_35;
  always @(posedge _EVAL_9) begin
    if (_EVAL_274) begin
      _EVAL_20 <= _EVAL_7;
    end
    if (_EVAL_274) begin
      _EVAL_26 <= _EVAL_10;
    end
    if (_EVAL_274) begin
      _EVAL_35 <= _EVAL_11;
    end
    if (_EVAL_100) begin
      _EVAL_122 <= _EVAL_12;
    end
    if (_EVAL_100) begin
      _EVAL_187 <= _EVAL_2;
    end
    if (_EVAL_8) begin
      _EVAL_204 <= 6'h0;
    end else if (_EVAL_300) begin
      if (_EVAL_276) begin
        if (_EVAL_28) begin
          _EVAL_204 <= _EVAL_258;
        end else begin
          _EVAL_204 <= 6'h0;
        end
      end else begin
        _EVAL_204 <= _EVAL_62;
      end
    end
    if (_EVAL_8) begin
      _EVAL_205 <= 6'h0;
    end else if (_EVAL_108) begin
      if (_EVAL_273) begin
        if (_EVAL_52) begin
          _EVAL_205 <= _EVAL_237;
        end else begin
          _EVAL_205 <= 6'h0;
        end
      end else begin
        _EVAL_205 <= _EVAL_314;
      end
    end
    if (_EVAL_8) begin
      _EVAL_212 <= 32'h0;
    end else if (_EVAL_308) begin
      _EVAL_212 <= 32'h0;
    end else begin
      _EVAL_212 <= _EVAL_151;
    end
    if (_EVAL_8) begin
      _EVAL_240 <= 6'h0;
    end else if (_EVAL_300) begin
      if (_EVAL_91) begin
        if (_EVAL_28) begin
          _EVAL_240 <= _EVAL_258;
        end else begin
          _EVAL_240 <= 6'h0;
        end
      end else begin
        _EVAL_240 <= _EVAL_25;
      end
    end
    if (_EVAL_274) begin
      _EVAL_263 <= _EVAL_1;
    end
    if (_EVAL_274) begin
      _EVAL_285 <= _EVAL_15;
    end
    if (_EVAL_100) begin
      _EVAL_287 <= _EVAL_6;
    end
    if (_EVAL_8) begin
      _EVAL_290 <= 2'h0;
    end else begin
      _EVAL_290 <= _EVAL_92;
    end
    if (_EVAL_8) begin
      _EVAL_302 <= 6'h0;
    end else if (_EVAL_108) begin
      if (_EVAL_57) begin
        if (_EVAL_52) begin
          _EVAL_302 <= _EVAL_237;
        end else begin
          _EVAL_302 <= 6'h0;
        end
      end else begin
        _EVAL_302 <= _EVAL_130;
      end
    end
    if (_EVAL_100) begin
      _EVAL_311 <= _EVAL_0;
    end
    if (_EVAL_100) begin
      _EVAL_326 <= _EVAL_17;
    end
    if (_EVAL_274) begin
      _EVAL_347 <= _EVAL_4;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b89ee5e1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_248) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(af98b544)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba0c689a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_166) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_244) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6b6ed1a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_292) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8b7b7742)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_296) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(16e2c774)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_48) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b425311f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(78dccd4d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_330) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bc5df332)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7bf91190)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_66) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d82cfb5c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a3fe0f66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_257 & _EVAL_166) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(86fe575a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_321) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b8567bdd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1d9a5927)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_292) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_146) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1716f46)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d68e1cff)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_245) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4965884b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_344) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cb74aef3)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5098eeb9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1515931c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf18667)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_66) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_99) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(12e82b18)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_142) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_270) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2cc4c8ad)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_301) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b4c43ff4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_344) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a228683e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c83bc2bb)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_48) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc92f8fe)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b61e7c11)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b3c3832c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_180) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_344) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a59fcd76)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_248) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2bac9332)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8960701a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_344) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_344) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(69c3f14e)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_246) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e09c0a1a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f27aa2a1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_304) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(126d057a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(866d1427)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8f31f87f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8c52c166)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(6c83d618)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(428a8031)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_292) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5cdc8723)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_161) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(26005506)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d488a9b2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_80 & _EVAL_330) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_252) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2ea753dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_124) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(270ee79b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_304) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(50dbcb66)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(380484fa)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_304) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(487ed2a0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_304) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db72bd6d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e2944ab2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_244) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f0c5e0ac)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(673025e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_341) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5e911f3b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_321) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_301) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_301) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(7aa4e25a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_301) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ca9c913c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_341) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_231) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_41) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a5b3da55)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_32) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_245) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a74b8f6f)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_147) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_214) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ba9d95a9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_259) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5afe4a02)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(ebcfdb69)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_113) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(1760bfe4)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_246) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL & _EVAL_241) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dc9e5fc2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(cd32edb0)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_99) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_161) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_348) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_344) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_292) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(dd1d627b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_190) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(bf40a209)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_342) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b52ab7e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_201) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_56) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(196cbe9d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_292) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(74d7a379)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_252) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_104) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4cd65140)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_113) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(925a94f2)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_55) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(20b10ecf)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_281 & _EVAL_124) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(41f888d6)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_104) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_56) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(db284749)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_154 & _EVAL_41) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_235 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_231) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8450a04a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_282 & _EVAL_147) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a9dab4af)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_83 & _EVAL_292) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_208 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL & _EVAL_241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_323 & _EVAL_55) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(d2f46065)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_185) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_196) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(77084b9)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_142) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(f68e7df8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_214) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(8bd69cdd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(4355f22a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(673025e8)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_271) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_271) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(372680bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_197 & _EVAL_185) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(a520eb5b)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_196) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_169 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(b33fb96d)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_342) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_32) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(9c823235)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_289 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(239265bd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_201) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(668c1373)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_296) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(2604591a)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_284 & _EVAL_292) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_128 & _EVAL_259) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_50) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(5c693ccd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_37 & _EVAL_348) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(c4b8a785)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_EVAL_157 & _EVAL_50) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_94 & _EVAL_160) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(e5d7f0dd)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_EVAL_222 & _EVAL_180) begin
          $fwrite(32'h80000002,"Obfuscated Simulation Output(704a3c6c)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _EVAL_20 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  _EVAL_26 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  _EVAL_35 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _EVAL_122 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  _EVAL_187 = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  _EVAL_204 = _RAND_5[5:0];
  _RAND_6 = {1{`RANDOM}};
  _EVAL_205 = _RAND_6[5:0];
  _RAND_7 = {1{`RANDOM}};
  _EVAL_212 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  _EVAL_240 = _RAND_8[5:0];
  _RAND_9 = {1{`RANDOM}};
  _EVAL_263 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  _EVAL_285 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _EVAL_287 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  _EVAL_290 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  _EVAL_302 = _RAND_13[5:0];
  _RAND_14 = {1{`RANDOM}};
  _EVAL_311 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _EVAL_326 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  _EVAL_347 = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS

endmodule
